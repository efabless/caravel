* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for mprj2_logic_high abstract view
.subckt mprj2_logic_high HI vccd2 vssd2
.ends

* Black-box entry subcircuit for mprj_logic_high abstract view
.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46]
+ HI[47] HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57]
+ HI[58] HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68]
+ HI[69] HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79]
+ HI[7] HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8]
+ HI[90] HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1
+ vssd1
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv mprj2_vdd_logic1 mprj_vdd_logic1 vccd vssd vdda1 vssa1 vdda2
+ vssa2
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd vccd1_uq1 vccd2_uq0 vdda1_uq0 vdda2_uq0 vssd vssd2_uq0
+ vssa1_uq0 vssa2_uq0 vssd1_uq1
XFILLER_3_3168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1343__B _1343_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_166 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0703__A _0703_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1237__C _1237_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1253__B _1253_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input127_A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3390 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input92_A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0613__A _0613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[8\] mprj_dat_i_user[8] _0870_/X vssd vssd vccd vccd _0584_/A sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2903 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1444__A _1444_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1270_ _1270_/A vssd vssd vccd vccd _1270_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1163__B _1163_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output513_A _1024_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output882_A _0586_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3198 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] _0658_/X vssd vssd vccd vccd _0470_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_36_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0985_ _0985_/A _0985_/B vssd vssd vccd vccd _0986_/A sky130_fd_sc_hd__and2_2
XFILLER_9_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0523__A _0523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_29_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1057__C _1057_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput467 _1226_/X vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__buf_12
Xoutput478 _1246_/X vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__buf_12
XFILLER_9_3399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput489 _1266_/X vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__buf_12
X_1537_ _1537_/A vssd vssd vccd vccd _1537_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1468_ _1468_/A vssd vssd vccd vccd _1468_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1073__B _1073_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1399_ _1399_/A _1399_/B vssd vssd vccd vccd _1400_/A sky130_fd_sc_hd__and2_4
XFILLER_27_203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1529__A _1529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_847 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1264__A _1264_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input244_A la_iena_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input411_A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1439__A _1439_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0770_ _0770_/A vssd vssd vccd vccd _0770_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output463_A _1020_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_674 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0997__B _0997_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output728_A _1492_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1174__A _1174_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1322_ _1322_/A vssd vssd vccd vccd _1322_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1253_ _1509_/A _1253_/B _1253_/C vssd vssd vccd vccd _1254_/A sky130_fd_sc_hd__and3b_2
XFILLER_0_3127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1184_ _1184_/A vssd vssd vccd vccd _1184_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0518__A _0518_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1349__A _1349_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0968_ _0968_/A vssd vssd vccd vccd _0968_/X sky130_fd_sc_hd__buf_8
XFILLER_44_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0899_ _0899_/A _0899_/B vssd vssd vccd vccd _0900_/A sky130_fd_sc_hd__and2_2
XFILLER_48_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2083 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_740 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_75 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input194_A la_iena_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2578 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input361_A la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input459_A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input55_A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3386 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1441__B _1441_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output580_A _1200_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0822_ _0822_/A vssd vssd vccd vccd _0822_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output845_A _1474_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0753_ _0753_/A _0753_/B vssd vssd vccd vccd _0754_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0801__A _0801_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0684_ _0684_/A vssd vssd vccd vccd _0684_/X sky130_fd_sc_hd__clkbuf_1
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] _0792_/X vssd vssd vccd vccd _0537_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_45_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1305_ _1305_/A _1305_/B vssd vssd vccd vccd _1306_/A sky130_fd_sc_hd__and2_4
XFILLER_42_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1236_ _1236_/A vssd vssd vccd vccd _1236_/X sky130_fd_sc_hd__buf_2
XFILLER_42_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1351__B _1351_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1167_ _1423_/A _1167_/B _1167_/C vssd vssd vccd vccd _1168_/A sky130_fd_sc_hd__and3b_1
XFILLER_39_2935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1098_ _1098_/A vssd vssd vccd vccd _1098_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1298 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0711__A _0711_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3938 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1245__C _1245_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1261__B _1261_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input207_A la_iena_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0621__A _0621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1155__C _1155_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1171__B _1171_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1021_ _1277_/A _1021_/B _1021_/C vssd vssd vccd vccd _1022_/A sky130_fd_sc_hd__and3b_2
XFILLER_47_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2598 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output795_A _1382_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[20\] mprj_dat_i_user[20] _0870_/X vssd vssd vccd vccd _0596_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_12_3853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0805_ _0805_/A _0805_/B vssd vssd vccd vccd _0806_/A sky130_fd_sc_hd__and2_4
XANTENNA__0531__A _0531_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0736_ _0736_/A vssd vssd vccd vccd _0736_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0667_ _0667_/A _0667_/B vssd vssd vccd vccd _0668_/A sky130_fd_sc_hd__and2_1
XFILLER_6_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1968 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0598_ _0598_/A vssd vssd vccd vccd _0598_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_2432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1362__A _1362_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1045__A_N _1301_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1081__B _1081_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1219_ _1475_/A _1219_/B input5/X vssd vssd vccd vccd _1220_/A sky130_fd_sc_hd__and3b_4
XTAP_2919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1195__A_N _1451_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input157_A la_iena_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput301 la_oenb_mprj[21] vssd vssd vccd vccd _1317_/A sky130_fd_sc_hd__buf_2
Xinput312 la_oenb_mprj[31] vssd vssd vccd vccd _1337_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput323 la_oenb_mprj[41] vssd vssd vccd vccd _1357_/A sky130_fd_sc_hd__buf_2
XFILLER_44_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput334 la_oenb_mprj[51] vssd vssd vccd vccd _1377_/A sky130_fd_sc_hd__clkbuf_4
Xinput345 la_oenb_mprj[61] vssd vssd vccd vccd _1397_/A sky130_fd_sc_hd__buf_2
XANTENNA__1272__A _1272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput356 la_oenb_mprj[71] vssd vssd vccd vccd _1417_/A sky130_fd_sc_hd__clkbuf_4
Xinput367 la_oenb_mprj[81] vssd vssd vccd vccd _1437_/A sky130_fd_sc_hd__buf_4
XANTENNA_input324_A la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput378 la_oenb_mprj[91] vssd vssd vccd vccd _1457_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput389 mprj_adr_o_core[10] vssd vssd vccd vccd _0911_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input18_A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1447__A _1447_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput808 _1406_/X vssd vssd vccd vccd la_oenb_core[65] sky130_fd_sc_hd__buf_12
Xoutput819 _1426_/X vssd vssd vccd vccd la_oenb_core[75] sky130_fd_sc_hd__buf_12
X_0521_ _0521_/A vssd vssd vccd vccd _0521_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] _0718_/X vssd vssd vccd vccd _0500_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_26_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1004_ _1004_/A vssd vssd vccd vccd _1004_/X sky130_fd_sc_hd__buf_6
XFILLER_1_2395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0526__A _0526_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1357__A _1357_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0719_ _0719_/A _0719_/B vssd vssd vccd vccd _0720_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1092__A _1092_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input274_A la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input441_A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput120 la_data_out_mprj[8] vssd vssd vccd vccd _1035_/C sky130_fd_sc_hd__clkbuf_1
Xinput131 la_data_out_mprj[9] vssd vssd vccd vccd _1037_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput142 la_iena_mprj[109] vssd vssd vccd vccd _0825_/B sky130_fd_sc_hd__clkbuf_4
Xinput153 la_iena_mprj[119] vssd vssd vccd vccd _0845_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput164 la_iena_mprj[13] vssd vssd vccd vccd _0633_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput175 la_iena_mprj[23] vssd vssd vccd vccd _0653_/B sky130_fd_sc_hd__clkbuf_2
Xinput186 la_iena_mprj[33] vssd vssd vccd vccd _0673_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_18_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput197 la_iena_mprj[43] vssd vssd vccd vccd _0693_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output660_A _0492_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output758_A _1278_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput605 _0557_/Y vssd vssd vccd vccd la_data_in_mprj[112] sky130_fd_sc_hd__buf_12
XFILLER_9_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput616 _0567_/Y vssd vssd vccd vccd la_data_in_mprj[122] sky130_fd_sc_hd__buf_12
XFILLER_29_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput627 _0462_/Y vssd vssd vccd vccd la_data_in_mprj[17] sky130_fd_sc_hd__buf_12
Xoutput638 _0472_/Y vssd vssd vccd vccd la_data_in_mprj[27] sky130_fd_sc_hd__buf_12
XANTENNA_output925_A _0996_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput649 _0482_/Y vssd vssd vccd vccd la_data_in_mprj[37] sky130_fd_sc_hd__buf_12
X_0504_ _0504_/A vssd vssd vccd vccd _0504_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1484_ _1484_/A vssd vssd vccd vccd _1484_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1233__A_N _1489_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0703__B _0703_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1253__C _1253_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_974 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input391_A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input85_A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0613__B _0613_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_2503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1163__C _1163_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output506_A _1066_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1460__A _1460_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output875_A _0902_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] _0644_/X vssd vssd vccd vccd _0463_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__0804__A _0804_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0984_ _0984_/A vssd vssd vccd vccd _0984_/X sky130_fd_sc_hd__buf_6
XFILLER_31_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[100\]_B _0808_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput468 _1228_/X vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__buf_12
X_1536_ _1536_/A vssd vssd vccd vccd _1536_/Y sky130_fd_sc_hd__inv_2
Xoutput479 _1248_/X vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__buf_12
XFILLER_5_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1467_ _1467_/A _1467_/B vssd vssd vccd vccd _1468_/A sky130_fd_sc_hd__and2_1
XFILLER_25_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1073__C _1073_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1398_ _1398_/A vssd vssd vccd vccd _1398_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_3760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1370__A _1370_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1529__B _1529_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1129__A_N _1385_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input237_A la_iena_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1280__A _1280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input404_A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1439__B _1439_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1455__A _1455_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2723 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1321_ _1321_/A _1321_/B vssd vssd vccd vccd _1322_/A sky130_fd_sc_hd__and2_4
XFILLER_25_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output623_A _1546_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1252_ _1252_/A vssd vssd vccd vccd _1252_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1183_ _1439_/A _1183_/B _1183_/C vssd vssd vccd vccd _1184_/A sky130_fd_sc_hd__and3b_1
XFILLER_4_2596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1190__A _1190_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0534__A _0534_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1349__B _1349_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0967_ _0967_/A _0967_/B vssd vssd vccd vccd _0968_/A sky130_fd_sc_hd__and2_1
XFILLER_31_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0898_ _0898_/A vssd vssd vccd vccd _0898_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_44_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1365__A _1365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1519_ _1519_/A _1519_/B vssd vssd vccd vccd _1520_/A sky130_fd_sc_hd__and2_1
XFILLER_26_3991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0709__A _0709_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3590 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1259__B _1259_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input187_A la_iena_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1275__A _1275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input354_A la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input48_A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0619__A _0619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1169__B _1169_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0821_ _0821_/A _0821_/B vssd vssd vccd vccd _0822_/A sky130_fd_sc_hd__and2_1
XANTENNA_output573_A _1188_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0752_ _0752_/A vssd vssd vccd vccd _0752_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0801__B _0801_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0683_ _0683_/A _0683_/B vssd vssd vccd vccd _0684_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] _0778_/X vssd vssd vccd vccd _0530_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1304_ _1304_/A vssd vssd vccd vccd _1304_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_3061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0529__A _0529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1235_ _1491_/A _1235_/B _1235_/C vssd vssd vccd vccd _1236_/A sky130_fd_sc_hd__and3b_2
XFILLER_49_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1166_ _1166_/A vssd vssd vccd vccd _1166_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_2925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2947 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1097_ _1353_/A _1097_/B _1097_/C vssd vssd vccd vccd _1098_/A sky130_fd_sc_hd__and3b_2
XFILLER_52_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1079__B _1079_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0711__B _0711_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1261__C _1261_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input102_A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0902__A _0902_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0621__B _0621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_998 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1171__C _1171_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1020_ _1020_/A vssd vssd vccd vccd _1020_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output955_A _0874_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[13\] mprj_dat_i_user[13] _0870_/X vssd vssd vccd vccd _0589_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_28_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3906 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0804_ _0804_/A vssd vssd vccd vccd _0804_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__0812__A _0812_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0735_ _0735_/A _0735_/B vssd vssd vccd vccd _0736_/A sky130_fd_sc_hd__and2_1
XFILLER_45_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0666_ _0666_/A vssd vssd vccd vccd _0666_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0597_ _0597_/A vssd vssd vccd vccd _0597_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_wb_dat_gates\[1\]_A mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] _0830_/X vssd vssd vccd vccd _0556_/A
+ sky130_fd_sc_hd__nand2_1
X_1218_ _1218_/A vssd vssd vccd vccd _1218_/X sky130_fd_sc_hd__buf_4
XTAP_2909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1149_ _1405_/A _1149_/B _1149_/C vssd vssd vccd vccd _1150_/A sky130_fd_sc_hd__and3b_2
XFILLER_0_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1962 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput302 la_oenb_mprj[22] vssd vssd vccd vccd _1319_/A sky130_fd_sc_hd__buf_2
Xinput313 la_oenb_mprj[32] vssd vssd vccd vccd _1339_/A sky130_fd_sc_hd__clkbuf_2
Xinput324 la_oenb_mprj[42] vssd vssd vccd vccd _1359_/A sky130_fd_sc_hd__buf_2
XFILLER_0_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput335 la_oenb_mprj[52] vssd vssd vccd vccd _1379_/A sky130_fd_sc_hd__buf_2
XFILLER_40_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput346 la_oenb_mprj[62] vssd vssd vccd vccd _1399_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput357 la_oenb_mprj[72] vssd vssd vccd vccd _1419_/A sky130_fd_sc_hd__clkbuf_4
Xinput368 la_oenb_mprj[82] vssd vssd vccd vccd _1439_/A sky130_fd_sc_hd__buf_4
XFILLER_5_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput379 la_oenb_mprj[92] vssd vssd vccd vccd _1459_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input317_A la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_880 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1447__B _1447_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput809 _1408_/X vssd vssd vccd vccd la_oenb_core[66] sky130_fd_sc_hd__buf_12
XFILLER_46_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0520_ _0520_/A vssd vssd vccd vccd _0520_/Y sky130_fd_sc_hd__inv_2
XTAP_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output536_A _1120_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1463__A _1463_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output703_A _0531_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1003_ _1003_/A _1003_/B vssd vssd vccd vccd _1004_/A sky130_fd_sc_hd__and2_4
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] _0704_/X vssd vssd vccd vccd _0493_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__0807__A _0807_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0542__A _0542_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1357__B _1357_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0718_ _0718_/A vssd vssd vccd vccd _0718_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0649_ _0649_/A _0649_/B vssd vssd vccd vccd _0650_/A sky130_fd_sc_hd__and2_1
XANTENNA__1373__A _1373_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0717__A _0717_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1267__B _1267_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input267_A la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1283__A _1283_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input434_A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput110 la_data_out_mprj[80] vssd vssd vccd vccd _1179_/C sky130_fd_sc_hd__buf_4
Xinput121 la_data_out_mprj[90] vssd vssd vccd vccd _1199_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_41_3880 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input30_A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput132 la_iena_mprj[0] vssd vssd vccd vccd _1531_/B sky130_fd_sc_hd__clkbuf_1
Xinput143 la_iena_mprj[10] vssd vssd vccd vccd _0627_/B sky130_fd_sc_hd__buf_2
XFILLER_27_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput154 la_iena_mprj[11] vssd vssd vccd vccd _0629_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_2_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput165 la_iena_mprj[14] vssd vssd vccd vccd _0635_/B sky130_fd_sc_hd__clkbuf_1
Xinput176 la_iena_mprj[24] vssd vssd vccd vccd _0655_/B sky130_fd_sc_hd__clkbuf_1
Xinput187 la_iena_mprj[34] vssd vssd vccd vccd _0675_/B sky130_fd_sc_hd__clkbuf_1
Xinput198 la_iena_mprj[44] vssd vssd vccd vccd _0695_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0627__A _0627_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output486_A _1260_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1458__A _1458_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1035__A_N _1291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1177__B _1177_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput606 _0558_/Y vssd vssd vccd vccd la_data_in_mprj[113] sky130_fd_sc_hd__buf_12
Xoutput617 _0568_/Y vssd vssd vccd vccd la_data_in_mprj[123] sky130_fd_sc_hd__buf_12
Xoutput628 _0463_/Y vssd vssd vccd vccd la_data_in_mprj[18] sky130_fd_sc_hd__buf_12
Xoutput639 _0473_/Y vssd vssd vccd vccd la_data_in_mprj[28] sky130_fd_sc_hd__buf_12
XFILLER_29_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0503_ _0503_/A vssd vssd vccd vccd _0503_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output820_A _1428_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1185__A_N _1441_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1483_ _1483_/A _1483_/B vssd vssd vccd vccd _1484_/A sky130_fd_sc_hd__and2_1
XANTENNA_output918_A _0984_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2386 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0537__A _0537_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1368__A _1368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1087__B _1087_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3234 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1278__A _1278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input384_A la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input78_A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0910__A _0910_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0983_ _0983_/A _0983_/B vssd vssd vccd vccd _0984_/A sky130_fd_sc_hd__and2_2
XANTENNA_output868_A _0948_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1188__A _1188_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0820__A _0820_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput469 _1230_/X vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__buf_12
X_1535_ _1535_/A vssd vssd vccd vccd _1535_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1466_ _1466_/A vssd vssd vccd vccd _1466_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_1955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1397_ _1397_/A _1397_/B vssd vssd vccd vccd _1398_/A sky130_fd_sc_hd__and2_4
XFILLER_3_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1098__A _1098_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1139 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0730__A _0730_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input132_A la_iena_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0905__A _0905_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1455__B _1455_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2735 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1320_ _1320_/A vssd vssd vccd vccd _1320_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1251_ _1507_/A _1251_/B _1251_/C vssd vssd vccd vccd _1252_/A sky130_fd_sc_hd__and3b_1
XFILLER_42_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output616_A _0567_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1471__A _1471_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1223__A_N _1479_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1182_ _1182_/A vssd vssd vccd vccd _1182_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] _0668_/X vssd vssd vccd vccd _0475_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_33_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0815__A _0815_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0966_ _0966_/A vssd vssd vccd vccd _0966_/X sky130_fd_sc_hd__buf_6
XFILLER_31_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0897_ _0897_/A _0897_/B vssd vssd vccd vccd _0898_/A sky130_fd_sc_hd__and2_1
XFILLER_31_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0550__A _0550_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1365__B _1365_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1518_ _1518_/A vssd vssd vccd vccd _1518_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1449_ _1449_/A _1449_/B vssd vssd vccd vccd _1450_/A sky130_fd_sc_hd__and2_1
XFILLER_25_2289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1381__A _1381_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0709__B _0709_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_ack_gate_A mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0725__A _0725_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1259__C _1259_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1275__B _1275_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input347_A la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1291__A _1291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0619__B _0619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0635__A _0635_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0820_ _0820_/A vssd vssd vccd vccd _0820_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1169__C _1169_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0751_ _0751_/A _0751_/B vssd vssd vccd vccd _0752_/A sky130_fd_sc_hd__and2_2
XANTENNA_output566_A _1176_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0682_ _0682_/A vssd vssd vccd vccd _0682_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1185__B _1185_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output733_A _1500_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] _0764_/X vssd vssd vccd vccd _0523_/A
+ sky130_fd_sc_hd__nand2_8
X_1303_ _1303_/A _1303_/B vssd vssd vccd vccd _1304_/A sky130_fd_sc_hd__and2_2
XFILLER_22_2418 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1234_ _1234_/A vssd vssd vccd vccd _1234_/X sky130_fd_sc_hd__buf_2
XFILLER_4_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1165_ _1421_/A _1165_/B _1165_/C vssd vssd vccd vccd _1166_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1096_ _1096_/A vssd vssd vccd vccd _1096_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0545__A _0545_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1119__A_N _1375_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0949_ _0949_/A _0949_/B vssd vssd vccd vccd _0950_/A sky130_fd_sc_hd__and2_1
XANTENNA__1376__A _1376_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1269__A_N _1525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1839 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input297_A la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1286__A _1286_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input60_A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output850_A _0914_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0803_ _0803_/A _0803_/B vssd vssd vccd vccd _0804_/A sky130_fd_sc_hd__and2_4
XFILLER_11_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output948_A _0890_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1196__A _1196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0734_ _0734_/A vssd vssd vccd vccd _0734_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0665_ _0665_/A _0665_/B vssd vssd vccd vccd _0666_/A sky130_fd_sc_hd__and2_1
XFILLER_45_3686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0596_ _0596_/A vssd vssd vccd vccd _0596_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1217_ _1473_/A _1217_/B _1217_/C vssd vssd vccd vccd _1218_/A sky130_fd_sc_hd__and3b_1
XFILLER_39_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] _0816_/X vssd vssd vccd vccd _0549_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_26_826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1148_ _1148_/A vssd vssd vccd vccd _1148_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1079_ _1335_/A _1079_/B _1079_/C vssd vssd vccd vccd _1080_/A sky130_fd_sc_hd__and3b_2
XFILLER_33_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4066 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1996 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput303 la_oenb_mprj[23] vssd vssd vccd vccd _1321_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput314 la_oenb_mprj[33] vssd vssd vccd vccd _1341_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_2091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput325 la_oenb_mprj[43] vssd vssd vccd vccd _1361_/A sky130_fd_sc_hd__buf_6
Xinput336 la_oenb_mprj[53] vssd vssd vccd vccd _1381_/A sky130_fd_sc_hd__clkbuf_2
Xinput347 la_oenb_mprj[63] vssd vssd vccd vccd _1401_/A sky130_fd_sc_hd__buf_4
XFILLER_40_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput358 la_oenb_mprj[73] vssd vssd vccd vccd _1421_/A sky130_fd_sc_hd__clkbuf_4
Xinput369 la_oenb_mprj[83] vssd vssd vccd vccd _1441_/A sky130_fd_sc_hd__buf_4
XFILLER_28_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input212_A la_iena_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0913__A _0913_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1463__B _1463_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output529_A _1108_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1002_ _1002_/A vssd vssd vccd vccd _1002_/X sky130_fd_sc_hd__buf_6
XFILLER_53_3911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0823__A _0823_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0717_ _0717_/A _0717_/B vssd vssd vccd vccd _0718_/A sky130_fd_sc_hd__and2_1
XFILLER_41_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0648_ _0648_/A vssd vssd vccd vccd _0648_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1839 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1778 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0579_ _0579_/A vssd vssd vccd vccd _0579_/Y sky130_fd_sc_hd__inv_2
XTAP_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0717__B _0717_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1267__C _1267_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input162_A la_iena_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1283__B _1283_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput100 la_data_out_mprj[71] vssd vssd vccd vccd _1161_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput111 la_data_out_mprj[81] vssd vssd vccd vccd _1181_/C sky130_fd_sc_hd__buf_4
XFILLER_40_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput122 la_data_out_mprj[91] vssd vssd vccd vccd _1201_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_2_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput133 la_iena_mprj[100] vssd vssd vccd vccd _0807_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_41_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input427_A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput144 la_iena_mprj[110] vssd vssd vccd vccd _0827_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_2_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput155 la_iena_mprj[120] vssd vssd vccd vccd _0847_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput166 la_iena_mprj[15] vssd vssd vccd vccd _0637_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_input23_A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput177 la_iena_mprj[25] vssd vssd vccd vccd _0657_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput188 la_iena_mprj[35] vssd vssd vccd vccd _0677_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__0908__A _0908_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput199 la_iena_mprj[45] vssd vssd vccd vccd _0697_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0627__B _0627_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_656 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0643__A _0643_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output479_A _1248_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__1177__C _1177_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput607 _0559_/Y vssd vssd vccd vccd la_data_in_mprj[114] sky130_fd_sc_hd__buf_12
XFILLER_9_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput618 _0569_/Y vssd vssd vccd vccd la_data_in_mprj[124] sky130_fd_sc_hd__buf_12
Xoutput629 _0464_/Y vssd vssd vccd vccd la_data_in_mprj[19] sky130_fd_sc_hd__buf_12
XFILLER_25_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output646_A _0479_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1474__A _1474_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0502_ _0502_/A vssd vssd vccd vccd _0502_/Y sky130_fd_sc_hd__inv_2
X_1482_ _1482_/A vssd vssd vccd vccd _1482_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1193__B _1193_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] _0728_/X vssd vssd vccd vccd _0505_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_3_1703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0818__A _0818_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0553__A _0553_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_50_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1384__A _1384_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input377_A la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1294__A _1294_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output596_A _0549_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1469__A _1469_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0982_ _0982_/A vssd vssd vccd vccd _0982_/X sky130_fd_sc_hd__buf_6
XFILLER_35_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output930_A _1006_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1534_ _1534_/A vssd vssd vccd vccd _1534_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_3139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1923 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1465_ _1465_/A _1465_/B vssd vssd vccd vccd _1466_/A sky130_fd_sc_hd__and2_1
XFILLER_29_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1396_ _1396_/A vssd vssd vccd vccd _1396_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0548__A _0548_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3784 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1379__A _1379_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput960 _0872_/X vssd vssd vccd vccd user_reset sky130_fd_sc_hd__buf_12
XFILLER_28_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1025__A_N _1281_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input125_A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_968 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0905__B _0905_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1289__A _1289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1175__A_N _1431_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input90_A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0921__A _0921_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[6\] mprj_dat_i_user[6] _0870_/X vssd vssd vccd vccd _0582_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2747 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1250_ _1250_/A vssd vssd vccd vccd _1250_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_3266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1471__B _1471_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output511_A _1076_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1181_ _1437_/A _1181_/B _1181_/C vssd vssd vccd vccd _1182_/A sky130_fd_sc_hd__and3b_1
XANTENNA_output609_A _0561_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output880_A _0878_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__0815__B _0815_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] _0654_/X vssd vssd vccd vccd _0468_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_36_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0965_ _0965_/A _0965_/B vssd vssd vccd vccd _0966_/A sky130_fd_sc_hd__and2_1
XANTENNA__0831__A _0831_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0896_ _0896_/A vssd vssd vccd vccd _0896_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1517_ _1517_/A _1517_/B vssd vssd vccd vccd _1518_/A sky130_fd_sc_hd__and2_1
XFILLER_47_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1448_ _1448_/A vssd vssd vccd vccd _1448_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1381__B _1381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1379_ _1379_/A _1379_/B vssd vssd vccd vccd _1380_/A sky130_fd_sc_hd__and2_4
XFILLER_0_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0725__B _0725_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_45 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3058 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput790 _1374_/X vssd vssd vccd vccd la_oenb_core[49] sky130_fd_sc_hd__buf_12
XANTENNA_input242_A la_iena_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1291__B _1291_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0651__A _0651_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0750_ _0750_/A vssd vssd vccd vccd _0750_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0681_ _0681_/A _0681_/B vssd vssd vccd vccd _0682_/A sky130_fd_sc_hd__and2_2
XANTENNA_output559_A _1162_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1185__C _1185_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output726_A _1488_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1482__A _1482_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1302_ _1302_/A vssd vssd vccd vccd _1302_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1233_ _1489_/A _1233_/B _1233_/C vssd vssd vccd vccd _1234_/A sky130_fd_sc_hd__and3b_4
XFILLER_49_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1164_ _1164_/A vssd vssd vccd vccd _1164_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0826__A _0826_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1095_ _1351_/A _1095_/B _1095_/C vssd vssd vccd vccd _1096_/A sky130_fd_sc_hd__and3b_2
XFILLER_18_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_746 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0948_ _0948_/A vssd vssd vccd vccd _0948_/X sky130_fd_sc_hd__buf_4
XFILLER_44_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0879_ _0879_/A _0879_/B vssd vssd vccd vccd _0880_/A sky130_fd_sc_hd__and2_2
XFILLER_31_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1095__C _1095_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1392__A _1392_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4090 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input192_A la_iena_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1213__A_N _1469_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input457_A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input53_A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2831 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0646__A _0646_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1477__A _1477_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0802_ _0802_/A vssd vssd vccd vccd _0802_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0733_ _0733_/A _0733_/B vssd vssd vccd vccd _0734_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0664_ _0664_/A vssd vssd vccd vccd _0664_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] _0788_/X vssd vssd vccd vccd _0535_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_28_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0595_ _0595_/A vssd vssd vccd vccd _0595_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1216_ _1216_/A vssd vssd vccd vccd _1216_/X sky130_fd_sc_hd__buf_4
XFILLER_38_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1147_ _1403_/A _1147_/B _1147_/C vssd vssd vccd vccd _1148_/A sky130_fd_sc_hd__and3b_4
XFILLER_0_1322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1078_ _1078_/A vssd vssd vccd vccd _1078_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1387__A _1387_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput304 la_oenb_mprj[24] vssd vssd vccd vccd _1323_/A sky130_fd_sc_hd__clkbuf_2
Xinput315 la_oenb_mprj[34] vssd vssd vccd vccd _1343_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_44_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput326 la_oenb_mprj[44] vssd vssd vccd vccd _1363_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_2_3523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput337 la_oenb_mprj[54] vssd vssd vccd vccd _1383_/A sky130_fd_sc_hd__buf_6
XFILLER_29_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput348 la_oenb_mprj[64] vssd vssd vccd vccd _1403_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_2811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput359 la_oenb_mprj[74] vssd vssd vccd vccd _1423_/A sky130_fd_sc_hd__buf_4
XFILLER_40_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1036 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input205_A la_iena_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0913__B _0913_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1297__A _1297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_B _0718_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1109__A_N _1365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1001_ _1001_/A _1001_/B vssd vssd vccd vccd _1002_/A sky130_fd_sc_hd__and2_2
XFILLER_47_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1259__A_N _1515_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output793_A _1378_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output960_A _0872_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__0823__B _0823_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1000__A _1000_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0716_ _0716_/A vssd vssd vccd vccd _0716_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0647_ _0647_/A _0647_/B vssd vssd vccd vccd _0648_/A sky130_fd_sc_hd__and2_1
XFILLER_48_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0578_ _0578_/A vssd vssd vccd vccd _0578_/Y sky130_fd_sc_hd__inv_2
XTAP_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0733__B _0733_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input155_A la_iena_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput101 la_data_out_mprj[72] vssd vssd vccd vccd _1163_/C sky130_fd_sc_hd__buf_2
XFILLER_7_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput112 la_data_out_mprj[82] vssd vssd vccd vccd _1183_/C sky130_fd_sc_hd__buf_4
Xinput123 la_data_out_mprj[92] vssd vssd vccd vccd _1203_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput134 la_iena_mprj[101] vssd vssd vccd vccd _0809_/B sky130_fd_sc_hd__clkbuf_2
Xinput145 la_iena_mprj[111] vssd vssd vccd vccd _0829_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput156 la_iena_mprj[121] vssd vssd vccd vccd _0849_/B sky130_fd_sc_hd__buf_2
XFILLER_40_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input322_A la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput167 la_iena_mprj[16] vssd vssd vccd vccd _0639_/B sky130_fd_sc_hd__clkbuf_1
Xinput178 la_iena_mprj[26] vssd vssd vccd vccd _0659_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 la_iena_mprj[36] vssd vssd vccd vccd _0679_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[30\]_A mprj_dat_i_user[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0643__B _0643_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput608 _0560_/Y vssd vssd vccd vccd la_data_in_mprj[115] sky130_fd_sc_hd__buf_12
XFILLER_29_2723 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput619 _0570_/Y vssd vssd vccd vccd la_data_in_mprj[125] sky130_fd_sc_hd__buf_12
XFILLER_45_2002 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0501_ _0501_/A vssd vssd vccd vccd _0501_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1481_ _1481_/A _1481_/B vssd vssd vccd vccd _1482_/A sky130_fd_sc_hd__and2_1
XFILLER_46_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output639_A _0473_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1193__C _1193_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output806_A _1402_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] _0714_/X vssd vssd vccd vccd _0498_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_48_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_A mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0834__A _0834_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1414 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[103\]_B _0814_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input8_A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[12\]_A mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input272_A la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0919__A _0919_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1469__B _1469_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output491_A _1270_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0981_ _0981_/A _0981_/B vssd vssd vccd vccd _0982_/A sky130_fd_sc_hd__and2_4
XANTENNA_output589_A _1218_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output756_A _1312_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1485__A _1485_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1533_ _1533_/A vssd vssd vccd vccd _1533_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output923_A _0994_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2658 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1464_ _1464_/A vssd vssd vccd vccd _1464_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_1935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0829__A _0829_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1395_ _1395_/A _1395_/B vssd vssd vccd vccd _1396_/A sky130_fd_sc_hd__and2_4
XFILLER_7_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3763 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1379__B _1379_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1395__A _1395_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput950 _0882_/X vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__buf_12
XFILLER_47_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0474__A _0474_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1289__B _1289_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input83_A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0921__B _0921_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0649__A _0649_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1180_ _1180_/A vssd vssd vccd vccd _1180_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1199__B _1199_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output873_A _0898_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] _0640_/X vssd vssd vccd vccd _1549_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_18_2298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[29\] mprj_dat_i_user[29] _0870_/X vssd vssd vccd vccd _0605_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_31_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0964_ _0964_/A vssd vssd vccd vccd _0964_/X sky130_fd_sc_hd__buf_6
XFILLER_9_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0831__B _0831_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0895_ _0895_/A _0895_/B vssd vssd vccd vccd _0896_/A sky130_fd_sc_hd__and2_1
XFILLER_12_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1516_ _1516_/A vssd vssd vccd vccd _1516_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3919 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1447_ _1447_/A _1447_/B vssd vssd vccd vccd _1448_/A sky130_fd_sc_hd__and2_1
XFILLER_29_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] _0862_/X vssd vssd vccd vccd _0572_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_9_1787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1378_ _1378_/A vssd vssd vccd vccd _1378_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_3560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0741__B _0741_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput780 _1282_/X vssd vssd vccd vccd la_oenb_core[3] sky130_fd_sc_hd__buf_12
Xoutput791 _1284_/X vssd vssd vccd vccd la_oenb_core[4] sky130_fd_sc_hd__buf_12
XFILLER_47_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input235_A la_iena_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input402_A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0932__A _0932_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0651__B _0651_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0680_ _0680_/A vssd vssd vccd vccd _0680_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1301_ _1301_/A _1301_/B vssd vssd vccd vccd _1302_/A sky130_fd_sc_hd__and2_4
XANTENNA_output621_A _0572_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output719_A _1276_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1232_ _1232_/A vssd vssd vccd vccd _1232_/X sky130_fd_sc_hd__buf_2
XFILLER_38_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1163_ _1419_/A _1163_/B _1163_/C vssd vssd vccd vccd _1164_/A sky130_fd_sc_hd__and3b_1
XFILLER_37_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1094_ _1094_/A vssd vssd vccd vccd _1094_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1003__A _1003_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_758 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0947_ _0947_/A _0947_/B vssd vssd vccd vccd _0948_/A sky130_fd_sc_hd__and2_1
XFILLER_31_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0878_ _0878_/A vssd vssd vccd vccd _0878_/X sky130_fd_sc_hd__buf_6
XFILLER_44_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[4\]_A mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1165__A_N _1421_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0752__A _0752_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input185_A la_iena_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input352_A la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input46_A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3110 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2887 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0927__A _0927_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0662__A _0662_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1477__B _1477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3879 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0801_ _0801_/A _0801_/B vssd vssd vccd vccd _0802_/A sky130_fd_sc_hd__and2_4
XANTENNA_output571_A _1184_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0732_ _0732_/A vssd vssd vccd vccd _0732_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0663_ _0663_/A _0663_/B vssd vssd vccd vccd _0664_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1493__A _1493_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0594_ _0594_/A vssd vssd vccd vccd _0594_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] _0774_/X vssd vssd vccd vccd _0528_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1215_ _1471_/A _1215_/B _1215_/C vssd vssd vccd vccd _1216_/A sky130_fd_sc_hd__and3b_1
XFILLER_39_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0837__A _0837_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1146_ _1146_/A vssd vssd vccd vccd _1146_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1077_ _1333_/A _1077_/B _1077_/C vssd vssd vccd vccd _1078_/A sky130_fd_sc_hd__and3b_4
XFILLER_41_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1387__B _1387_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput305 la_oenb_mprj[25] vssd vssd vccd vccd _1325_/A sky130_fd_sc_hd__clkbuf_2
Xinput316 la_oenb_mprj[35] vssd vssd vccd vccd _1345_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput327 la_oenb_mprj[45] vssd vssd vccd vccd _1365_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput338 la_oenb_mprj[55] vssd vssd vccd vccd _1385_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput349 la_oenb_mprj[65] vssd vssd vccd vccd _1405_/A sky130_fd_sc_hd__buf_2
XFILLER_25_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0747__A _0747_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1048 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3234 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input100_A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1297__B _1297_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2695 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0657__A _0657_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1000_ _1000_/A vssd vssd vccd vccd _1000_/X sky130_fd_sc_hd__buf_6
XFILLER_1_3089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output786_A _1366_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output953_A output953/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[11\] mprj_dat_i_user[11] _0870_/X vssd vssd vccd vccd _0587_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_15_1375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0715_ _0715_/A _0715_/B vssd vssd vccd vccd _0716_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0646_ _0646_/A vssd vssd vccd vccd _0646_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0577_ _0577_/A vssd vssd vccd vccd _0577_/Y sky130_fd_sc_hd__clkinv_2
XTAP_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1203__A_N _1459_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1129_ _1385_/A _1129_/B _1129_/C vssd vssd vccd vccd _1130_/A sky130_fd_sc_hd__and3b_4
XFILLER_39_3289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1398__A _1398_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput102 la_data_out_mprj[73] vssd vssd vccd vccd _1165_/C sky130_fd_sc_hd__buf_2
XFILLER_0_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput113 la_data_out_mprj[83] vssd vssd vccd vccd _1185_/C sky130_fd_sc_hd__buf_4
XFILLER_7_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput124 la_data_out_mprj[93] vssd vssd vccd vccd _1205_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_0_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input148_A la_iena_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput135 la_iena_mprj[102] vssd vssd vccd vccd _0811_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput146 la_iena_mprj[112] vssd vssd vccd vccd _0831_/B sky130_fd_sc_hd__clkbuf_4
Xinput157 la_iena_mprj[122] vssd vssd vccd vccd _0851_/B sky130_fd_sc_hd__buf_2
Xinput168 la_iena_mprj[17] vssd vssd vccd vccd _0641_/B sky130_fd_sc_hd__clkbuf_1
XTAP_3900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0477__A _0477_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 la_iena_mprj[27] vssd vssd vccd vccd _0661_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_29_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input315_A la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[30\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0940__A _0940_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput609 _0561_/Y vssd vssd vccd vccd la_data_in_mprj[116] sky130_fd_sc_hd__buf_12
XFILLER_49_2161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0500_ _0500_/A vssd vssd vccd vccd _0500_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1480_ _1480_/A vssd vssd vccd vccd _1480_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output534_A _1118_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] _0700_/X vssd vssd vccd vccd _0491_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_47_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[21\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1011__A _1011_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] _0624_/X vssd vssd vccd vccd _1541_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_28_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0629_ _0629_/A _0629_/B vssd vssd vccd vccd _0630_/A sky130_fd_sc_hd__and2_1
XFILLER_41_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1880 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3616 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[12\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2672 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0760__A _0760_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input265_A la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1249__A_N _1505_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input432_A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0919__B _0919_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0935__A _0935_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0980_ _0980_/A vssd vssd vccd vccd _0980_/X sky130_fd_sc_hd__buf_6
XFILLER_31_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output484_A _1258_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0670__A _0670_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1485__B _1485_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output651_A _0484_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1532_ _1532_/A vssd vssd vccd vccd _1532_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output916_A _0980_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1463_ _1463_/A _1463_/B vssd vssd vccd vccd _1464_/A sky130_fd_sc_hd__and2_1
XFILLER_45_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1394_ _1394_/A vssd vssd vccd vccd _1394_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0829__B _0829_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1006__A _1006_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0845__A _0845_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1395__B _1395_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput940 _0966_/X vssd vssd vccd vccd mprj_dat_o_user[5] sky130_fd_sc_hd__buf_12
Xoutput951 output951/A vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_12
XFILLER_47_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1828 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0739__B _0739_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0755__A _0755_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input382_A la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1071__A_N _1327_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input76_A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0665__A _0665_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output866_A _0944_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0963_ _0963_/A _0963_/B vssd vssd vccd vccd _0964_/A sky130_fd_sc_hd__and2_1
XFILLER_31_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0894_ _0894_/A vssd vssd vccd vccd _0894_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1515_ _1515_/A _1515_/B vssd vssd vccd vccd _1516_/A sky130_fd_sc_hd__and2_1
XFILLER_9_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1755 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1446_ _1446_/A vssd vssd vccd vccd _1446_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_2011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1377_ _1377_/A _1377_/B vssd vssd vccd vccd _1378_/A sky130_fd_sc_hd__and2_1
XFILLER_28_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1919 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput770 _1336_/X vssd vssd vccd vccd la_oenb_core[30] sky130_fd_sc_hd__buf_12
Xoutput781 _1356_/X vssd vssd vccd vccd la_oenb_core[40] sky130_fd_sc_hd__buf_12
XFILLER_47_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput792 _1376_/X vssd vssd vccd vccd la_oenb_core[50] sky130_fd_sc_hd__buf_12
XFILLER_5_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input130_A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input228_A la_iena_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3822 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0485__A _0485_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1300_ _1300_/A vssd vssd vccd vccd _1300_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1231_ _1487_/A _1231_/B _1231_/C vssd vssd vccd vccd _1232_/A sky130_fd_sc_hd__and3b_4
XFILLER_4_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output614_A _0565_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1162_ _1162_/A vssd vssd vccd vccd _1162_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1093_ _1349_/A _1093_/B _1093_/C vssd vssd vccd vccd _1094_/A sky130_fd_sc_hd__and3b_1
XFILLER_52_317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1003__B _1003_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0946_ _0946_/A vssd vssd vccd vccd _0946_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_53_1297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0877_ _0877_/A _0877_/B vssd vssd vccd vccd _0878_/A sky130_fd_sc_hd__and2_1
XFILLER_44_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[4\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1429_ _1429_/A _1429_/B vssd vssd vccd vccd _1430_/A sky130_fd_sc_hd__and2_2
XFILLER_42_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_936 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input178_A la_iena_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input345_A la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3122 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input39_A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2432 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_314 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0927__B _0927_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1104__A _1104_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0800_ _0800_/A vssd vssd vccd vccd _0800_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0731_ _0731_/A _0731_/B vssd vssd vccd vccd _0732_/A sky130_fd_sc_hd__and2_1
XANTENNA_output564_A _1172_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0662_ _0662_/A vssd vssd vccd vccd _0662_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1493__B _1493_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output731_A _1496_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output829_A _1444_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0593_ _0593_/A vssd vssd vccd vccd _0593_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] _0760_/X vssd vssd vccd vccd _0521_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_23_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1214_ _1214_/A vssd vssd vccd vccd _1214_/X sky130_fd_sc_hd__buf_2
XFILLER_1_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0837__B _0837_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1145_ _1401_/A _1145_/B _1145_/C vssd vssd vccd vccd _1146_/A sky130_fd_sc_hd__and3b_4
XANTENNA__1014__A _1014_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1076_ _1076_/A vssd vssd vccd vccd _1076_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0853__A _0853_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0929_ _0929_/A _0929_/B vssd vssd vccd vccd _0930_/A sky130_fd_sc_hd__and2_1
XFILLER_11_1911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput306 la_oenb_mprj[26] vssd vssd vccd vccd _1327_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput317 la_oenb_mprj[36] vssd vssd vccd vccd _1347_/A sky130_fd_sc_hd__clkbuf_1
Xinput328 la_oenb_mprj[46] vssd vssd vccd vccd _1367_/A sky130_fd_sc_hd__buf_4
Xinput339 la_oenb_mprj[56] vssd vssd vccd vccd _1387_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0747__B _0747_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0763__A _0763_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1702 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_8_516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input295_A la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input462_A user_irq_ena[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0938__A _0938_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0657__B _0657_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0673__A _0673_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output779_A _1354_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1155__A_N _1411_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_37_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output946_A _0886_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0714_ _0714_/A vssd vssd vccd vccd _0714_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0645_ _0645_/A _0645_/B vssd vssd vccd vccd _0646_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1009__A _1009_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0576_ _0576_/A vssd vssd vccd vccd _0576_/Y sky130_fd_sc_hd__clkinv_2
XTAP_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] _0812_/X vssd vssd vccd vccd _0547_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1128_ _1128_/A vssd vssd vccd vccd _1128_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1059_ _1315_/A _1059_/B _1059_/C vssd vssd vccd vccd _1060_/A sky130_fd_sc_hd__and3b_2
XFILLER_41_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_16_1118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput103 la_data_out_mprj[74] vssd vssd vccd vccd _1167_/C sky130_fd_sc_hd__buf_4
Xinput114 la_data_out_mprj[84] vssd vssd vccd vccd _1187_/C sky130_fd_sc_hd__buf_4
XANTENNA__0758__A _0758_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput125 la_data_out_mprj[94] vssd vssd vccd vccd _1207_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput136 la_iena_mprj[103] vssd vssd vccd vccd _0813_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput147 la_iena_mprj[113] vssd vssd vccd vccd _0833_/B sky130_fd_sc_hd__clkbuf_4
Xinput158 la_iena_mprj[123] vssd vssd vccd vccd _0853_/B sky130_fd_sc_hd__buf_2
XFILLER_5_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput169 la_iena_mprj[18] vssd vssd vccd vccd _0643_/B sky130_fd_sc_hd__clkbuf_1
XTAP_3901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input210_A la_iena_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input308_A la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1101__B _1101_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1499__A _1499_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] _0686_/X vssd vssd vccd vccd _0484_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_36_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1011__B _1011_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2306 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0628_ _0628_/A vssd vssd vccd vccd _0628_/X sky130_fd_sc_hd__clkbuf_1
XTAP_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0559_ _0559_/A vssd vssd vccd vccd _0559_/Y sky130_fd_sc_hd__clkinv_4
XTAP_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1202__A _1202_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input160_A la_iena_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input258_A la_iena_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input425_A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input21_A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0935__B _0935_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1112__A _1112_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output477_A _1244_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1531_ _1531_/A _1531_/B vssd vssd vccd vccd _1532_/A sky130_fd_sc_hd__and2_1
XFILLER_29_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output644_A _0477_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1462_ _1462_/A vssd vssd vccd vccd _1462_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output909_A _0582_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1393_ _1393_/A _1393_/B vssd vssd vccd vccd _1394_/A sky130_fd_sc_hd__and2_1
XFILLER_20_3710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3798 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0845__B _0845_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1022__A _1022_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1847 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0861__A _0861_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput930 _1006_/X vssd vssd vccd vccd mprj_dat_o_user[25] sky130_fd_sc_hd__buf_12
Xoutput941 _0968_/X vssd vssd vccd vccd mprj_dat_o_user[6] sky130_fd_sc_hd__buf_12
XFILLER_9_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput952 output952/A vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_12
XFILLER_43_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0755__B _0755_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0771__A _0771_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2334 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input375_A la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input69_A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0665__B _0665_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3812 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0681__A _0681_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0962_ _0962_/A vssd vssd vccd vccd _0962_/X sky130_fd_sc_hd__buf_6
XFILLER_53_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output859_A _0894_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0893_ _0893_/A _0893_/B vssd vssd vccd vccd _0894_/A sky130_fd_sc_hd__and2_2
XFILLER_9_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3930 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1514_ _1514_/A vssd vssd vccd vccd _1514_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1445_ _1445_/A _1445_/B vssd vssd vccd vccd _1446_/A sky130_fd_sc_hd__and2_1
XFILLER_29_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1017__A _1017_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1376_ _1376_/A vssd vssd vccd vccd _1376_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1239__A_N _1495_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0591__A _0591_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1839 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput760 _1318_/X vssd vssd vccd vccd la_oenb_core[21] sky130_fd_sc_hd__buf_12
Xoutput771 _1338_/X vssd vssd vccd vccd la_oenb_core[31] sky130_fd_sc_hd__buf_12
XFILLER_40_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput782 _1358_/X vssd vssd vccd vccd la_oenb_core[41] sky130_fd_sc_hd__buf_12
XFILLER_8_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput793 _1378_/X vssd vssd vccd vccd la_oenb_core[51] sky130_fd_sc_hd__buf_12
XFILLER_47_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0766__A _0766_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input123_A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[4\] mprj_dat_i_user[4] _0870_/X vssd vssd vccd vccd _0580_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1230_ _1230_/A vssd vssd vccd vccd _1230_/X sky130_fd_sc_hd__buf_2
XFILLER_4_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0676__A _0676_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1161_ _1417_/A _1161_/B _1161_/C vssd vssd vccd vccd _1162_/A sky130_fd_sc_hd__and3b_1
XANTENNA_output607_A _0559_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1092_ _1092_/A vssd vssd vccd vccd _1092_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] _0650_/X vssd vssd vccd vccd _0466_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_37_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1300__A _1300_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0945_ _0945_/A _0945_/B vssd vssd vccd vccd _0946_/A sky130_fd_sc_hd__and2_1
XFILLER_31_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0876_ _0876_/A vssd vssd vccd vccd _0876_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1428_ _1428_/A vssd vssd vccd vccd _1428_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1359_ _1359_/A _1359_/B vssd vssd vccd vccd _1360_/A sky130_fd_sc_hd__and2_1
XFILLER_28_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1061__A_N _1317_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1210__A _1210_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput590 _1038_/X vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__buf_12
XFILLER_44_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input240_A la_iena_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input338_A la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0496__A _0496_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_2455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_863 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0943__B _0943_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1120__A _1120_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[58\]_B _0724_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0730_ _0730_/A vssd vssd vccd vccd _0730_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0661_ _0661_/A _0661_/B vssd vssd vccd vccd _0662_/A sky130_fd_sc_hd__and2_1
XANTENNA_output557_A _1032_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0592_ _0592_/A vssd vssd vccd vccd _0592_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_3911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output724_A _1484_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1213_ _1469_/A _1213_/B _1213_/C vssd vssd vccd vccd _1214_/A sky130_fd_sc_hd__and3b_4
XFILLER_38_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] _0746_/X vssd vssd vccd vccd _0514_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_39_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1144_ _1144_/A vssd vssd vccd vccd _1144_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_3795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1075_ _1331_/A _1075_/B _1075_/C vssd vssd vccd vccd _1076_/A sky130_fd_sc_hd__and3b_1
XFILLER_20_1275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0853__B _0853_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0928_ _0928_/A vssd vssd vccd vccd _0928_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0859_ _0859_/A _0859_/B vssd vssd vccd vccd _0860_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput307 la_oenb_mprj[27] vssd vssd vccd vccd _1329_/A sky130_fd_sc_hd__buf_2
XFILLER_6_3673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput318 la_oenb_mprj[37] vssd vssd vccd vccd _1349_/A sky130_fd_sc_hd__buf_4
Xinput329 la_oenb_mprj[47] vssd vssd vccd vccd _1369_/A sky130_fd_sc_hd__buf_6
XFILLER_40_2319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_863 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0763__B _0763_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1714 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input190_A la_iena_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input288_A la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input455_A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input51_A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0673__B _0673_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0713_ _0713_/A _0713_/B vssd vssd vccd vccd _0714_/A sky130_fd_sc_hd__and2_1
XANTENNA_output841_A _1466_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output939_A _0964_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0644_ _0644_/A vssd vssd vccd vccd _0644_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1009__B _1009_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0575_ _0575_/A vssd vssd vccd vccd _0575_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[24\]_A mprj_dat_i_user[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1127_ _1383_/A _1127_/B _1127_/C vssd vssd vccd vccd _1128_/A sky130_fd_sc_hd__and3b_4
XFILLER_17_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1058_ _1058_/A vssd vssd vccd vccd _1058_/X sky130_fd_sc_hd__buf_4
XFILLER_0_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput104 la_data_out_mprj[75] vssd vssd vccd vccd _1169_/C sky130_fd_sc_hd__buf_2
XFILLER_4_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput115 la_data_out_mprj[85] vssd vssd vccd vccd _1189_/C sky130_fd_sc_hd__buf_4
XFILLER_41_3874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput126 la_data_out_mprj[95] vssd vssd vccd vccd _1209_/C sky130_fd_sc_hd__clkbuf_1
Xinput137 la_iena_mprj[104] vssd vssd vccd vccd _0815_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_3345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput148 la_iena_mprj[114] vssd vssd vccd vccd _0835_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput159 la_iena_mprj[124] vssd vssd vccd vccd _0855_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_40_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[15\]_A mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0774__A _0774_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input203_A la_iena_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1101__C _1101_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input99_A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1499__B _1499_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output791_A _1284_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3898 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0627_ _0627_/A _0627_/B vssd vssd vccd vccd _0628_/A sky130_fd_sc_hd__and2_1
XFILLER_5_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0859__A _0859_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0558_ _0558_/A vssd vssd vccd vccd _0558_/Y sky130_fd_sc_hd__inv_4
XFILLER_6_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0489_ _0489_/A vssd vssd vccd vccd _0489_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_41_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0594__A _0594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3542 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0769__A _0769_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input153_A la_iena_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_2509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1145__A_N _1401_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input320_A la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input418_A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0951__B _0951_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1530_ _1530_/A vssd vssd vccd vccd _1530_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0679__A _0679_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1461_ _1461_/A _1461_/B vssd vssd vccd vccd _1462_/A sky130_fd_sc_hd__and2_1
XFILLER_46_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output637_A _0471_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1392_ _1392_/A vssd vssd vccd vccd _1392_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] _0710_/X vssd vssd vccd vccd _0496_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_40_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1303__A _1303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1859 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput920 _0988_/X vssd vssd vccd vccd mprj_dat_o_user[16] sky130_fd_sc_hd__buf_12
XFILLER_2_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput931 _1008_/X vssd vssd vccd vccd mprj_dat_o_user[26] sky130_fd_sc_hd__buf_12
Xoutput942 _0970_/X vssd vssd vccd vccd mprj_dat_o_user[7] sky130_fd_sc_hd__buf_12
Xoutput953 output953/A vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_12
XFILLER_45_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input6_A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2346 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input270_A la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4030 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input368_A la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0499__A _0499_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1107__B _1107_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3824 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0681__B _0681_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0961_ _0961_/A _0961_/B vssd vssd vccd vccd _0962_/A sky130_fd_sc_hd__and2_1
XANTENNA_output587_A _1214_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0892_ _0892_/A vssd vssd vccd vccd _0892_/X sky130_fd_sc_hd__buf_2
XFILLER_48_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output921_A _0990_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1513_ _1513_/A _1513_/B vssd vssd vccd vccd _1514_/A sky130_fd_sc_hd__and2_1
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] _0806_/X vssd vssd vccd vccd _0544_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_29_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3942 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1444_ _1444_/A vssd vssd vccd vccd _1444_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_3828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1017__B _1017_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1375_ _1375_/A _1375_/B vssd vssd vccd vccd _1376_/A sky130_fd_sc_hd__and2_4
XFILLER_0_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[7\]_A mprj_dat_i_user[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput750 _1300_/X vssd vssd vccd vccd la_oenb_core[12] sky130_fd_sc_hd__buf_12
XANTENNA__1208__A _1208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput761 _1320_/X vssd vssd vccd vccd la_oenb_core[22] sky130_fd_sc_hd__buf_12
Xoutput772 _1340_/X vssd vssd vccd vccd la_oenb_core[32] sky130_fd_sc_hd__buf_12
Xoutput783 _1360_/X vssd vssd vccd vccd la_oenb_core[42] sky130_fd_sc_hd__buf_12
XFILLER_5_3535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput794 _1380_/X vssd vssd vccd vccd la_oenb_core[52] sky130_fd_sc_hd__buf_12
XFILLER_5_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0782__A _0782_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input81_A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1118__A _1118_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1160_ _1160_/A vssd vssd vccd vccd _1160_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output502_A _1022_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1091_ _1347_/A _1091_/B _1091_/C vssd vssd vccd vccd _1092_/A sky130_fd_sc_hd__and3b_2
XTAP_4082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output871_A _0952_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[27\] mprj_dat_i_user[27] _0870_/X vssd vssd vccd vccd _0603_/A
+ sky130_fd_sc_hd__nand2_1
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] _0636_/X vssd vssd vccd vccd _1547_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_18_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0944_ _0944_/A vssd vssd vccd vccd _0944_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0875_ _0875_/A input2/X vssd vssd vccd vccd _0876_/A sky130_fd_sc_hd__and2_1
XFILLER_44_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1427_ _1427_/A _1427_/B vssd vssd vccd vccd _1428_/A sky130_fd_sc_hd__and2_1
XANTENNA__0867__A _0867_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] _0858_/X vssd vssd vccd vccd _0570_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_9_1587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1358_ _1358_/A vssd vssd vccd vccd _1358_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_3371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1289_ _1289_/A _1289_/B vssd vssd vccd vccd _1290_/A sky130_fd_sc_hd__and2_4
XFILLER_23_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput580 _1200_/X vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__buf_12
XFILLER_40_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput591 _1533_/Y vssd vssd vccd vccd la_data_in_mprj[0] sky130_fd_sc_hd__buf_12
XFILLER_43_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0777__A _0777_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input233_A la_iena_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input400_A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3930 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3086 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1401__A _1401_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0660_ _0660_/A vssd vssd vccd vccd _0660_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0591_ _0591_/A vssd vssd vccd vccd _0591_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1229__A_N _1485_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0687__A _0687_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1212_ _1212_/A vssd vssd vccd vccd _1212_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_38_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1143_ _1399_/A _1143_/B _1143_/C vssd vssd vccd vccd _1144_/A sky130_fd_sc_hd__and3b_4
XFILLER_38_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1074_ _1074_/A vssd vssd vccd vccd _1074_/X sky130_fd_sc_hd__buf_4
XFILLER_19_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1311__A _1311_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0927_ _0927_/A _0927_/B vssd vssd vccd vccd _0928_/A sky130_fd_sc_hd__and2_1
XFILLER_31_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0858_ _0858_/A vssd vssd vccd vccd _0858_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0789_ _0789_/A _0789_/B vssd vssd vccd vccd _0790_/A sky130_fd_sc_hd__and2_4
XFILLER_28_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput308 la_oenb_mprj[28] vssd vssd vccd vccd _1331_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput319 la_oenb_mprj[38] vssd vssd vccd vccd _1351_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_3685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1205__B _1205_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input183_A la_iena_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input350_A la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input448_A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input44_A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1115__B _1115_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0970__A _0970_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output667_A _0498_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0712_ _0712_/A vssd vssd vccd vccd _0712_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1051__A_N _1307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0643_ _0643_/A _0643_/B vssd vssd vccd vccd _0644_/A sky130_fd_sc_hd__and2_1
XFILLER_10_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0574_ _0574_/A vssd vssd vccd vccd _0574_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] _0770_/X vssd vssd vccd vccd _0526_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1306__A _1306_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1025__B _1025_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[24\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1126_ _1126_/A vssd vssd vccd vccd _1126_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1057_ _1313_/A _1057_/B _1057_/C vssd vssd vccd vccd _1058_/A sky130_fd_sc_hd__and3b_1
XFILLER_15_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3270 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0880__A _0880_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput105 la_data_out_mprj[76] vssd vssd vccd vccd _1171_/C sky130_fd_sc_hd__buf_4
Xinput116 la_data_out_mprj[86] vssd vssd vccd vccd _1191_/C sky130_fd_sc_hd__buf_4
XFILLER_44_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput127 la_data_out_mprj[96] vssd vssd vccd vccd _1211_/C sky130_fd_sc_hd__clkbuf_1
Xinput138 la_iena_mprj[105] vssd vssd vccd vccd _0817_/B sky130_fd_sc_hd__clkbuf_1
Xinput149 la_iena_mprj[115] vssd vssd vccd vccd _0837_/B sky130_fd_sc_hd__buf_4
XFILLER_22_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[15\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_466 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0790__A _0790_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input398_A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_576 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0949__B _0949_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1126__A _1126_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0965__A _0965_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_A user_irq_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output951_A output951/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0626_ _0626_/A vssd vssd vccd vccd _0626_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0859__B _0859_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0557_ _0557_/A vssd vssd vccd vccd _0557_/Y sky130_fd_sc_hd__clkinv_4
XTAP_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1036__A _1036_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0488_ _0488_/A vssd vssd vccd vccd _0488_/Y sky130_fd_sc_hd__clkinv_2
XTAP_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0875__A _0875_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1109_ _1365_/A _1109_/B _1109_/C vssd vssd vccd vccd _1110_/A sky130_fd_sc_hd__and3b_2
XFILLER_26_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input146_A la_iena_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0785__A _0785_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input313_A la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3730 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1460_ _1460_/A vssd vssd vccd vccd _1460_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0679__B _0679_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1391_ _1391_/A _1391_/B vssd vssd vccd vccd _1392_/A sky130_fd_sc_hd__and2_4
XFILLER_7_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3986 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0695__A _0695_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1303__B _1303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] _0696_/X vssd vssd vccd vccd _0489_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_1_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput910 _0583_/Y vssd vssd vccd vccd mprj_dat_i_core[7] sky130_fd_sc_hd__buf_12
XFILLER_28_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput921 _0990_/X vssd vssd vccd vccd mprj_dat_o_user[17] sky130_fd_sc_hd__buf_12
Xoutput932 _1010_/X vssd vssd vccd vccd mprj_dat_o_user[27] sky130_fd_sc_hd__buf_12
Xoutput943 _0972_/X vssd vssd vccd vccd mprj_dat_o_user[8] sky130_fd_sc_hd__buf_12
XFILLER_47_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] _0620_/X vssd vssd vccd vccd _1539_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_25_2900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput954 output954/A vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_12
XFILLER_45_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0609_ _0609_/A _0609_/B vssd vssd vccd vccd _0610_/A sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1213__B _1213_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input263_A la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input430_A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1107__C _1107_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1404__A _1404_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1123__B _1123_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0960_ _0960_/A vssd vssd vccd vccd _0960_/X sky130_fd_sc_hd__buf_6
XFILLER_53_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output482_A _1254_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0891_ _0891_/A _0891_/B vssd vssd vccd vccd _0892_/A sky130_fd_sc_hd__and2_1
XFILLER_51_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1512_ _1512_/A vssd vssd vccd vccd _1512_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output914_A _0976_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1443_ _1443_/A _1443_/B vssd vssd vccd vccd _1444_/A sky130_fd_sc_hd__and2_2
XFILLER_42_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1374_ _1374_/A vssd vssd vccd vccd _1374_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1314__A _1314_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1033__B _1033_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_954 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1135__A_N _1391_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[7\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput740 _1514_/X vssd vssd vccd vccd la_oenb_core[119] sky130_fd_sc_hd__buf_12
Xoutput751 _1302_/X vssd vssd vccd vccd la_oenb_core[13] sky130_fd_sc_hd__buf_12
XFILLER_47_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput762 _1322_/X vssd vssd vccd vccd la_oenb_core[23] sky130_fd_sc_hd__buf_12
Xoutput773 _1342_/X vssd vssd vccd vccd la_oenb_core[33] sky130_fd_sc_hd__buf_12
XFILLER_9_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput784 _1362_/X vssd vssd vccd vccd la_oenb_core[43] sky130_fd_sc_hd__buf_12
XFILLER_25_2730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput795 _1382_/X vssd vssd vccd vccd la_oenb_core[53] sky130_fd_sc_hd__buf_12
XFILLER_5_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1224__A _1224_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2534 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input109_A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input380_A la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input74_A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0957__B _0957_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1134__A _1134_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1090_ _1090_/A vssd vssd vccd vccd _1090_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0973__A _0973_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0943_ _0943_/A _0943_/B vssd vssd vccd vccd _0944_/A sky130_fd_sc_hd__and2_1
XANTENNA_output864_A _0940_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3390 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0874_ _0874_/A vssd vssd vccd vccd _0874_/X sky130_fd_sc_hd__buf_6
XFILLER_31_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1309__A _1309_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1426_ _1426_/A vssd vssd vccd vccd _1426_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0867__B _0867_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1357_ _1357_/A _1357_/B vssd vssd vccd vccd _1358_/A sky130_fd_sc_hd__and2_4
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] _0844_/X vssd vssd vccd vccd _0563_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_3_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1288_ _1288_/A vssd vssd vccd vccd _1288_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__0883__A _0883_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput570 _1182_/X vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__buf_12
XFILLER_44_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput581 _1202_/X vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__buf_12
XFILLER_47_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput592 _0545_/Y vssd vssd vccd vccd la_data_in_mprj[100] sky130_fd_sc_hd__buf_12
XFILLER_5_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input226_A la_iena_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0793__A _0793_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XTAP_1243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1401__B _1401_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1863 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1251 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3604 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0590_ _0590_/A vssd vssd vccd vccd _0590_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1211_ _1467_/A _1211_/B _1211_/C vssd vssd vccd vccd _1212_/A sky130_fd_sc_hd__and3b_4
XFILLER_46_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output612_A _0564_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1142_ _1142_/A vssd vssd vccd vccd _1142_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1073_ _1329_/A _1073_/B _1073_/C vssd vssd vccd vccd _1074_/A sky130_fd_sc_hd__and3b_1
XFILLER_52_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__1311__B _1311_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0926_ _0926_/A vssd vssd vccd vccd _0926_/X sky130_fd_sc_hd__buf_6
XFILLER_31_2052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1974 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0857_ _0857_/A _0857_/B vssd vssd vccd vccd _0858_/A sky130_fd_sc_hd__and2_1
XFILLER_11_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0788_ _0788_/A vssd vssd vccd vccd _0788_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput309 la_oenb_mprj[29] vssd vssd vccd vccd _1333_/A sky130_fd_sc_hd__buf_4
XFILLER_29_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1409_ _1409_/A _1409_/B vssd vssd vccd vccd _1410_/A sky130_fd_sc_hd__and2_1
XFILLER_26_2891 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__1221__B _1221_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input176_A la_iena_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0788__A _0788_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input343_A la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input37_A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1115__C _1115_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1412__A _1412_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1131__B _1131_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0711_ _0711_/A _0711_/B vssd vssd vccd vccd _0712_/A sky130_fd_sc_hd__and2_1
XANTENNA_output562_A _1168_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0642_ _0642_/A vssd vssd vccd vccd _0642_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0698__A _0698_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output827_A _1440_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0573_ _0573_/A vssd vssd vccd vccd _0573_/Y sky130_fd_sc_hd__inv_2
XTAP_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] _0756_/X vssd vssd vccd vccd _0519_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1025__C _1025_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1125_ _1381_/A _1125_/B _1125_/C vssd vssd vccd vccd _1126_/A sky130_fd_sc_hd__and3b_4
XFILLER_38_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1322__A _1322_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1056_ _1056_/A vssd vssd vccd vccd _1056_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1041__B _1041_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0909_ _0909_/A _0909_/B vssd vssd vccd vccd _0910_/A sky130_fd_sc_hd__and2_1
XFILLER_50_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput106 la_data_out_mprj[77] vssd vssd vccd vccd _1173_/C sky130_fd_sc_hd__buf_4
XFILLER_41_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput117 la_data_out_mprj[87] vssd vssd vccd vccd _1193_/C sky130_fd_sc_hd__buf_6
XFILLER_2_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput128 la_data_out_mprj[97] vssd vssd vccd vccd _1213_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_48_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput139 la_iena_mprj[106] vssd vssd vccd vccd _0819_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_478 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1232__A _1232_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1219__A_N _1475_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input293_A la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input460_A user_irq_ena[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_94 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1407__A _1407_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0965__B _0965_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1142__A _1142_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_990 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0981__A _0981_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output944_A _0974_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0625_ _0625_/A _0625_/B vssd vssd vccd vccd _0626_/A sky130_fd_sc_hd__and2_1
XFILLER_25_3827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1317__A _1317_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0556_ _0556_/A vssd vssd vccd vccd _0556_/Y sky130_fd_sc_hd__inv_4
XFILLER_3_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0487_ _0487_/A vssd vssd vccd vccd _0487_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] _0808_/X vssd vssd vccd vccd _0545_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_3_2999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1052__A _1052_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2334 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1108_ _1108_/A vssd vssd vccd vccd _1108_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0891__A _0891_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1039_ _1295_/A _1039_/B _1039_/C vssd vssd vccd vccd _1040_/A sky130_fd_sc_hd__and3b_4
XFILLER_17_2621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input139_A la_iena_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1041__A_N _1297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input306_A la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1191__A_N _1447_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1390_ _1390_/A vssd vssd vccd vccd _1390_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0976__A _0976_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output525_A _1100_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0695__B _0695_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] _0682_/X vssd vssd vccd vccd _0482_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_36_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput900 _0603_/Y vssd vssd vccd vccd mprj_dat_i_core[27] sky130_fd_sc_hd__buf_12
XFILLER_47_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput911 _0584_/Y vssd vssd vccd vccd mprj_dat_i_core[8] sky130_fd_sc_hd__buf_12
XFILLER_9_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput922 _0992_/X vssd vssd vccd vccd mprj_dat_o_user[18] sky130_fd_sc_hd__buf_12
Xoutput933 _1012_/X vssd vssd vccd vccd mprj_dat_o_user[28] sky130_fd_sc_hd__buf_12
Xoutput944 _0974_/X vssd vssd vccd vccd mprj_dat_o_user[9] sky130_fd_sc_hd__buf_12
XFILLER_8_2107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput955 _0874_/X vssd vssd vccd vccd user_clock sky130_fd_sc_hd__buf_12
XFILLER_47_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0608_ _0608_/A vssd vssd vccd vccd _0608_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_28_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0886__A _0886_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ _0539_/A vssd vssd vccd vccd _0539_/Y sky130_fd_sc_hd__inv_2
XTAP_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1510__A _1510_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3959 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_4054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3882 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input256_A la_iena_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0796__A _0796_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input423_A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1123__C _1123_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[88\]_B _0784_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1420__A _1420_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0890_ _0890_/A vssd vssd vccd vccd _0890_/X sky130_fd_sc_hd__buf_8
XFILLER_48_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output475_A _1240_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1511_ _1511_/A _1511_/B vssd vssd vccd vccd _1512_/A sky130_fd_sc_hd__and2_1
XFILLER_29_3067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output642_A _0475_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1442_ _1442_/A vssd vssd vccd vccd _1442_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[12\]_B _0632_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1373_ _1373_/A _1373_/B vssd vssd vccd vccd _1374_/A sky130_fd_sc_hd__and2_1
XFILLER_42_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output907_A _0580_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1033__C _1033_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1330__A _1330_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1046 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_966 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput730 _1296_/X vssd vssd vccd vccd la_oenb_core[10] sky130_fd_sc_hd__buf_12
Xoutput741 _1298_/X vssd vssd vccd vccd la_oenb_core[11] sky130_fd_sc_hd__buf_12
Xoutput752 _1304_/X vssd vssd vccd vccd la_oenb_core[14] sky130_fd_sc_hd__buf_12
XFILLER_47_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput763 _1324_/X vssd vssd vccd vccd la_oenb_core[24] sky130_fd_sc_hd__buf_12
Xoutput774 _1344_/X vssd vssd vccd vccd la_oenb_core[34] sky130_fd_sc_hd__buf_12
Xoutput785 _1364_/X vssd vssd vccd vccd la_oenb_core[44] sky130_fd_sc_hd__buf_12
XFILLER_25_3465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput796 _1384_/X vssd vssd vccd vccd la_oenb_core[54] sky130_fd_sc_hd__buf_12
XFILLER_25_3487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1505__A _1505_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1240__A _1240_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input373_A la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input67_A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1415__A _1415_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0973__B _0973_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1150__A _1150_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0942_ _0942_/A vssd vssd vccd vccd _0942_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output857_A _0928_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0873_ _0873_/A input1/X vssd vssd vccd vccd _0874_/A sky130_fd_sc_hd__and2_2
XFILLER_31_1544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1309__B _1309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1425_ _1425_/A _1425_/B vssd vssd vccd vccd _1426_/A sky130_fd_sc_hd__and2_1
XFILLER_6_3879 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1325__A _1325_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1356_ _1356_/A vssd vssd vccd vccd _1356_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1287_ _1287_/A _1287_/B vssd vssd vccd vccd _1288_/A sky130_fd_sc_hd__and2_4
XFILLER_37_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1060__A _1060_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1219__B _1219_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput560 _1164_/X vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__buf_12
XFILLER_5_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput571 _1184_/X vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__buf_12
XFILLER_43_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput582 _1204_/X vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__buf_12
XFILLER_44_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput593 _0546_/Y vssd vssd vccd vccd la_data_in_mprj[101] sky130_fd_sc_hd__buf_12
XFILLER_8_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input121_A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input219_A la_iena_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[2\] mprj_dat_i_user[2] _0870_/X vssd vssd vccd vccd _0578_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3616 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1129__B _1129_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1210_ _1210_/A vssd vssd vccd vccd _1210_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_3743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1125__A_N _1381_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1141_ _1397_/A _1141_/B _1141_/C vssd vssd vccd vccd _1142_/A sky130_fd_sc_hd__and3b_4
XANTENNA_output605_A _0557_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__0984__A _0984_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2198 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1072_ _1072_/A vssd vssd vccd vccd _1072_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0925_ _0925_/A _0925_/B vssd vssd vccd vccd _0926_/A sky130_fd_sc_hd__and2_1
XFILLER_11_2627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0856_ _0856_/A vssd vssd vccd vccd _0856_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1039__B _1039_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0787_ _0787_/A _0787_/B vssd vssd vccd vccd _0788_/A sky130_fd_sc_hd__and2_4
XFILLER_48_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1270 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[27\]_A mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1408_ _1408_/A vssd vssd vccd vccd _1408_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0894__A _0894_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1339_ _1339_/A _1339_/B vssd vssd vccd vccd _1340_/A sky130_fd_sc_hd__and2_2
XFILLER_25_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input169_A la_iena_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[18\]_A mprj_dat_i_user[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input336_A la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1131__C _1131_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0710_ _0710_/A vssd vssd vccd vccd _0710_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0641_ _0641_/A _0641_/B vssd vssd vccd vccd _0642_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0979__A _0979_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output555_A _1156_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0572_ _0572_/A vssd vssd vccd vccd _0572_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output722_A _1480_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] _0742_/X vssd vssd vccd vccd _0512_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_39_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1124_ _1124_/A vssd vssd vccd vccd _1124_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_3595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1055_ _1311_/A _1055_/B _1055_/C vssd vssd vccd vccd _1056_/A sky130_fd_sc_hd__and3b_4
XFILLER_53_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1041__C _1041_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0908_ _0908_/A vssd vssd vccd vccd _0908_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0889__A _0889_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0839_ _0839_/A _0839_/B vssd vssd vccd vccd _0840_/A sky130_fd_sc_hd__and2_2
XFILLER_8_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput107 la_data_out_mprj[78] vssd vssd vccd vccd _1175_/C sky130_fd_sc_hd__buf_4
XFILLER_22_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput118 la_data_out_mprj[88] vssd vssd vccd vccd _1195_/C sky130_fd_sc_hd__buf_2
XFILLER_2_3326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput129 la_data_out_mprj[98] vssd vssd vccd vccd _1215_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1513__A _1513_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input286_A la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0799__A _0799_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_73 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input453_A mprj_iena_wb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1407__B _1407_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1423__A _1423_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0981__B _0981_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output937_A _1018_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0502__A _0502_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0624_ _0624_/A vssd vssd vccd vccd _0624_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_3839 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1317__B _1317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0555_ _0555_/A vssd vssd vccd vccd _0555_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_28_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0486_ _0486_/A vssd vssd vccd vccd _0486_/Y sky130_fd_sc_hd__clkinv_2
XTAP_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1333__A _1333_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1107_ _1363_/A _1107_/B _1107_/C vssd vssd vccd vccd _1108_/A sky130_fd_sc_hd__and3b_2
XFILLER_39_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0891__B _0891_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1038_ _1038_/A vssd vssd vccd vccd _1038_/X sky130_fd_sc_hd__buf_2
XFILLER_17_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3990 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1227__B _1227_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2074 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input201_A la_iena_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input97_A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1418__A _1418_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1137__B _1137_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3922 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output518_A _1088_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput460 user_irq_ena[0] vssd vssd vccd vccd _0863_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_40_3195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0992__A _0992_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3632 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output887_A _0591_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1328__A _1328_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput901 _0604_/Y vssd vssd vccd vccd mprj_dat_i_core[28] sky130_fd_sc_hd__buf_12
Xoutput912 _0585_/Y vssd vssd vccd vccd mprj_dat_i_core[9] sky130_fd_sc_hd__buf_12
Xoutput923 _0994_/X vssd vssd vccd vccd mprj_dat_o_user[19] sky130_fd_sc_hd__buf_12
XFILLER_9_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput934 _1014_/X vssd vssd vccd vccd mprj_dat_o_user[29] sky130_fd_sc_hd__buf_12
XFILLER_47_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput945 _0884_/X vssd vssd vccd vccd mprj_sel_o_user[0] sky130_fd_sc_hd__buf_12
Xoutput956 _0876_/X vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__buf_12
XFILLER_8_2119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1047__B _1047_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0607_ _0607_/A vssd vssd vccd vccd _0607_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1209__A_N _1465_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0538_ _0538_/A vssd vssd vccd vccd _0538_/Y sky130_fd_sc_hd__inv_2
XTAP_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0469_ _0469_/A vssd vssd vccd vccd _0469_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_39_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3142 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_783 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1238__A _1238_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4066 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3894 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input151_A la_iena_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input249_A la_iena_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input416_A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output468_A _1228_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1148__A _1148_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1510_ _1510_/A vssd vssd vccd vccd _1510_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0987__A _0987_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1441_ _1441_/A _1441_/B vssd vssd vccd vccd _1442_/A sky130_fd_sc_hd__and2_1
XFILLER_26_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output635_A _0469_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1372_ _1372_/A vssd vssd vccd vccd _1372_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output802_A _1286_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput290 la_oenb_mprj[127] vssd vssd vccd vccd _1529_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1031__A_N _1287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput720 _1476_/X vssd vssd vccd vccd la_oenb_core[100] sky130_fd_sc_hd__buf_12
XFILLER_47_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput731 _1496_/X vssd vssd vccd vccd la_oenb_core[110] sky130_fd_sc_hd__buf_12
XFILLER_9_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput742 _1516_/X vssd vssd vccd vccd la_oenb_core[120] sky130_fd_sc_hd__buf_12
Xoutput753 _1306_/X vssd vssd vccd vccd la_oenb_core[15] sky130_fd_sc_hd__buf_12
XANTENNA__0897__A _0897_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput764 _1326_/X vssd vssd vccd vccd la_oenb_core[25] sky130_fd_sc_hd__buf_12
XFILLER_47_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput775 _1346_/X vssd vssd vccd vccd la_oenb_core[35] sky130_fd_sc_hd__buf_12
XFILLER_5_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput786 _1366_/X vssd vssd vccd vccd la_oenb_core[45] sky130_fd_sc_hd__buf_12
XFILLER_5_3538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput797 _1386_/X vssd vssd vccd vccd la_oenb_core[55] sky130_fd_sc_hd__buf_12
XFILLER_21_3308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1505__B _1505_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1181__A_N _1437_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1521__A _1521_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input199_A la_iena_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input366_A la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_irq_gates\[1\] user_irq_core[1] _0866_/X vssd vssd vccd vccd _0574_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1415__B _1415_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1431__A _1431_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0941_ _0941_/A _0941_/B vssd vssd vccd vccd _0942_/A sky130_fd_sc_hd__and2_1
XANTENNA_output585_A _1210_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0872_ _0872_/A vssd vssd vccd vccd _0872_/X sky130_fd_sc_hd__buf_2
XFILLER_35_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] _0802_/X vssd vssd vccd vccd _0542_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_42_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0510__A _0510_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1424_ _1424_/A vssd vssd vccd vccd _1424_/X sky130_fd_sc_hd__buf_2
XFILLER_25_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1325__B _1325_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1355_ _1355_/A _1355_/B vssd vssd vccd vccd _1356_/A sky130_fd_sc_hd__and2_1
XFILLER_4_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1286_ _1286_/A vssd vssd vccd vccd _1286_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1341__A _1341_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput550 _1146_/X vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__buf_12
XFILLER_5_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput561 _1166_/X vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__buf_12
XANTENNA__1516__A _1516_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput572 _1186_/X vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__buf_12
XFILLER_5_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput583 _1206_/X vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__buf_12
XFILLER_5_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput594 _0547_/Y vssd vssd vccd vccd la_data_in_mprj[102] sky130_fd_sc_hd__buf_12
XFILLER_8_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1235__B _1235_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input114_A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1077__A_N _1333_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3628 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1129__C _1129_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1145__B _1145_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2662 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1140_ _1140_/A vssd vssd vccd vccd _1140_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1071_ _1327_/A _1071_/B _1071_/C vssd vssd vccd vccd _1072_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3590 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] _0632_/X vssd vssd vccd vccd _1545_/A
+ sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_gates\[25\] mprj_dat_i_user[25] _0870_/X vssd vssd vccd vccd _0601_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_50_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0505__A _0505_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0924_ _0924_/A vssd vssd vccd vccd _0924_/X sky130_fd_sc_hd__buf_2
XFILLER_11_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0855_ _0855_/A _0855_/B vssd vssd vccd vccd _0856_/A sky130_fd_sc_hd__and2_1
XFILLER_11_1927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1039__C _1039_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0786_ _0786_/A vssd vssd vccd vccd _0786_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_2011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1336__A _1336_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1055__B _1055_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1407_ _1407_/A _1407_/B vssd vssd vccd vccd _1408_/A sky130_fd_sc_hd__and2_2
XANTENNA_user_wb_dat_gates\[27\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] _0854_/X vssd vssd vccd vccd _0568_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_29_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1338_ _1338_/A vssd vssd vccd vccd _1338_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1269_ _1525_/A _1269_/B _1269_/C vssd vssd vccd vccd _1270_/A sky130_fd_sc_hd__and3b_1
XFILLER_25_801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_322 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1246__A _1246_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[18\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input231_A la_iena_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input329_A la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0640_ _0640_/A vssd vssd vccd vccd _0640_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0979__B _0979_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0571_ _0571_/A vssd vssd vccd vccd _0571_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_49_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1156__A _1156_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0995__A _0995_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1123_ _1379_/A _1123_/B _1123_/C vssd vssd vccd vccd _1124_/A sky130_fd_sc_hd__and3b_4
XFILLER_1_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1054_ _1054_/A vssd vssd vccd vccd _1054_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0907_ _0907_/A _0907_/B vssd vssd vccd vccd _0908_/A sky130_fd_sc_hd__and2_2
X_0838_ _0838_/A vssd vssd vccd vccd _0838_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0889__B _0889_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0769_ _0769_/A _0769_/B vssd vssd vccd vccd _0770_/A sky130_fd_sc_hd__and2_4
XANTENNA__1066__A _1066_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput108 la_data_out_mprj[79] vssd vssd vccd vccd _1177_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput119 la_data_out_mprj[89] vssd vssd vccd vccd _1197_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2751 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1513__B _1513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1115__A_N _1371_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input181_A la_iena_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input279_A la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input446_A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1265__A_N _1521_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input42_A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1423__B _1423_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output498_A _1052_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output665_A _0496_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output832_A _1450_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0623_ _0623_/A _0623_/B vssd vssd vccd vccd _0624_/A sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0554_ _0554_/A vssd vssd vccd vccd _0554_/Y sky130_fd_sc_hd__clkinv_4
XTAP_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0485_ _0485_/A vssd vssd vccd vccd _0485_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_2902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1333__B _1333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1106_ _1106_/A vssd vssd vccd vccd _1106_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1037_ _1293_/A _1037_/B _1037_/C vssd vssd vccd vccd _1038_/A sky130_fd_sc_hd__and3b_2
XFILLER_22_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3008 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput90 la_data_out_mprj[62] vssd vssd vccd vccd _1143_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2086 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1243__B _1243_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input396_A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0603__A _0603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1137__C _1137_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3934 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1434__A _1434_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput450 mprj_dat_o_core[7] vssd vssd vccd vccd _0969_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput461 user_irq_ena[1] vssd vssd vccd vccd _0865_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1153__B _1153_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3644 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output782_A _1358_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0513__A _0513_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput902 _0605_/Y vssd vssd vccd vccd mprj_dat_i_core[29] sky130_fd_sc_hd__buf_12
XFILLER_29_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput913 _0956_/X vssd vssd vccd vccd mprj_dat_o_user[0] sky130_fd_sc_hd__buf_12
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput924 _0958_/X vssd vssd vccd vccd mprj_dat_o_user[1] sky130_fd_sc_hd__buf_12
Xoutput935 _0960_/X vssd vssd vccd vccd mprj_dat_o_user[2] sky130_fd_sc_hd__buf_12
XFILLER_9_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput946 _0886_/X vssd vssd vccd vccd mprj_sel_o_user[1] sky130_fd_sc_hd__buf_12
XFILLER_5_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0606_ _0606_/A vssd vssd vccd vccd _0606_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1047__C _1047_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput957 _0573_/Y vssd vssd vccd vccd user_irq[0] sky130_fd_sc_hd__buf_12
XFILLER_23_4040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0537_ _0537_/A vssd vssd vccd vccd _0537_/Y sky130_fd_sc_hd__inv_2
XTAP_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1344__A _1344_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0468_ _0468_/A vssd vssd vccd vccd _0468_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1063__B _1063_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1519__A _1519_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1254__A _1254_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input144_A la_iena_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input311_A la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input409_A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1429__A _1429_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1440_ _1440_/A vssd vssd vccd vccd _1440_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0987__B _0987_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output530_A _1110_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1371_ _1371_/A _1371_/B vssd vssd vccd vccd _1372_/A sky130_fd_sc_hd__and2_2
XFILLER_42_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output628_A _0463_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput280 la_oenb_mprj[118] vssd vssd vccd vccd _1511_/A sky130_fd_sc_hd__buf_2
Xinput291 la_oenb_mprj[12] vssd vssd vccd vccd _1299_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] _0692_/X vssd vssd vccd vccd _0487_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__0508__A _0508_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1339__A _1339_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput710 _0537_/Y vssd vssd vccd vccd la_data_in_mprj[92] sky130_fd_sc_hd__buf_12
Xoutput721 _1478_/X vssd vssd vccd vccd la_oenb_core[101] sky130_fd_sc_hd__buf_12
XFILLER_25_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput732 _1498_/X vssd vssd vccd vccd la_oenb_core[111] sky130_fd_sc_hd__buf_12
XFILLER_47_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput743 _1518_/X vssd vssd vccd vccd la_oenb_core[121] sky130_fd_sc_hd__buf_12
XFILLER_9_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput754 _1308_/X vssd vssd vccd vccd la_oenb_core[16] sky130_fd_sc_hd__buf_12
XANTENNA__0897__B _0897_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput765 _1328_/X vssd vssd vccd vccd la_oenb_core[26] sky130_fd_sc_hd__buf_12
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] _0616_/X vssd vssd vccd vccd _1537_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput776 _1348_/X vssd vssd vccd vccd la_oenb_core[36] sky130_fd_sc_hd__buf_12
XFILLER_28_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput787 _1368_/X vssd vssd vccd vccd la_oenb_core[46] sky130_fd_sc_hd__buf_12
XFILLER_25_2733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput798 _1388_/X vssd vssd vccd vccd la_oenb_core[56] sky130_fd_sc_hd__buf_12
XANTENNA__1074__A _1074_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2490 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1521__B _1521_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input261_A la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input359_A la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1783 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3898 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1431__B _1431_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3658 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0940_ _0940_/A vssd vssd vccd vccd _0940_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output480_A _1250_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0871_ input3/X _0871_/B vssd vssd vccd vccd _0872_/A sky130_fd_sc_hd__and2b_1
XANTENNA_output578_A _1198_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0998__A _0998_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1423_ _1423_/A _1423_/B vssd vssd vccd vccd _1424_/A sky130_fd_sc_hd__and2_1
XFILLER_20_4010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1354_ _1354_/A vssd vssd vccd vccd _1354_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_20_4054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1285_ _1285_/A _1285_/B vssd vssd vccd vccd _1286_/A sky130_fd_sc_hd__and2_4
XFILLER_37_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1341__B _1341_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0701__A _0701_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput540 _1128_/X vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__buf_12
XFILLER_47_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput551 _1148_/X vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__buf_12
XFILLER_9_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput562 _1168_/X vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__buf_12
Xoutput573 _1188_/X vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__buf_12
XFILLER_43_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput584 _1208_/X vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__buf_12
Xoutput595 _0548_/Y vssd vssd vccd vccd la_data_in_mprj[103] sky130_fd_sc_hd__buf_12
XFILLER_5_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1235__C _1235_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1251__B _1251_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input72_A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0611__A _0611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1145__C _1145_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2674 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1442__A _1442_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1070_ _1070_/A vssd vssd vccd vccd _1070_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_1225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1161__B _1161_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1021__A_N _1277_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output862_A _0936_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0923_ _0923_/A _0923_/B vssd vssd vccd vccd _0924_/A sky130_fd_sc_hd__and2_1
XFILLER_14_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1171__A_N _1427_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_gates\[18\] mprj_dat_i_user[18] _0870_/X vssd vssd vccd vccd _0594_/A
+ sky130_fd_sc_hd__nand2_2
X_0854_ _0854_/A vssd vssd vccd vccd _0854_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0785_ _0785_/A _0785_/B vssd vssd vccd vccd _0786_/A sky130_fd_sc_hd__and2_4
XFILLER_48_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0521__A _0521_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3656 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1055__C _1055_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1406_ _1406_/A vssd vssd vccd vccd _1406_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1337_ _1337_/A _1337_/B vssd vssd vccd vccd _1338_/A sky130_fd_sc_hd__and2_2
XFILLER_29_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1352__A _1352_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] _0840_/X vssd vssd vccd vccd _0561_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_39_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1268_ _1268_/A vssd vssd vccd vccd _1268_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1071__B _1071_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1199_ _1455_/A _1199_/B _1199_/C vssd vssd vccd vccd _1200_/A sky130_fd_sc_hd__and3b_2
XFILLER_52_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1527__A _1527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1262__A _1262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input224_A la_iena_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2943 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1437__A _1437_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0570_ _0570_/A vssd vssd vccd vccd _0570_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0995__B _0995_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output610_A _0562_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1122_ _1122_/A vssd vssd vccd vccd _1122_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1053_ _1309_/A _1053_/B _1053_/C vssd vssd vccd vccd _1054_/A sky130_fd_sc_hd__and3b_4
XFILLER_20_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0516__A _0516_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0906_ _0906_/A vssd vssd vccd vccd _0906_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0837_ _0837_/A _0837_/B vssd vssd vccd vccd _0838_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3646 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0768_ _0768_/A vssd vssd vccd vccd _0768_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_gates\[60\]_B _0728_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0699_ _0699_/A _0699_/B vssd vssd vccd vccd _0700_/A sky130_fd_sc_hd__and2_1
XFILLER_2_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput109 la_data_out_mprj[7] vssd vssd vccd vccd _1033_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__1067__A_N _1323_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1082__A _1082_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input174_A la_iena_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input341_A la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3908 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input439_A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input35_A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output658_A _0490_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0622_ _0622_/A vssd vssd vccd vccd _0622_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0553_ _0553_/A vssd vssd vccd vccd _0553_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output825_A _1436_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0484_ _0484_/A vssd vssd vccd vccd _0484_/Y sky130_fd_sc_hd__clkinv_2
XTAP_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] _0752_/X vssd vssd vccd vccd _0517_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_23_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1105_ _1361_/A _1105_/B _1105_/C vssd vssd vccd vccd _1106_/A sky130_fd_sc_hd__and3b_4
XFILLER_38_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1036_ _1036_/A vssd vssd vccd vccd _1036_/X sky130_fd_sc_hd__buf_2
XFILLER_39_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput80 la_data_out_mprj[53] vssd vssd vccd vccd _1125_/C sky130_fd_sc_hd__clkbuf_2
Xinput91 la_data_out_mprj[63] vssd vssd vccd vccd _1145_/C sky130_fd_sc_hd__buf_2
XFILLER_43_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1243__C _1243_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input291_A la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input389_A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_878 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput440 mprj_dat_o_core[27] vssd vssd vccd vccd _1009_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput451 mprj_dat_o_core[8] vssd vssd vccd vccd _0971_/B sky130_fd_sc_hd__clkbuf_4
Xinput462 user_irq_ena[2] vssd vssd vccd vccd _0867_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1153__C _1153_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output942_A _0970_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput903 _0578_/Y vssd vssd vccd vccd mprj_dat_i_core[2] sky130_fd_sc_hd__buf_12
XFILLER_7_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput914 _0976_/X vssd vssd vccd vccd mprj_dat_o_user[10] sky130_fd_sc_hd__buf_12
Xoutput925 _0996_/X vssd vssd vccd vccd mprj_dat_o_user[20] sky130_fd_sc_hd__buf_12
XFILLER_47_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput936 _1016_/X vssd vssd vccd vccd mprj_dat_o_user[30] sky130_fd_sc_hd__buf_12
XFILLER_25_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput947 _0888_/X vssd vssd vccd vccd mprj_sel_o_user[2] sky130_fd_sc_hd__buf_12
X_0605_ _0605_/A vssd vssd vccd vccd _0605_/Y sky130_fd_sc_hd__inv_2
Xoutput958 _0574_/Y vssd vssd vccd vccd user_irq[1] sky130_fd_sc_hd__buf_12
XFILLER_23_4052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0536_ _0536_/A vssd vssd vccd vccd _0536_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_3340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2959 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0467_ _0467_/A vssd vssd vccd vccd _0467_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_3384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1050 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2722 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1063__C _1063_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1105__A_N _1361_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1019_ _1275_/A _1019_/B input4/X vssd vssd vccd vccd _1020_/A sky130_fd_sc_hd__and3b_1
XFILLER_23_933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1255__A_N _1511_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1519__B _1519_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input137_A la_iena_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input304_A la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1429__B _1429_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1445__A _1445_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1370_ _1370_/A vssd vssd vccd vccd _1370_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_1729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output523_A _1098_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput270 la_oenb_mprj[109] vssd vssd vccd vccd _1493_/A sky130_fd_sc_hd__clkbuf_4
Xinput281 la_oenb_mprj[119] vssd vssd vccd vccd _1513_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput292 la_oenb_mprj[13] vssd vssd vccd vccd _1301_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output892_A _0577_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] _0678_/X vssd vssd vccd vccd _0480_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_20_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0524__A _0524_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1339__B _1339_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput700 _0528_/Y vssd vssd vccd vccd la_data_in_mprj[83] sky130_fd_sc_hd__buf_12
XFILLER_9_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput711 _0538_/Y vssd vssd vccd vccd la_data_in_mprj[93] sky130_fd_sc_hd__buf_12
Xoutput722 _1480_/X vssd vssd vccd vccd la_oenb_core[102] sky130_fd_sc_hd__buf_12
Xoutput733 _1500_/X vssd vssd vccd vccd la_oenb_core[112] sky130_fd_sc_hd__buf_12
Xoutput744 _1520_/X vssd vssd vccd vccd la_oenb_core[122] sky130_fd_sc_hd__buf_12
XFILLER_28_1101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput755 _1310_/X vssd vssd vccd vccd la_oenb_core[17] sky130_fd_sc_hd__buf_12
XFILLER_47_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1355__A _1355_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput766 _1330_/X vssd vssd vccd vccd la_oenb_core[27] sky130_fd_sc_hd__buf_12
Xoutput777 _1350_/X vssd vssd vccd vccd la_oenb_core[37] sky130_fd_sc_hd__buf_12
XFILLER_5_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput788 _1370_/X vssd vssd vccd vccd la_oenb_core[47] sky130_fd_sc_hd__buf_12
Xoutput799 _1390_/X vssd vssd vccd vccd la_oenb_core[57] sky130_fd_sc_hd__buf_12
XFILLER_28_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0519_ _0519_/A vssd vssd vccd vccd _0519_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1499_/A _1499_/B vssd vssd vccd vccd _1500_/A sky130_fd_sc_hd__and2_1
XFILLER_25_2789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1090__A _1090_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1249__B _1249_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input254_A la_iena_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input421_A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0609__A _0609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0870_ _0870_/A vssd vssd vccd vccd _0870_/X sky130_fd_sc_hd__buf_12
XANTENNA__1159__B _1159_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output473_A _1238_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output640_A _0474_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3755 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1422_ _1422_/A vssd vssd vccd vccd _1422_/X sky130_fd_sc_hd__buf_2
XFILLER_42_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1353_ _1353_/A _1353_/B vssd vssd vccd vccd _1354_/A sky130_fd_sc_hd__and2_1
XFILLER_24_3490 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4066 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1632 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1284_ _1284_/A vssd vssd vccd vccd _1284_/X sky130_fd_sc_hd__buf_2
XFILLER_49_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0519__A _0519_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1069__B _1069_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0999_ _0999_/A _0999_/B vssd vssd vccd vccd _1000_/A sky130_fd_sc_hd__and2_2
XFILLER_31_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2807 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0701__B _0701_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput530 _1110_/X vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__buf_12
Xoutput541 _1130_/X vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__buf_12
Xoutput552 _1150_/X vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__buf_12
Xoutput563 _1170_/X vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__buf_12
XFILLER_47_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput574 _1190_/X vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__buf_12
Xoutput585 _1210_/X vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__buf_12
XFILLER_25_2531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput596 _0549_/Y vssd vssd vccd vccd la_data_in_mprj[104] sky130_fd_sc_hd__buf_12
XFILLER_25_3287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1251__C _1251_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_582 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input371_A la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input65_A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2306 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1161__C _1161_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output590_A _1038_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0922_ _0922_/A vssd vssd vccd vccd _0922_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output855_A _0924_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0853_ _0853_/A _0853_/B vssd vssd vccd vccd _0854_/A sky130_fd_sc_hd__and2_1
XFILLER_48_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0802__A _0802_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0784_ _0784_/A vssd vssd vccd vccd _0784_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1405_ _1405_/A _1405_/B vssd vssd vccd vccd _1406_/A sky130_fd_sc_hd__and2_4
XFILLER_26_2873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[0\]_A mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1336_ _1336_/A vssd vssd vccd vccd _1336_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1080 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput1 caravel_clk vssd vssd vccd vccd input1/X sky130_fd_sc_hd__buf_6
X_1267_ _1523_/A _1267_/B _1267_/C vssd vssd vccd vccd _1268_/A sky130_fd_sc_hd__and3b_1
XFILLER_37_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] _0826_/X vssd vssd vccd vccd _0554_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_39_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1071__C _1071_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1198_ _1198_/A vssd vssd vccd vccd _1198_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1527__B _1527_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input217_A la_iena_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[0\] mprj_dat_i_user[0] _0870_/X vssd vssd vccd vccd _0576_/A sky130_fd_sc_hd__nand2_1
XFILLER_49_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1437__B _1437_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1121_ _1377_/A _1121_/B _1121_/C vssd vssd vccd vccd _1122_/A sky130_fd_sc_hd__and3b_4
XANTENNA_output603_A _0555_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1052_ _1052_/A vssd vssd vccd vccd _1052_/X sky130_fd_sc_hd__buf_4
XFILLER_4_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[30\] mprj_dat_i_user[30] _0870_/X vssd vssd vccd vccd _0606_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_33_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0905_ _0905_/A _0905_/B vssd vssd vccd vccd _0906_/A sky130_fd_sc_hd__and2_2
XFILLER_11_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0532__A _0532_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0836_ _0836_/A vssd vssd vccd vccd _0836_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1347__B _1347_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_4050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0767_ _0767_/A _0767_/B vssd vssd vccd vccd _0768_/A sky130_fd_sc_hd__and2_2
XFILLER_28_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0698_ _0698_/A vssd vssd vccd vccd _0698_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1319_ _1319_/A _1319_/B vssd vssd vccd vccd _1320_/A sky130_fd_sc_hd__and2_2
XFILLER_29_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0707__A _0707_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1257__B _1257_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input167_A la_iena_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input334_A la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input28_A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1161__A_N _1417_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0617__A _0617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1448__A _1448_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1167__B _1167_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0621_ _0621_/A _0621_/B vssd vssd vccd vccd _0622_/A sky130_fd_sc_hd__and2_1
XFILLER_45_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0552_ _0552_/A vssd vssd vccd vccd _0552_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output720_A _1476_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output818_A _1424_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0483_ _0483_/A vssd vssd vccd vccd _0483_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] _0738_/X vssd vssd vccd vccd _0510_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_3_2948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1104_ _1104_/A vssd vssd vccd vccd _1104_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0527__A _0527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1035_ _1291_/A _1035_/B _1035_/C vssd vssd vccd vccd _1036_/A sky130_fd_sc_hd__and3b_2
XFILLER_35_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_934 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1358__A _1358_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1077__B _1077_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput70 la_data_out_mprj[44] vssd vssd vccd vccd _1107_/C sky130_fd_sc_hd__clkbuf_1
X_0819_ _0819_/A _0819_/B vssd vssd vccd vccd _0820_/A sky130_fd_sc_hd__and2_2
Xinput81 la_data_out_mprj[54] vssd vssd vccd vccd _1127_/C sky130_fd_sc_hd__clkbuf_4
Xinput92 la_data_out_mprj[64] vssd vssd vccd vccd _1147_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_24_3308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1268__A _1268_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input284_A la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1066 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input451_A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__0900__A _0900_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput430 mprj_dat_o_core[18] vssd vssd vccd vccd _0991_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput441 mprj_dat_o_core[28] vssd vssd vccd vccd _1011_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_48_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput452 mprj_dat_o_core[9] vssd vssd vccd vccd _0973_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1057__A_N _1313_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output670_A _0501_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1178__A _1178_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output935_A _0960_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput904 _0606_/Y vssd vssd vccd vccd mprj_dat_i_core[30] sky130_fd_sc_hd__buf_12
XFILLER_28_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput915 _0978_/X vssd vssd vccd vccd mprj_dat_o_user[11] sky130_fd_sc_hd__buf_12
XFILLER_28_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput926 _0998_/X vssd vssd vccd vccd mprj_dat_o_user[21] sky130_fd_sc_hd__buf_12
Xoutput937 _1018_/X vssd vssd vccd vccd mprj_dat_o_user[31] sky130_fd_sc_hd__buf_12
XFILLER_45_3043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0604_ _0604_/A vssd vssd vccd vccd _0604_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0810__A _0810_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput948 _0890_/X vssd vssd vccd vccd mprj_sel_o_user[3] sky130_fd_sc_hd__buf_12
XFILLER_25_3639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput959 _0575_/Y vssd vssd vccd vccd user_irq[2] sky130_fd_sc_hd__buf_12
XTAP_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0535_ _0535_/A vssd vssd vccd vccd _0535_/Y sky130_fd_sc_hd__inv_2
XTAP_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4064 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0466_ _0466_/A vssd vssd vccd vccd _0466_/Y sky130_fd_sc_hd__inv_2
XTAP_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2662 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1018_ _1018_/A vssd vssd vccd vccd _1018_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_36_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1088__A _1088_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1954 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_783 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input95_A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1445__B _1445_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output516_A _1084_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput260 la_oenb_mprj[0] vssd vssd vccd vccd _1275_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1461__A _1461_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput271 la_oenb_mprj[10] vssd vssd vccd vccd _1295_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput282 la_oenb_mprj[11] vssd vssd vccd vccd _1297_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput293 la_oenb_mprj[14] vssd vssd vccd vccd _1303_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_1279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] _0664_/X vssd vssd vccd vccd _0473_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_53_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0805__A _0805_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput701 _0529_/Y vssd vssd vccd vccd la_data_in_mprj[84] sky130_fd_sc_hd__buf_12
Xoutput712 _0539_/Y vssd vssd vccd vccd la_data_in_mprj[94] sky130_fd_sc_hd__buf_12
XFILLER_9_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0540__A _0540_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput723 _1482_/X vssd vssd vccd vccd la_oenb_core[103] sky130_fd_sc_hd__buf_12
Xoutput734 _1502_/X vssd vssd vccd vccd la_oenb_core[113] sky130_fd_sc_hd__buf_12
XFILLER_29_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput745 _1522_/X vssd vssd vccd vccd la_oenb_core[123] sky130_fd_sc_hd__buf_12
Xoutput756 _1312_/X vssd vssd vccd vccd la_oenb_core[18] sky130_fd_sc_hd__buf_12
XANTENNA__1355__B _1355_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput767 _1332_/X vssd vssd vccd vccd la_oenb_core[28] sky130_fd_sc_hd__buf_12
XFILLER_5_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput778 _1352_/X vssd vssd vccd vccd la_oenb_core[38] sky130_fd_sc_hd__buf_12
XFILLER_29_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput789 _1372_/X vssd vssd vccd vccd la_oenb_core[48] sky130_fd_sc_hd__buf_12
XFILLER_28_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0518_ _0518_/A vssd vssd vccd vccd _0518_/Y sky130_fd_sc_hd__clkinv_2
XTAP_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1498_/A vssd vssd vccd vccd _1498_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_2779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1371__A _1371_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0715__A _0715_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1249__C _1249_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1265__B _1265_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input247_A la_iena_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1281__A _1281_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input414_A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0625__A _0625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1662 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1159__C _1159_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1456__A _1456_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1175__B _1175_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1421_ _1421_/A _1421_/B vssd vssd vccd vccd _1422_/A sky130_fd_sc_hd__and2_2
XANTENNA_output633_A _0467_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1352_ _1352_/A vssd vssd vccd vccd _1352_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1245__A_N _1501_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4078 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1283_ _1283_/A _1283_/B vssd vssd vccd vccd _1284_/A sky130_fd_sc_hd__and2_2
XFILLER_23_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0535__A _0535_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1069__C _1069_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0998_ _0998_/A vssd vssd vccd vccd _0998_/X sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1366__A _1366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput520 _1092_/X vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__buf_12
Xoutput531 _1112_/X vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__buf_12
XFILLER_9_3452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2819 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1085__B _1085_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput542 _1132_/X vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__buf_12
Xoutput553 _1152_/X vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__buf_12
XFILLER_43_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput564 _1172_/X vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__buf_12
Xoutput575 _1192_/X vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__buf_12
XFILLER_47_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2510 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput586 _1212_/X vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__buf_12
Xoutput597 _0550_/Y vssd vssd vccd vccd la_data_in_mprj[105] sky130_fd_sc_hd__buf_12
XFILLER_5_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input2_A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input197_A la_iena_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1276__A _1276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input364_A la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input58_A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1330 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0921_ _0921_/A _0921_/B vssd vssd vccd vccd _0922_/A sky130_fd_sc_hd__and2_1
XFILLER_35_2171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output583_A _1206_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0852_ _0852_/A vssd vssd vccd vccd _0852_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output848_A _0892_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0783_ _0783_/A _0783_/B vssd vssd vccd vccd _0784_/A sky130_fd_sc_hd__and2_4
XFILLER_48_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] _0798_/X vssd vssd vccd vccd _0540_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1404_ _1404_/A vssd vssd vccd vccd _1404_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[0\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1335_ _1335_/A _1335_/B vssd vssd vccd vccd _1336_/A sky130_fd_sc_hd__and2_2
XFILLER_29_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput2 caravel_clk2 vssd vssd vccd vccd input2/X sky130_fd_sc_hd__clkbuf_1
X_1266_ _1266_/A vssd vssd vccd vccd _1266_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1197_ _1453_/A _1197_/B _1197_/C vssd vssd vccd vccd _1198_/A sky130_fd_sc_hd__and3b_1
XFILLER_37_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1096__A _1096_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input112_A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1453__B _1453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1120_ _1120_/A vssd vssd vccd vccd _1120_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1051_ _1307_/A _1051_/B _1051_/C vssd vssd vccd vccd _1052_/A sky130_fd_sc_hd__and3b_1
XFILLER_18_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output798_A _1388_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[23\] mprj_dat_i_user[23] _0870_/X vssd vssd vccd vccd _0599_/A
+ sky130_fd_sc_hd__nand2_1
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] _0628_/X vssd vssd vccd vccd _1543_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_15_3298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0904_ _0904_/A vssd vssd vccd vccd _0904_/X sky130_fd_sc_hd__buf_6
XANTENNA__0813__A _0813_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0835_ _0835_/A _0835_/B vssd vssd vccd vccd _0836_/A sky130_fd_sc_hd__and2_2
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0766_ _0766_/A vssd vssd vccd vccd _0766_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0697_ _0697_/A _0697_/B vssd vssd vccd vccd _0698_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1363__B _1363_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] _0850_/X vssd vssd vccd vccd _0566_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_29_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1318_ _1318_/A vssd vssd vccd vccd _1318_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1249_ _1505_/A _1249_/B _1249_/C vssd vssd vccd vccd _1250_/A sky130_fd_sc_hd__and3b_2
XFILLER_38_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0707__B _0707_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0723__A _0723_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1257__C _1257_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1273__B _1273_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input327_A la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0617__B _0617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0633__A _0633_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_49_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0620_ _0620_/A vssd vssd vccd vccd _0620_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1167__C _1167_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0551_ _0551_/A vssd vssd vccd vccd _0551_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_output546_A _1030_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1464__A _1464_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1823 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0482_ _0482_/A vssd vssd vccd vccd _0482_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_3534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1183__B _1183_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1103_ _1359_/A _1103_/B _1103_/C vssd vssd vccd vccd _1104_/A sky130_fd_sc_hd__and3b_2
XFILLER_17_4006 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] _0724_/X vssd vssd vccd vccd _0503_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__0808__A _0808_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1034_ _1034_/A vssd vssd vccd vccd _1034_/X sky130_fd_sc_hd__buf_2
XFILLER_39_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_946 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0543__A _0543_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_28_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput60 la_data_out_mprj[35] vssd vssd vccd vccd _1089_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1077__C _1077_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput71 la_data_out_mprj[45] vssd vssd vccd vccd _1109_/C sky130_fd_sc_hd__clkbuf_1
X_0818_ _0818_/A vssd vssd vccd vccd _0818_/X sky130_fd_sc_hd__clkbuf_2
Xinput82 la_data_out_mprj[55] vssd vssd vccd vccd _1129_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput93 la_data_out_mprj[65] vssd vssd vccd vccd _1149_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0749_ _0749_/A _0749_/B vssd vssd vccd vccd _0750_/A sky130_fd_sc_hd__and2_1
XFILLER_48_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1374__A _1374_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1093__B _1093_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0718__A _0718_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input277_A la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1807 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1284__A _1284_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input444_A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input40_A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput420 mprj_cyc_o_core vssd vssd vccd vccd _0877_/B sky130_fd_sc_hd__clkbuf_8
Xinput431 mprj_dat_o_core[19] vssd vssd vccd vccd _0993_/B sky130_fd_sc_hd__clkbuf_4
Xinput442 mprj_dat_o_core[29] vssd vssd vccd vccd _1013_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_3177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput453 mprj_iena_wb vssd vssd vccd vccd _0869_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_48_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output496_A _1048_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1459__A _1459_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_2534 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput905 _0607_/Y vssd vssd vccd vccd mprj_dat_i_core[31] sky130_fd_sc_hd__buf_12
XFILLER_49_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput916 _0980_/X vssd vssd vccd vccd mprj_dat_o_user[12] sky130_fd_sc_hd__buf_12
XFILLER_29_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output830_A _1446_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput927 _1000_/X vssd vssd vccd vccd mprj_dat_o_user[22] sky130_fd_sc_hd__buf_12
X_0603_ _0603_/A vssd vssd vccd vccd _0603_/Y sky130_fd_sc_hd__inv_2
Xoutput938 _0962_/X vssd vssd vccd vccd mprj_dat_o_user[3] sky130_fd_sc_hd__buf_12
XANTENNA_output928_A _1002_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput949 _0880_/X vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__buf_12
XFILLER_45_3055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1194__A _1194_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2906 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0534_ _0534_/A vssd vssd vccd vccd _0534_/Y sky130_fd_sc_hd__clkinv_2
XTAP_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0465_ _0465_/A vssd vssd vccd vccd _0465_/Y sky130_fd_sc_hd__inv_2
XTAP_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1074 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2674 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0538__A _0538_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1017_ _1017_/A _1017_/B vssd vssd vccd vccd _1018_/A sky130_fd_sc_hd__and2_2
XFILLER_22_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1369__A _1369_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1151__A_N _1407_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1966 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1862 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1279__A _1279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input394_A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input88_A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0911__A _0911_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3684 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput250 la_iena_mprj[91] vssd vssd vccd vccd _0789_/B sky130_fd_sc_hd__clkbuf_1
Xinput261 la_oenb_mprj[100] vssd vssd vccd vccd _1475_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1461__B _1461_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput272 la_oenb_mprj[110] vssd vssd vccd vccd _1495_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput283 la_oenb_mprj[120] vssd vssd vccd vccd _1515_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output509_A _1072_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput294 la_oenb_mprj[15] vssd vssd vccd vccd _1305_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output780_A _1282_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output878_A _0908_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1690 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0821__A _0821_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput702 _0530_/Y vssd vssd vccd vccd la_data_in_mprj[85] sky130_fd_sc_hd__buf_12
Xoutput713 _0540_/Y vssd vssd vccd vccd la_data_in_mprj[95] sky130_fd_sc_hd__buf_12
Xoutput724 _1484_/X vssd vssd vccd vccd la_oenb_core[104] sky130_fd_sc_hd__buf_12
Xoutput735 _1504_/X vssd vssd vccd vccd la_oenb_core[114] sky130_fd_sc_hd__buf_12
Xoutput746 _1524_/X vssd vssd vccd vccd la_oenb_core[124] sky130_fd_sc_hd__buf_12
Xoutput757 _1314_/X vssd vssd vccd vccd la_oenb_core[19] sky130_fd_sc_hd__buf_12
XFILLER_47_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput768 _1334_/X vssd vssd vccd vccd la_oenb_core[29] sky130_fd_sc_hd__buf_12
Xoutput779 _1354_/X vssd vssd vccd vccd la_oenb_core[39] sky130_fd_sc_hd__buf_12
XFILLER_25_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2162 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0517_ _0517_/A vssd vssd vccd vccd _0517_/Y sky130_fd_sc_hd__inv_2
XTAP_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1497_ _1497_/A _1497_/B vssd vssd vccd vccd _1498_/A sky130_fd_sc_hd__and2_1
XTAP_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1371__B _1371_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1831 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0715__B _0715_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_242 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0731__A _0731_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1265__C _1265_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1047__A_N _1303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input142_A la_iena_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1281__B _1281_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input407_A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0906__A _0906_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0625__B _0625_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0641__A _0641_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1420_ _1420_/A vssd vssd vccd vccd _1420_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1175__C _1175_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1351_ _1351_/A _1351_/B vssd vssd vccd vccd _1352_/A sky130_fd_sc_hd__and2_2
XFILLER_20_4024 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1472__A _1472_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output626_A _1549_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1282_ _1282_/A vssd vssd vccd vccd _1282_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1191__B _1191_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] _0688_/X vssd vssd vccd vccd _0485_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__0816__A _0816_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0997_ _0997_/A _0997_/B vssd vssd vccd vccd _0998_/A sky130_fd_sc_hd__and2_2
XFILLER_30_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput510 _1074_/X vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__buf_12
Xoutput521 _1094_/X vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__buf_12
Xoutput532 _1114_/X vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__buf_12
XFILLER_44_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput543 _1134_/X vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__buf_12
XANTENNA__1085__C _1085_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput554 _1154_/X vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__buf_12
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] _0612_/X vssd vssd vccd vccd _1535_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput565 _1174_/X vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__buf_12
Xoutput576 _1194_/X vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__buf_12
XFILLER_25_2522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput587 _1214_/X vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__buf_12
XFILLER_47_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput598 _0551_/Y vssd vssd vccd vccd la_data_in_mprj[106] sky130_fd_sc_hd__buf_12
X_1549_ _1549_/A vssd vssd vccd vccd _1549_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__1382__A _1382_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_706 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input357_A la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1292__A _1292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ _0920_/A vssd vssd vccd vccd _0920_/X sky130_fd_sc_hd__buf_6
XFILLER_42_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0851_ _0851_/A _0851_/B vssd vssd vccd vccd _0852_/A sky130_fd_sc_hd__and2_1
XANTENNA_output576_A _1194_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2058 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1467__A _1467_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0782_ _0782_/A vssd vssd vccd vccd _0782_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output743_A _1518_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output910_A _0583_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1403_ _1403_/A _1403_/B vssd vssd vccd vccd _1404_/A sky130_fd_sc_hd__and2_1
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] _0784_/X vssd vssd vccd vccd _0533_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_3587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1334_ _1334_/A vssd vssd vccd vccd _1334_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1265_ _1521_/A _1265_/B _1265_/C vssd vssd vccd vccd _1266_/A sky130_fd_sc_hd__and3b_2
XFILLER_20_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput3 caravel_rstn vssd vssd vccd vccd input3/X sky130_fd_sc_hd__buf_12
XFILLER_7_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1196_ _1196_/A vssd vssd vccd vccd _1196_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0546__A _0546_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1377__A _1377_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3064 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2170 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input105_A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1235__A_N _1491_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__0903__B _0903_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1287__A _1287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input70_A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1050_ _1050_/A vssd vssd vccd vccd _1050_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output860_A _0932_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0903_ _0903_/A _0903_/B vssd vssd vccd vccd _0904_/A sky130_fd_sc_hd__and2_1
XANTENNA__0813__B _0813_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[16\] mprj_dat_i_user[16] _0870_/X vssd vssd vccd vccd _0592_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_31_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0834_ _0834_/A vssd vssd vccd vccd _0834_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0765_ _0765_/A _0765_/B vssd vssd vccd vccd _0766_/A sky130_fd_sc_hd__and2_4
XFILLER_6_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0696_ _0696_/A vssd vssd vccd vccd _0696_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3478 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1317_ _1317_/A _1317_/B vssd vssd vccd vccd _1318_/A sky130_fd_sc_hd__and2_2
XFILLER_29_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] _0836_/X vssd vssd vccd vccd _0559_/A
+ sky130_fd_sc_hd__nand2_1
X_1248_ _1248_/A vssd vssd vccd vccd _1248_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1179_ _1435_/A _1179_/B _1179_/C vssd vssd vccd vccd _1180_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0723__B _0723_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1273__C _1273_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input222_A la_iena_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0914__A _0914_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2142 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0633__B _0633_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0550_ _0550_/A vssd vssd vccd vccd _0550_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_3502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0481_ _0481_/A vssd vssd vccd vccd _0481_/Y sky130_fd_sc_hd__clkinv_2
XTAP_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1835 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1183__C _1183_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1868 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output706_A _0534_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1102_ _1102_/A vssd vssd vccd vccd _1102_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1033_ _1289_/A _1033_/B _1033_/C vssd vssd vccd vccd _1034_/A sky130_fd_sc_hd__and3b_2
XFILLER_35_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[20\]_A mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0824__A _0824_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_958 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3962 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput50 la_data_out_mprj[26] vssd vssd vccd vccd _1071_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0817_ _0817_/A _0817_/B vssd vssd vccd vccd _0818_/A sky130_fd_sc_hd__and2_4
Xinput61 la_data_out_mprj[36] vssd vssd vccd vccd _1091_/C sky130_fd_sc_hd__clkbuf_1
Xinput72 la_data_out_mprj[46] vssd vssd vccd vccd _1111_/C sky130_fd_sc_hd__clkbuf_1
Xinput83 la_data_out_mprj[56] vssd vssd vccd vccd _1131_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_28_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput94 la_data_out_mprj[66] vssd vssd vccd vccd _1151_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_28_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0748_ _0748_/A vssd vssd vccd vccd _0748_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0679_ _0679_/A _0679_/B vssd vssd vccd vccd _0680_/A sky130_fd_sc_hd__and2_1
XANTENNA__1093__C _1093_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1390__A _1390_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[11\]_A mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input172_A la_iena_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input437_A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput410 mprj_adr_o_core[2] vssd vssd vccd vccd _0895_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_40_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput421 mprj_dat_o_core[0] vssd vssd vccd vccd _0955_/B sky130_fd_sc_hd__buf_4
XFILLER_7_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input33_A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput432 mprj_dat_o_core[1] vssd vssd vccd vccd _0957_/B sky130_fd_sc_hd__buf_4
XFILLER_48_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput443 mprj_dat_o_core[2] vssd vssd vccd vccd _0959_/B sky130_fd_sc_hd__buf_2
XANTENNA__0909__A _0909_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput454 mprj_sel_o_core[0] vssd vssd vccd vccd _0883_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_5_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1459__B _1459_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output489_A _1266_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output656_A _0488_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1475__A _1475_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput906 _0579_/Y vssd vssd vccd vccd mprj_dat_i_core[3] sky130_fd_sc_hd__buf_12
Xoutput917 _0982_/X vssd vssd vccd vccd mprj_dat_o_user[13] sky130_fd_sc_hd__buf_12
X_0602_ _0602_/A vssd vssd vccd vccd _0602_/Y sky130_fd_sc_hd__inv_2
Xoutput928 _1002_/X vssd vssd vccd vccd mprj_dat_o_user[23] sky130_fd_sc_hd__buf_12
XFILLER_29_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput939 _0964_/X vssd vssd vccd vccd mprj_dat_o_user[4] sky130_fd_sc_hd__buf_12
XFILLER_45_3067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0533_ _0533_/A vssd vssd vccd vccd _0533_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4044 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0464_ _0464_/A vssd vssd vccd vccd _0464_/Y sky130_fd_sc_hd__inv_2
XTAP_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] _0748_/X vssd vssd vccd vccd _0515_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0819__A _0819_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1016_ _1016_/A vssd vssd vccd vccd _1016_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_23_903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1369__B _1369_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1385__A _1385_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2586 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0729__A _0729_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1279__B _1279_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input387_A la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__0911__B _0911_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1295__A _1295_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0639__A _0639_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput240 la_iena_mprj[82] vssd vssd vccd vccd _0771_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_48_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput251 la_iena_mprj[92] vssd vssd vccd vccd _0791_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput262 la_oenb_mprj[101] vssd vssd vccd vccd _1477_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput273 la_oenb_mprj[111] vssd vssd vccd vccd _1497_/A sky130_fd_sc_hd__buf_2
XFILLER_23_1259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput284 la_oenb_mprj[121] vssd vssd vccd vccd _1517_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput295 la_oenb_mprj[16] vssd vssd vccd vccd _1307_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1189__B _1189_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output940_A _0966_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0821__B _0821_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput703 _0531_/Y vssd vssd vccd vccd la_data_in_mprj[86] sky130_fd_sc_hd__buf_12
Xoutput714 _0541_/Y vssd vssd vccd vccd la_data_in_mprj[96] sky130_fd_sc_hd__buf_12
Xoutput725 _1486_/X vssd vssd vccd vccd la_oenb_core[105] sky130_fd_sc_hd__buf_12
XFILLER_47_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput736 _1506_/X vssd vssd vccd vccd la_oenb_core[115] sky130_fd_sc_hd__buf_12
XFILLER_29_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput747 _1526_/X vssd vssd vccd vccd la_oenb_core[125] sky130_fd_sc_hd__buf_12
Xoutput758 _1278_/X vssd vssd vccd vccd la_oenb_core[1] sky130_fd_sc_hd__buf_12
XFILLER_28_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput769 _1280_/X vssd vssd vccd vccd la_oenb_core[2] sky130_fd_sc_hd__buf_12
XFILLER_47_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0516_ _0516_/A vssd vssd vccd vccd _0516_/Y sky130_fd_sc_hd__inv_2
XTAP_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _1496_/A vssd vssd vccd vccd _1496_/X sky130_fd_sc_hd__clkbuf_2
XTAP_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_700 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1099__B _1099_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0731__B _0731_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input135_A la_iena_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input302_A la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0922__A _0922_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1350_ _1350_/A vssd vssd vccd vccd _1350_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output521_A _1094_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1281_ _1281_/A _1281_/B vssd vssd vccd vccd _1282_/A sky130_fd_sc_hd__and2_2
XFILLER_49_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output619_A _0570_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1191__C _1191_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1141__A_N _1397_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] _0674_/X vssd vssd vccd vccd _0478_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_18_3264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0996_ _0996_/A vssd vssd vccd vccd _0996_/X sky130_fd_sc_hd__buf_6
XFILLER_30_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput500 _1056_/X vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__buf_12
Xoutput511 _1076_/X vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__buf_12
Xoutput522 _1096_/X vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__buf_12
Xoutput533 _1116_/X vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__buf_12
XFILLER_47_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput544 _1136_/X vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__buf_12
Xoutput555 _1156_/X vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__buf_12
Xoutput566 _1176_/X vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__buf_12
XANTENNA_user_wb_dat_gates\[3\]_A mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput577 _1196_/X vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__buf_12
XFILLER_29_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput588 _1216_/X vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__buf_12
X_1548_ _1548_/A vssd vssd vccd vccd _1548_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_2534 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput599 _0552_/Y vssd vssd vccd vccd la_data_in_mprj[107] sky130_fd_sc_hd__buf_12
XFILLER_25_2556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1479_ _1479_/A _1479_/B vssd vssd vccd vccd _1480_/A sky130_fd_sc_hd__and2_1
XFILLER_41_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3684 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input252_A la_iena_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0850_ _0850_/A vssd vssd vccd vccd _0850_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1467__B _1467_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output471_A _1234_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0781_ _0781_/A _0781_/B vssd vssd vccd vccd _0782_/A sky130_fd_sc_hd__and2_1
XANTENNA_output569_A _1180_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1483__A _1483_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1402_ _1402_/A vssd vssd vccd vccd _1402_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_3649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2832 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output903_A _0578_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1333_ _1333_/A _1333_/B vssd vssd vccd vccd _1334_/A sky130_fd_sc_hd__and2_1
XFILLER_42_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1264_ _1264_/A vssd vssd vccd vccd _1264_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput4 la_data_out_mprj[0] vssd vssd vccd vccd input4/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__0827__A _0827_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1195_ _1451_/A _1195_/B _1195_/C vssd vssd vccd vccd _1196_/A sky130_fd_sc_hd__and3b_1
XFILLER_24_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0562__A _0562_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1037__A_N _1293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0979_ _0979_/A _0979_/B vssd vssd vccd vccd _0980_/A sky130_fd_sc_hd__and2_4
XFILLER_44_3600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1187__A_N _1443_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1393__A _1393_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1287__B _1287_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input63_A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3728 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0647__A _0647_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1478__A _1478_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0902_ _0902_/A vssd vssd vccd vccd _0902_/X sky130_fd_sc_hd__buf_4
XFILLER_15_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1197__B _1197_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0833_ _0833_/A _0833_/B vssd vssd vccd vccd _0834_/A sky130_fd_sc_hd__and2_1
XANTENNA_output853_A _0920_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0764_ _0764_/A vssd vssd vccd vccd _0764_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0695_ _0695_/A _0695_/B vssd vssd vccd vccd _0696_/A sky130_fd_sc_hd__and2_1
XFILLER_6_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1316_ _1316_/A vssd vssd vccd vccd _1316_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0557__A _0557_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1247_ _1503_/A _1247_/B _1247_/C vssd vssd vccd vccd _1248_/A sky130_fd_sc_hd__and3b_2
XFILLER_4_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] _0822_/X vssd vssd vccd vccd _0552_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_25_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1178_ _1178_/A vssd vssd vccd vccd _1178_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_606 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1388__A _1388_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3750 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input215_A la_iena_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1298__A _1298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0480_ _0480_/A vssd vssd vccd vccd _0480_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_3514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1101_ _1357_/A _1101_/B _1101_/C vssd vssd vccd vccd _1102_/A sky130_fd_sc_hd__and3b_4
XANTENNA_output601_A _0554_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1032_ _1032_/A vssd vssd vccd vccd _1032_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_47_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[20\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1001__A _1001_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput40 la_data_out_mprj[17] vssd vssd vccd vccd _1053_/C sky130_fd_sc_hd__clkbuf_1
X_0816_ _0816_/A vssd vssd vccd vccd _0816_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__0840__A _0840_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput51 la_data_out_mprj[27] vssd vssd vccd vccd _1073_/C sky130_fd_sc_hd__clkbuf_2
Xinput62 la_data_out_mprj[37] vssd vssd vccd vccd _1093_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput73 la_data_out_mprj[47] vssd vssd vccd vccd _1113_/C sky130_fd_sc_hd__clkbuf_2
Xinput84 la_data_out_mprj[57] vssd vssd vccd vccd _1133_/C sky130_fd_sc_hd__clkbuf_2
Xinput95 la_data_out_mprj[67] vssd vssd vccd vccd _1153_/C sky130_fd_sc_hd__buf_2
X_0747_ _0747_/A _0747_/B vssd vssd vccd vccd _0748_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0678_ _0678_/A vssd vssd vccd vccd _0678_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1225__A_N _1481_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[11\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input165_A la_iena_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput400 mprj_adr_o_core[20] vssd vssd vccd vccd _0931_/B sky130_fd_sc_hd__buf_6
Xinput411 mprj_adr_o_core[30] vssd vssd vccd vccd _0951_/B sky130_fd_sc_hd__buf_6
Xinput422 mprj_dat_o_core[10] vssd vssd vccd vccd _0975_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput433 mprj_dat_o_core[20] vssd vssd vccd vccd _0995_/B sky130_fd_sc_hd__buf_2
XFILLER_7_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input332_A la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput444 mprj_dat_o_core[30] vssd vssd vccd vccd _1015_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput455 mprj_sel_o_core[1] vssd vssd vccd vccd _0885_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__0909__B _0909_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input26_A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput907 _0580_/Y vssd vssd vccd vccd mprj_dat_i_core[4] sky130_fd_sc_hd__buf_12
X_0601_ _0601_/A vssd vssd vccd vccd _0601_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1475__B _1475_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput918 _0984_/X vssd vssd vccd vccd mprj_dat_o_user[14] sky130_fd_sc_hd__buf_12
Xoutput929 _1004_/X vssd vssd vccd vccd mprj_dat_o_user[24] sky130_fd_sc_hd__buf_12
XANTENNA_output649_A _0482_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0532_ _0532_/A vssd vssd vccd vccd _0532_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2919 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0463_ _0463_/A vssd vssd vccd vccd _0463_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_2389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1491__A _1491_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0819__B _0819_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] _0734_/X vssd vssd vccd vccd _0508_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_27_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1015_ _1015_/A _1015_/B vssd vssd vccd vccd _1016_/A sky130_fd_sc_hd__and2_2
XFILLER_35_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0835__A _0835_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1394 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1385__B _1385_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0729__B _0729_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0745__A _0745_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_414 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input282_A la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1295__B _1295_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput230 la_iena_mprj[73] vssd vssd vccd vccd _0753_/B sky130_fd_sc_hd__clkbuf_4
Xinput241 la_iena_mprj[83] vssd vssd vccd vccd _0773_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput252 la_iena_mprj[93] vssd vssd vccd vccd _0793_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_48_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput263 la_oenb_mprj[102] vssd vssd vccd vccd _1479_/A sky130_fd_sc_hd__clkbuf_4
Xinput274 la_oenb_mprj[112] vssd vssd vccd vccd _1499_/A sky130_fd_sc_hd__buf_2
XFILLER_49_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput285 la_oenb_mprj[122] vssd vssd vccd vccd _1519_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput296 la_oenb_mprj[17] vssd vssd vccd vccd _1309_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0655__A _0655_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_230 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output599_A _0552_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1189__C _1189_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output766_A _1330_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1486__A _1486_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output933_A _1012_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput704 _0532_/Y vssd vssd vccd vccd la_data_in_mprj[87] sky130_fd_sc_hd__buf_12
XFILLER_29_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput715 _0542_/Y vssd vssd vccd vccd la_data_in_mprj[97] sky130_fd_sc_hd__buf_12
Xoutput726 _1488_/X vssd vssd vccd vccd la_oenb_core[106] sky130_fd_sc_hd__buf_12
Xoutput737 _1508_/X vssd vssd vccd vccd la_oenb_core[116] sky130_fd_sc_hd__buf_12
XFILLER_47_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput748 _1528_/X vssd vssd vccd vccd la_oenb_core[126] sky130_fd_sc_hd__buf_12
XFILLER_7_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput759 _1316_/X vssd vssd vccd vccd la_oenb_core[20] sky130_fd_sc_hd__buf_12
XTAP_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0515_ _0515_/A vssd vssd vccd vccd _0515_/Y sky130_fd_sc_hd__inv_2
XTAP_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _1495_/A _1495_/B vssd vssd vccd vccd _1496_/A sky130_fd_sc_hd__and2_1
XFILLER_25_2749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1099__C _1099_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3866 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1396__A _1396_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input128_A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1093__A_N _1349_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input93_A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[9\] mprj_dat_i_user[9] _0870_/X vssd vssd vccd vccd _0585_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1280_ _1280_/A vssd vssd vccd vccd _1280_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_3336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output514_A _1080_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output883_A _0587_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] _0660_/X vssd vssd vccd vccd _0471_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_36_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0995_ _0995_/A _0995_/B vssd vssd vccd vccd _0996_/A sky130_fd_sc_hd__and2_4
XFILLER_53_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput501 _1058_/X vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__buf_12
Xoutput512 _1078_/X vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__buf_12
XFILLER_29_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput523 _1098_/X vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__buf_12
XFILLER_25_3203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput534 _1118_/X vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__buf_12
XFILLER_44_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput545 _1138_/X vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__buf_12
XFILLER_47_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput556 _1158_/X vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__buf_12
XANTENNA_user_wb_dat_gates\[3\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput567 _1178_/X vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__buf_12
XFILLER_5_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput578 _1198_/X vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__buf_12
Xoutput589 _1218_/X vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__buf_12
X_1547_ _1547_/A vssd vssd vccd vccd _1547_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_47_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1478_ _1478_/A vssd vssd vccd vccd _1478_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input245_A la_iena_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input412_A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0917__B _0917_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0933__A _0933_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0780_ _0780_/A vssd vssd vccd vccd _0780_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output464_A _1220_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1483__B _1483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1401_ _1401_/A _1401_/B vssd vssd vccd vccd _1402_/A sky130_fd_sc_hd__and2_2
XFILLER_29_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output631_A _0465_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1332_ _1332_/A vssd vssd vccd vccd _1332_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1263_ _1519_/A _1263_/B _1263_/C vssd vssd vccd vccd _1264_/A sky130_fd_sc_hd__and3b_2
XFILLER_20_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput5 la_data_out_mprj[100] vssd vssd vccd vccd input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_3177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0827__B _0827_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1194_ _1194_/A vssd vssd vccd vccd _1194_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1004__A _1004_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0843__A _0843_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0978_ _0978_/A vssd vssd vccd vccd _0978_/X sky130_fd_sc_hd__buf_6
XFILLER_27_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1393__B _1393_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0737__B _0737_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_306 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0753__A _0753_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_13_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input195_A la_iena_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1131__A_N _1387_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input362_A la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input56_A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3887 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0928__A _0928_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0647__B _0647_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0663__A _0663_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0901_ _0901_/A _0901_/B vssd vssd vccd vccd _0902_/A sky130_fd_sc_hd__and2_1
XANTENNA_output581_A _1202_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_32_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0832_ _0832_/A vssd vssd vccd vccd _0832_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0763_ _0763_/A _0763_/B vssd vssd vccd vccd _0764_/A sky130_fd_sc_hd__and2_4
XFILLER_31_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0694_ _0694_/A vssd vssd vccd vccd _0694_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] _0794_/X vssd vssd vccd vccd _0538_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_41_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1315_ _1315_/A _1315_/B vssd vssd vccd vccd _1316_/A sky130_fd_sc_hd__and2_4
XFILLER_42_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1246_ _1246_/A vssd vssd vccd vccd _1246_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1177_ _1433_/A _1177_/B _1177_/C vssd vssd vccd vccd _1178_/A sky130_fd_sc_hd__and3b_2
XFILLER_0_2378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_618 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_50_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3762 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input110_A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input208_A la_iena_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1763 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0658__A _0658_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1010 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1100_ _1100_/A vssd vssd vccd vccd _1100_/X sky130_fd_sc_hd__buf_4
XFILLER_1_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1027__A_N _1283_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1031_ _1287_/A _1031_/B _1031_/C vssd vssd vccd vccd _1032_/A sky130_fd_sc_hd__and3b_1
XFILLER_1_3399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1177__A_N _1433_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1489__A _1489_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[21\] mprj_dat_i_user[21] _0870_/X vssd vssd vccd vccd _0597_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_12_3953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1001__B _1001_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput30 la_data_out_mprj[123] vssd vssd vccd vccd _1265_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0815_ _0815_/A _0815_/B vssd vssd vccd vccd _0816_/A sky130_fd_sc_hd__and2_4
Xinput41 la_data_out_mprj[18] vssd vssd vccd vccd _1055_/C sky130_fd_sc_hd__clkbuf_2
Xinput52 la_data_out_mprj[28] vssd vssd vccd vccd _1075_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput63 la_data_out_mprj[38] vssd vssd vccd vccd _1095_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput74 la_data_out_mprj[48] vssd vssd vccd vccd _1115_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 la_data_out_mprj[58] vssd vssd vccd vccd _1135_/C sky130_fd_sc_hd__clkbuf_2
Xinput96 la_data_out_mprj[68] vssd vssd vccd vccd _1155_/C sky130_fd_sc_hd__clkbuf_4
X_0746_ _0746_/A vssd vssd vccd vccd _0746_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0677_ _0677_/A _0677_/B vssd vssd vccd vccd _0678_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0568__A _0568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1229_ _1485_/A _1229_/B _1229_/C vssd vssd vccd vccd _1230_/A sky130_fd_sc_hd__and3b_2
XFILLER_37_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1399__A _1399_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3886 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input158_A la_iena_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput401 mprj_adr_o_core[21] vssd vssd vccd vccd _0933_/B sky130_fd_sc_hd__clkbuf_16
Xinput412 mprj_adr_o_core[31] vssd vssd vccd vccd _0953_/B sky130_fd_sc_hd__buf_6
Xinput423 mprj_dat_o_core[11] vssd vssd vccd vccd _0977_/B sky130_fd_sc_hd__buf_2
Xinput434 mprj_dat_o_core[21] vssd vssd vccd vccd _0997_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput445 mprj_dat_o_core[31] vssd vssd vccd vccd _1017_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput456 mprj_sel_o_core[2] vssd vssd vccd vccd _0887_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input325_A la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input19_A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0925__B _0925_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1102__A _1102_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0941__A _0941_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0600_ _0600_/A vssd vssd vccd vccd _0600_/Y sky130_fd_sc_hd__inv_2
Xoutput908 _0581_/Y vssd vssd vccd vccd mprj_dat_i_core[5] sky130_fd_sc_hd__buf_12
Xoutput919 _0986_/X vssd vssd vccd vccd mprj_dat_o_user[15] sky130_fd_sc_hd__buf_12
XFILLER_45_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0531_ _0531_/A vssd vssd vccd vccd _0531_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_1571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output544_A _1136_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0462_ _0462_/A vssd vssd vccd vccd _0462_/Y sky130_fd_sc_hd__inv_2
XTAP_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1491__B _1491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output809_A _1408_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] _0720_/X vssd vssd vccd vccd _0501_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_35_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1014_ _1014_/A vssd vssd vccd vccd _1014_/X sky130_fd_sc_hd__buf_6
XANTENNA__0835__B _0835_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1012__A _1012_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0851__A _0851_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2074 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0729_ _0729_/A _0729_/B vssd vssd vccd vccd _0730_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4064 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0745__B _0745_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0761__A _0761_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input275_A la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input442_A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2931 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput220 la_iena_mprj[64] vssd vssd vccd vccd _0735_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput231 la_iena_mprj[74] vssd vssd vccd vccd _0755_/B sky130_fd_sc_hd__clkbuf_4
Xinput242 la_iena_mprj[84] vssd vssd vccd vccd _0775_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_2975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput253 la_iena_mprj[94] vssd vssd vccd vccd _0795_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput264 la_oenb_mprj[103] vssd vssd vccd vccd _1481_/A sky130_fd_sc_hd__buf_2
XFILLER_48_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput275 la_oenb_mprj[113] vssd vssd vccd vccd _1501_/A sky130_fd_sc_hd__buf_2
Xinput286 la_oenb_mprj[123] vssd vssd vccd vccd _1521_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput297 la_oenb_mprj[18] vssd vssd vccd vccd _1311_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__0936__A _0936_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output494_A _1044_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0671__A _0671_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1215__A_N _1471_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output661_A _0493_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output759_A _1316_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput705 _0533_/Y vssd vssd vccd vccd la_data_in_mprj[88] sky130_fd_sc_hd__buf_12
Xoutput716 _0543_/Y vssd vssd vccd vccd la_data_in_mprj[98] sky130_fd_sc_hd__buf_12
XFILLER_29_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput727 _1490_/X vssd vssd vccd vccd la_oenb_core[107] sky130_fd_sc_hd__buf_12
Xoutput738 _1510_/X vssd vssd vccd vccd la_oenb_core[117] sky130_fd_sc_hd__buf_12
Xoutput749 _1530_/X vssd vssd vccd vccd la_oenb_core[127] sky130_fd_sc_hd__buf_12
XANTENNA_output926_A _0998_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0514_ _0514_/A vssd vssd vccd vccd _0514_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _1494_/A vssd vssd vccd vccd _1494_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1007__A _1007_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3878 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[93\]_B _0794_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1744 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0756__A _0756_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_562 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input392_A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3366 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_B _0776_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input86_A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output876_A _0904_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1497__A _1497_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] _0646_/X vssd vssd vccd vccd _0464_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_32_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0994_ _0994_/A vssd vssd vccd vccd _0994_/X sky130_fd_sc_hd__buf_6
XFILLER_31_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput502 _1022_/X vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__buf_12
XFILLER_44_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput513 _1024_/X vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__buf_12
XFILLER_48_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput524 _1026_/X vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__buf_12
XFILLER_25_3215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput535 _1028_/X vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__buf_12
Xoutput546 _1030_/X vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__buf_12
XFILLER_44_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput557 _1032_/X vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__buf_12
XFILLER_5_3309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput568 _1034_/X vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__buf_12
XFILLER_47_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1546_ _1546_/A vssd vssd vccd vccd _1546_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_25_3259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput579 _1036_/X vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__buf_12
XFILLER_5_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1477_ _1477_/A _1477_/B vssd vssd vccd vccd _1478_/A sky130_fd_sc_hd__and2_1
XFILLER_3_3055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1200__A _1200_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input140_A la_iena_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input238_A la_iena_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input405_A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0933__B _0933_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1906 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[57\]_B _0722_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1110__A _1110_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1400_ _1400_/A vssd vssd vccd vccd _1400_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_2812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1331_ _1331_/A _1331_/B vssd vssd vccd vccd _1332_/A sky130_fd_sc_hd__and2_4
XFILLER_4_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output624_A _1547_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1262_ _1262_/A vssd vssd vccd vccd _1262_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput6 la_data_out_mprj[101] vssd vssd vccd vccd input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1193_ _1449_/A _1193_/B _1193_/C vssd vssd vccd vccd _1194_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0843__B _0843_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0977_ _0977_/A _0977_/B vssd vssd vccd vccd _0978_/A sky130_fd_sc_hd__and2_4
XFILLER_44_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] _1532_/X vssd vssd vccd vccd _1533_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_9_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1529_ _1529_/A _1529_/B vssd vssd vccd vccd _1530_/A sky130_fd_sc_hd__and2_1
XFILLER_47_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1083__A_N _1339_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0753__B _0753_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input188_A la_iena_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input355_A la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input49_A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0663__B _0663_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3258 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0900_ _0900_/A vssd vssd vccd vccd _0900_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0831_ _0831_/A _0831_/B vssd vssd vccd vccd _0832_/A sky130_fd_sc_hd__and2_1
XANTENNA_output574_A _1190_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0762_ _0762_/A vssd vssd vccd vccd _0762_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output741_A _1298_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output839_A _1462_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0693_ _0693_/A _0693_/B vssd vssd vccd vccd _0694_/A sky130_fd_sc_hd__and2_1
XFILLER_48_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] _0780_/X vssd vssd vccd vccd _0531_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_4_3150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1314_ _1314_/A vssd vssd vccd vccd _1314_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1245_ _1501_/A _1245_/B _1245_/C vssd vssd vccd vccd _1246_/A sky130_fd_sc_hd__and3b_1
XFILLER_49_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1015__A _1015_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[23\]_A mprj_dat_i_user[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1176_ _1176_/A vssd vssd vccd vccd _1176_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_B _0818_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_354 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[14\]_A mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0764__A _0764_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input103_A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1775 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0939__A _0939_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1226 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1022 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1030_ _1030_/A vssd vssd vccd vccd _1030_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0674__A _0674_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1489__B _1489_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output789_A _1372_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[14\] mprj_dat_i_user[14] _0870_/X vssd vssd vccd vccd _0590_/A
+ sky130_fd_sc_hd__nand2_1
Xinput20 la_data_out_mprj[114] vssd vssd vccd vccd _1247_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput31 la_data_out_mprj[124] vssd vssd vccd vccd _1267_/C sky130_fd_sc_hd__clkbuf_2
X_0814_ _0814_/A vssd vssd vccd vccd _0814_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput42 la_data_out_mprj[19] vssd vssd vccd vccd _1057_/C sky130_fd_sc_hd__clkbuf_1
Xinput53 la_data_out_mprj[29] vssd vssd vccd vccd _1077_/C sky130_fd_sc_hd__buf_2
Xinput64 la_data_out_mprj[39] vssd vssd vccd vccd _1097_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput75 la_data_out_mprj[49] vssd vssd vccd vccd _1117_/C sky130_fd_sc_hd__clkbuf_1
Xinput86 la_data_out_mprj[59] vssd vssd vccd vccd _1137_/C sky130_fd_sc_hd__clkbuf_2
X_0745_ _0745_/A _0745_/B vssd vssd vccd vccd _0746_/A sky130_fd_sc_hd__and2_1
Xinput97 la_data_out_mprj[69] vssd vssd vccd vccd _1157_/C sky130_fd_sc_hd__clkbuf_2
X_0676_ _0676_/A vssd vssd vccd vccd _0676_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0849__A _0849_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] _0832_/X vssd vssd vccd vccd _0557_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_26_903 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1228_ _1228_/A vssd vssd vccd vccd _1228_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_26_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1121__A_N _1377_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1159_ _1415_/A _1159_/B _1159_/C vssd vssd vccd vccd _1160_/A sky130_fd_sc_hd__and3b_1
XFILLER_39_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1399__B _1399_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3718 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3898 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1271__A_N _1527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0759__A _0759_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput402 mprj_adr_o_core[22] vssd vssd vccd vccd _0935_/B sky130_fd_sc_hd__buf_4
Xinput413 mprj_adr_o_core[3] vssd vssd vccd vccd _0897_/B sky130_fd_sc_hd__buf_6
XFILLER_2_3621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput424 mprj_dat_o_core[12] vssd vssd vccd vccd _0979_/B sky130_fd_sc_hd__clkbuf_2
Xinput435 mprj_dat_o_core[22] vssd vssd vccd vccd _0999_/B sky130_fd_sc_hd__clkbuf_4
Xinput446 mprj_dat_o_core[3] vssd vssd vccd vccd _0961_/B sky130_fd_sc_hd__buf_4
XFILLER_0_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput457 mprj_sel_o_core[3] vssd vssd vccd vccd _0889_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input220_A la_iena_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input318_A la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0494__A _0494_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0941__B _0941_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput909 _0582_/Y vssd vssd vccd vccd mprj_dat_i_core[6] sky130_fd_sc_hd__buf_12
XFILLER_45_3037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0530_ _0530_/A vssd vssd vccd vccd _0530_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0669__A _0669_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] _0706_/X vssd vssd vccd vccd _0494_/A
+ sky130_fd_sc_hd__nand2_1
X_1013_ _1013_/A _1013_/B vssd vssd vccd vccd _1014_/A sky130_fd_sc_hd__and2_2
XFILLER_34_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0851__B _0851_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2086 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0728_ _0728_/A vssd vssd vccd vccd _0728_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_2617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0659_ _0659_/A _0659_/B vssd vssd vccd vccd _0660_/A sky130_fd_sc_hd__and2_1
XFILLER_6_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4076 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0761__B _0761_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input170_A la_iena_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input268_A la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1167__A_N _1423_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input435_A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput210 la_iena_mprj[55] vssd vssd vccd vccd _0717_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input31_A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput221 la_iena_mprj[65] vssd vssd vccd vccd _0737_/B sky130_fd_sc_hd__clkbuf_1
Xinput232 la_iena_mprj[75] vssd vssd vccd vccd _0757_/B sky130_fd_sc_hd__buf_4
Xinput243 la_iena_mprj[85] vssd vssd vccd vccd _0777_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_2_3451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput254 la_iena_mprj[95] vssd vssd vccd vccd _0797_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput265 la_oenb_mprj[104] vssd vssd vccd vccd _1483_/A sky130_fd_sc_hd__buf_2
XFILLER_40_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput276 la_oenb_mprj[114] vssd vssd vccd vccd _1503_/A sky130_fd_sc_hd__clkbuf_4
Xinput287 la_oenb_mprj[124] vssd vssd vccd vccd _1523_/A sky130_fd_sc_hd__clkbuf_4
Xinput298 la_oenb_mprj[19] vssd vssd vccd vccd _1313_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3150 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output487_A _1262_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output654_A _0486_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput706 _0534_/Y vssd vssd vccd vccd la_data_in_mprj[89] sky130_fd_sc_hd__buf_12
Xoutput717 _0544_/Y vssd vssd vccd vccd la_data_in_mprj[99] sky130_fd_sc_hd__buf_12
XFILLER_10_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput728 _1492_/X vssd vssd vccd vccd la_oenb_core[108] sky130_fd_sc_hd__buf_12
Xoutput739 _1512_/X vssd vssd vccd vccd la_oenb_core[118] sky130_fd_sc_hd__buf_12
X_0513_ _0513_/A vssd vssd vccd vccd _0513_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output919_A _0986_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _1493_/A _1493_/B vssd vssd vccd vccd _1494_/A sky130_fd_sc_hd__and2_1
XTAP_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1007__B _1007_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0862__A _0862_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[6\]_A mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_574 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0772__A _0772_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1770 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input385_A la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input79_A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1108__A _1108_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0682__A _0682_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1497__B _1497_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0993_ _0993_/A _0993_/B vssd vssd vccd vccd _0994_/A sky130_fd_sc_hd__and2_4
XFILLER_34_1133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output869_A _0950_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput503 _1060_/X vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__buf_12
Xoutput514 _1080_/X vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__buf_12
XFILLER_44_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput525 _1100_/X vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__buf_12
XFILLER_48_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput536 _1120_/X vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__buf_12
XFILLER_47_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput547 _1140_/X vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__buf_12
XFILLER_5_990 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput558 _1160_/X vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__buf_12
X_1545_ _1545_/A vssd vssd vccd vccd _1545_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_2504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput569 _1180_/X vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__buf_12
XFILLER_47_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1018__A _1018_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1476_ _1476_/A vssd vssd vccd vccd _1476_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_1273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0857__A _0857_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0592__A _0592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0767__A _0767_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input133_A la_iena_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1205__A_N _1461_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input300_A la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1918 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1330_ _1330_/A vssd vssd vccd vccd _1330_/X sky130_fd_sc_hd__buf_2
XFILLER_8_3490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1582 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1261_ _1517_/A _1261_/B _1261_/C vssd vssd vccd vccd _1262_/A sky130_fd_sc_hd__and3b_1
XANTENNA__0677__A _0677_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output617_A _0568_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1192_ _1192_/A vssd vssd vccd vccd _1192_/X sky130_fd_sc_hd__clkbuf_4
Xinput7 la_data_out_mprj[102] vssd vssd vccd vccd input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] _0670_/X vssd vssd vccd vccd _0476_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_17_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1301__A _1301_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0976_ _0976_/A vssd vssd vccd vccd _0976_/X sky130_fd_sc_hd__buf_6
XFILLER_53_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1528_ _1528_/A vssd vssd vccd vccd _1528_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_1841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1459_ _1459_/A _1459_/B vssd vssd vccd vccd _1460_/A sky130_fd_sc_hd__and2_2
XFILLER_25_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input250_A la_iena_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input348_A la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0497__A _0497_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1105__B _1105_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0830_ _0830_/A vssd vssd vccd vccd _0830_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0960__A _0960_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0761_ _0761_/A _0761_/B vssd vssd vccd vccd _0762_/A sky130_fd_sc_hd__and2_4
XANTENNA_output567_A _1178_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0692_ _0692_/A vssd vssd vccd vccd _0692_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_2919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output734_A _1502_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1313_ _1313_/A _1313_/B vssd vssd vccd vccd _1314_/A sky130_fd_sc_hd__and2_2
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] _0766_/X vssd vssd vccd vccd _0524_/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_output901_A _0604_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1244_ _1244_/A vssd vssd vccd vccd _1244_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1015__B _1015_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1175_ _1431_/A _1175_/B _1175_/C vssd vssd vccd vccd _1176_/A sky130_fd_sc_hd__and3b_1
XANTENNA_user_wb_dat_gates\[23\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0959_ _0959_/A _0959_/B vssd vssd vccd vccd _0960_/A sky130_fd_sc_hd__and2_4
XFILLER_31_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1206__A _1206_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0780__A _0780_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input298_A la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input61_A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3686 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0939__B _0939_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1116__A _1116_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1073__A_N _1329_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput10 la_data_out_mprj[105] vssd vssd vccd vccd _1229_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_15_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output851_A _0916_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput21 la_data_out_mprj[115] vssd vssd vccd vccd _1249_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_0813_ _0813_/A _0813_/B vssd vssd vccd vccd _0814_/A sky130_fd_sc_hd__and2_4
Xinput32 la_data_out_mprj[125] vssd vssd vccd vccd _1269_/C sky130_fd_sc_hd__buf_2
XFILLER_11_1507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output949_A _0880_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput43 la_data_out_mprj[1] vssd vssd vccd vccd _1021_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput54 la_data_out_mprj[2] vssd vssd vccd vccd _1023_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput65 la_data_out_mprj[3] vssd vssd vccd vccd _1025_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 la_data_out_mprj[4] vssd vssd vccd vccd _1027_/C sky130_fd_sc_hd__clkbuf_1
X_0744_ _0744_/A vssd vssd vccd vccd _0744_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput87 la_data_out_mprj[5] vssd vssd vccd vccd _1029_/C sky130_fd_sc_hd__clkbuf_1
Xinput98 la_data_out_mprj[6] vssd vssd vccd vccd _1031_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0675_ _0675_/A _0675_/B vssd vssd vccd vccd _0676_/A sky130_fd_sc_hd__and2_1
XFILLER_48_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0849__B _0849_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1227_ _1483_/A _1227_/B input9/X vssd vssd vccd vccd _1228_/A sky130_fd_sc_hd__and3b_1
XANTENNA__0865__A _0865_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] _0818_/X vssd vssd vccd vccd _0550_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_17_3800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1158_ _1158_/A vssd vssd vccd vccd _1158_/X sky130_fd_sc_hd__buf_2
XFILLER_16_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj2_logic_high_inst output953/A vccd2_uq0 vssd2_uq0 mprj2_logic_high
X_1089_ _1345_/A _1089_/B _1089_/C vssd vssd vccd vccd _1090_/A sky130_fd_sc_hd__and3b_1
XFILLER_11_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0759__B _0759_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput403 mprj_adr_o_core[23] vssd vssd vccd vccd _0937_/B sky130_fd_sc_hd__buf_6
XFILLER_44_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput414 mprj_adr_o_core[4] vssd vssd vccd vccd _0899_/B sky130_fd_sc_hd__buf_8
XFILLER_0_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput425 mprj_dat_o_core[13] vssd vssd vccd vccd _0981_/B sky130_fd_sc_hd__clkbuf_2
Xinput436 mprj_dat_o_core[23] vssd vssd vccd vccd _1001_/B sky130_fd_sc_hd__clkbuf_4
Xinput447 mprj_dat_o_core[4] vssd vssd vccd vccd _0963_/B sky130_fd_sc_hd__buf_4
XFILLER_40_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput458 mprj_stb_o_core vssd vssd vccd vccd _0879_/B sky130_fd_sc_hd__buf_2
XFILLER_2_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0775__A _0775_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input213_A la_iena_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0685__A _0685_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1012_ _1012_/A vssd vssd vccd vccd _1012_/X sky130_fd_sc_hd__buf_6
XFILLER_19_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0727_ _0727_/A _0727_/B vssd vssd vccd vccd _0728_/A sky130_fd_sc_hd__and2_1
XFILLER_28_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0658_ _0658_/A vssd vssd vccd vccd _0658_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0589_ _0589_/A vssd vssd vccd vccd _0589_/Y sky130_fd_sc_hd__inv_2
XTAP_951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high_inst _0871_/B _1071_/B _1073_/B _1075_/B _1077_/B _1079_/B _1081_/B
+ _1083_/B _1085_/B _1087_/B _1089_/B _0891_/A _1091_/B _1093_/B _1095_/B _1097_/B
+ _1099_/B _1101_/B _1103_/B _1105_/B _1107_/B _1109_/B _0893_/A _1111_/B _1113_/B
+ _1115_/B _1117_/B _1119_/B _1121_/B _1123_/B _1125_/B _1127_/B _1129_/B _0895_/A
+ _1131_/B _1133_/B _1135_/B _1137_/B _1139_/B _1141_/B _1143_/B _1145_/B _1147_/B
+ _1149_/B _0897_/A _1151_/B _1153_/B _1155_/B _1157_/B _1159_/B _1161_/B _1163_/B
+ _1165_/B _1167_/B _1169_/B _0899_/A _1171_/B _1173_/B _1175_/B _1177_/B _1179_/B
+ _1181_/B _1183_/B _1185_/B _1187_/B _1189_/B _0901_/A _1191_/B _1193_/B _1195_/B
+ _1197_/B _1199_/B _1201_/B _1203_/B _1205_/B _1207_/B _1209_/B _0903_/A _1211_/B
+ _1213_/B _1215_/B _1217_/B _1219_/B _1221_/B _1223_/B _1225_/B _1227_/B _1229_/B
+ _0905_/A _1231_/B _1233_/B _1235_/B _1237_/B _1239_/B _1241_/B _1243_/B _1245_/B
+ _1247_/B _1249_/B _0907_/A _1251_/B _1253_/B _1255_/B _1257_/B _1259_/B _1261_/B
+ _1263_/B _1265_/B _1267_/B _1269_/B _0909_/A _0873_/A _1271_/B _1273_/B _1275_/B
+ _1277_/B _1279_/B _1281_/B _1283_/B _1285_/B _1287_/B _1289_/B _0911_/A _1291_/B
+ _1293_/B _1295_/B _1297_/B _1299_/B _1301_/B _1303_/B _1305_/B _1307_/B _1309_/B
+ _0913_/A _1311_/B _1313_/B _1315_/B _1317_/B _1319_/B _1321_/B _1323_/B _1325_/B
+ _1327_/B _1329_/B _0915_/A _1331_/B _1333_/B _1335_/B _1337_/B _1339_/B _1341_/B
+ _1343_/B _1345_/B _1347_/B _1349_/B _0917_/A _1351_/B _1353_/B _1355_/B _1357_/B
+ _1359_/B _1361_/B _1363_/B _1365_/B _1367_/B _1369_/B _0919_/A _1371_/B _1373_/B
+ _1375_/B _1377_/B _1379_/B _1381_/B _1383_/B _1385_/B _1387_/B _1389_/B _0921_/A
+ _1391_/B _1393_/B _1395_/B _1397_/B _1399_/B _1401_/B _1403_/B _1405_/B _1407_/B
+ _1409_/B _0923_/A _1411_/B _1413_/B _1415_/B _1417_/B _1419_/B _1421_/B _1423_/B
+ _1425_/B _1427_/B _1429_/B _0925_/A _1431_/B _1433_/B _1435_/B _1437_/B _1439_/B
+ _1441_/B _1443_/B _1445_/B _1447_/B _1449_/B _0927_/A _1451_/B _1453_/B _1455_/B
+ _1457_/B _1459_/B _1461_/B _1463_/B _1465_/B _1467_/B _1469_/B _0929_/A _0875_/A
+ _1471_/B _1473_/B _1475_/B _1477_/B _1479_/B _1481_/B _1483_/B _1485_/B _1487_/B
+ _1489_/B _0931_/A _1491_/B _1493_/B _1495_/B _1497_/B _1499_/B _1501_/B _1503_/B
+ _1505_/B _1507_/B _1509_/B _0933_/A _1511_/B _1513_/B _1515_/B _1517_/B _1519_/B
+ _1521_/B _1523_/B _1525_/B _1527_/B _1529_/B _0935_/A _1531_/A _0609_/A _0611_/A
+ _0613_/A _0615_/A _0617_/A _0619_/A _0621_/A _0623_/A _0625_/A _0937_/A _0627_/A
+ _0629_/A _0631_/A _0633_/A _0635_/A _0637_/A _0639_/A _0641_/A _0643_/A _0645_/A
+ _0939_/A _0647_/A _0649_/A _0651_/A _0653_/A _0655_/A _0657_/A _0659_/A _0661_/A
+ _0663_/A _0665_/A _0941_/A _0667_/A _0669_/A _0671_/A _0673_/A _0675_/A _0677_/A
+ _0679_/A _0681_/A _0683_/A _0685_/A _0943_/A _0687_/A _0689_/A _0691_/A _0693_/A
+ _0695_/A _0697_/A _0699_/A _0701_/A _0703_/A _0705_/A _0945_/A _0707_/A _0709_/A
+ _0711_/A _0713_/A _0715_/A _0717_/A _0719_/A _0721_/A _0723_/A _0725_/A _0947_/A
+ _0727_/A _0729_/A _0731_/A _0733_/A _0735_/A _0737_/A _0739_/A _0741_/A _0743_/A
+ _0745_/A _0949_/A _0877_/A _0747_/A _0749_/A _0751_/A _0753_/A _0755_/A _0757_/A
+ _0759_/A _0761_/A _0763_/A _0765_/A _0951_/A _0767_/A _0769_/A _0771_/A _0773_/A
+ _0775_/A _0777_/A _0779_/A _0781_/A _0783_/A _0785_/A _0953_/A _0787_/A _0789_/A
+ _0791_/A _0793_/A _0795_/A _0797_/A _0799_/A _0801_/A _0803_/A _0805_/A _0955_/A
+ _0807_/A _0809_/A _0811_/A _0813_/A _0815_/A _0817_/A _0819_/A _0821_/A _0823_/A
+ _0825_/A _0957_/A _0827_/A _0829_/A _0831_/A _0833_/A _0835_/A _0837_/A _0839_/A
+ _0841_/A _0843_/A _0845_/A _0959_/A _0847_/A _0849_/A _0851_/A _0853_/A _0855_/A
+ _0857_/A _0859_/A _0861_/A _0863_/A _0865_/A _0961_/A _0867_/A output951/A _0869_/A
+ _0963_/A _0965_/A _0967_/A _0969_/A _0879_/A _0971_/A _0973_/A _0975_/A _0977_/A
+ _0979_/A _0981_/A _0983_/A _0985_/A _0987_/A _0989_/A _0881_/A _0991_/A _0993_/A
+ _0995_/A _0997_/A _0999_/A _1001_/A _1003_/A _1005_/A _1007_/A _1009_/A _0883_/A
+ _1011_/A _1013_/A _1015_/A _1017_/A _1019_/B _1021_/B _1023_/B _1025_/B _1027_/B
+ _1029_/B _0885_/A _1031_/B _1033_/B _1035_/B _1037_/B _1039_/B _1041_/B _1043_/B
+ _1045_/B _1047_/B _1049_/B _0887_/A _1051_/B _1053_/B _1055_/B _1057_/B _1059_/B
+ _1061_/B _1063_/B _1065_/B _1067_/B _1069_/B _0889_/A vccd1_uq1 vssd1_uq1 mprj_logic_high
XFILLER_39_4033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0595__A _0595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1203__B _1203_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input163_A la_iena_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3634 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput200 la_iena_mprj[46] vssd vssd vccd vccd _0699_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput211 la_iena_mprj[56] vssd vssd vccd vccd _0719_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput222 la_iena_mprj[66] vssd vssd vccd vccd _0739_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput233 la_iena_mprj[76] vssd vssd vccd vccd _0759_/B sky130_fd_sc_hd__buf_2
XANTENNA_input330_A la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input428_A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput244 la_iena_mprj[86] vssd vssd vccd vccd _0779_/B sky130_fd_sc_hd__clkbuf_1
Xinput255 la_iena_mprj[96] vssd vssd vccd vccd _0799_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput266 la_oenb_mprj[105] vssd vssd vccd vccd _1485_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input24_A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput277 la_oenb_mprj[115] vssd vssd vccd vccd _1505_/A sky130_fd_sc_hd__buf_2
XFILLER_40_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput288 la_oenb_mprj[125] vssd vssd vccd vccd _1525_/A sky130_fd_sc_hd__buf_2
XFILLER_40_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput299 la_oenb_mprj[1] vssd vssd vccd vccd _1277_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1113__B _1113_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput707 _1541_/Y vssd vssd vccd vccd la_data_in_mprj[8] sky130_fd_sc_hd__buf_12
XFILLER_10_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput718 _1542_/Y vssd vssd vccd vccd la_data_in_mprj[9] sky130_fd_sc_hd__buf_12
Xoutput729 _1494_/X vssd vssd vccd vccd la_oenb_core[109] sky130_fd_sc_hd__buf_12
XFILLER_10_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output647_A _0480_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1111__A_N _1367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0512_ _0512_/A vssd vssd vccd vccd _0512_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1492_ _1492_/A vssd vssd vccd vccd _1492_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1261__A_N _1517_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] _0730_/X vssd vssd vccd vccd _0506_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_3_2548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1304__A _1304_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1023__B _1023_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[6\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1214__A _1214_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input280_A la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input378_A la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0947__B _0947_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1124__A _1124_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output597_A _0550_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0992_ _0992_/A vssd vssd vccd vccd _0992_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_35_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output931_A _1008_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput504 _1062_/X vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__buf_12
XFILLER_29_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput515 _1082_/X vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__buf_12
XFILLER_44_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput526 _1102_/X vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__buf_12
Xoutput537 _1122_/X vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__buf_12
Xoutput548 _1142_/X vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__buf_12
XFILLER_5_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput559 _1162_/X vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__buf_12
X_1544_ _1544_/A vssd vssd vccd vccd _1544_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_3239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1475_ _1475_/A _1475_/B vssd vssd vccd vccd _1476_/A sky130_fd_sc_hd__and2_1
XFILLER_42_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0857__B _0857_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1034__A _1034_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0873__A _0873_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1157__A_N _1413_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3604 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0767__B _0767_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input126_A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0783__A _0783_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XTAP_1777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input91_A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[7\] mprj_dat_i_user[7] _0870_/X vssd vssd vccd vccd _0583_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1260_ _1260_/A vssd vssd vccd vccd _1260_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0677__B _0677_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output512_A _1078_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1191_ _1447_/A _1191_/B _1191_/C vssd vssd vccd vccd _1192_/A sky130_fd_sc_hd__and3b_1
XFILLER_20_3169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput8 la_data_out_mprj[103] vssd vssd vccd vccd input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0693__A _0693_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output881_A _0576_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_33_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] _0656_/X vssd vssd vccd vccd _0469_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__1301__B _1301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0975_ _0975_/A _0975_/B vssd vssd vccd vccd _0976_/A sky130_fd_sc_hd__and2_2
XFILLER_31_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1527_ _1527_/A _1527_/B vssd vssd vccd vccd _1528_/A sky130_fd_sc_hd__and2_2
XFILLER_47_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1458_ _1458_/A vssd vssd vccd vccd _1458_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1389_ _1389_/A _1389_/B vssd vssd vccd vccd _1390_/A sky130_fd_sc_hd__and2_1
XFILLER_42_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_23_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1211__B _1211_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0778__A _0778_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput890 _0594_/Y vssd vssd vccd vccd mprj_dat_i_core[18] sky130_fd_sc_hd__buf_12
XFILLER_43_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input243_A la_iena_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2170 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input410_A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1105__C _1105_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1402__A _1402_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1121__B _1121_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0760_ _0760_/A vssd vssd vccd vccd _0760_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0691_ _0691_/A _0691_/B vssd vssd vccd vccd _0692_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output727_A _1490_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1312_ _1312_/A vssd vssd vccd vccd _1312_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_2688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1243_ _1499_/A _1243_/B _1243_/C vssd vssd vccd vccd _1244_/A sky130_fd_sc_hd__and3b_2
XFILLER_49_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1174_ _1174_/A vssd vssd vccd vccd _1174_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1312__A _1312_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1031__B _1031_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0958_ _0958_/A vssd vssd vccd vccd _0958_/X sky130_fd_sc_hd__buf_6
XFILLER_21_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0889_ _0889_/A _0889_/B vssd vssd vccd vccd _0890_/A sky130_fd_sc_hd__and2_4
XFILLER_31_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1222__A _1222_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input193_A la_iena_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input360_A la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input458_A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input54_A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2931 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3990 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0955__B _0955_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xpowergood_check output954/A output952/A vccd vssd vdda1_uq0 vssa1_uq0 vdda2_uq0 vssa2_uq0
+ mgmt_protect_hv
XFILLER_46_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1132__A _1132_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0971__A _0971_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput11 la_data_out_mprj[106] vssd vssd vccd vccd _1231_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_0812_ _0812_/A vssd vssd vccd vccd _0812_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput22 la_data_out_mprj[116] vssd vssd vccd vccd _1251_/C sky130_fd_sc_hd__clkbuf_2
Xinput33 la_data_out_mprj[126] vssd vssd vccd vccd _1271_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput44 la_data_out_mprj[20] vssd vssd vccd vccd _1059_/C sky130_fd_sc_hd__clkbuf_2
Xinput55 la_data_out_mprj[30] vssd vssd vccd vccd _1079_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_10_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output844_A _1472_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput66 la_data_out_mprj[40] vssd vssd vccd vccd _1099_/C sky130_fd_sc_hd__clkbuf_2
X_0743_ _0743_/A _0743_/B vssd vssd vccd vccd _0744_/A sky130_fd_sc_hd__and2_1
Xinput77 la_data_out_mprj[50] vssd vssd vccd vccd _1119_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_28_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput88 la_data_out_mprj[60] vssd vssd vccd vccd _1139_/C sky130_fd_sc_hd__buf_2
Xinput99 la_data_out_mprj[70] vssd vssd vccd vccd _1159_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0674_ _0674_/A vssd vssd vccd vccd _0674_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] _0790_/X vssd vssd vccd vccd _0536_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_48_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1307__A _1307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1226_ _1226_/A vssd vssd vccd vccd _1226_/X sky130_fd_sc_hd__buf_2
XFILLER_6_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0865__B _0865_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1157_ _1413_/A _1157_/B _1157_/C vssd vssd vccd vccd _1158_/A sky130_fd_sc_hd__and3b_1
XANTENNA__1042__A _1042_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1088_ _1088_/A vssd vssd vccd vccd _1088_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_12_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0881__A _0881_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput404 mprj_adr_o_core[24] vssd vssd vccd vccd _0939_/B sky130_fd_sc_hd__buf_8
Xinput415 mprj_adr_o_core[5] vssd vssd vccd vccd _0901_/B sky130_fd_sc_hd__buf_8
XFILLER_40_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput426 mprj_dat_o_core[14] vssd vssd vccd vccd _0983_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_6_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput437 mprj_dat_o_core[24] vssd vssd vccd vccd _1003_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput448 mprj_dat_o_core[5] vssd vssd vccd vccd _0965_/B sky130_fd_sc_hd__buf_4
XFILLER_40_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput459 mprj_we_o_core vssd vssd vccd vccd _0881_/B sky130_fd_sc_hd__buf_2
XFILLER_2_2911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0775__B _0775_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input206_A la_iena_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0791__A _0791_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0685__B _0685_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1011_ _1011_/A _1011_/B vssd vssd vccd vccd _1012_/A sky130_fd_sc_hd__and2_2
XFILLER_47_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0726_ _0726_/A vssd vssd vccd vccd _0726_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0657_ _0657_/A _0657_/B vssd vssd vccd vccd _0658_/A sky130_fd_sc_hd__and2_1
XFILLER_41_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0588_ _0588_/A vssd vssd vccd vccd _0588_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_3_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0876__A _0876_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1209_ _1465_/A _1209_/B _1209_/C vssd vssd vccd vccd _1210_/A sky130_fd_sc_hd__and3b_4
XTAP_2819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_628 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input156_A la_iena_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput201 la_iena_mprj[47] vssd vssd vccd vccd _0701_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_3679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput212 la_iena_mprj[57] vssd vssd vccd vccd _0721_/B sky130_fd_sc_hd__buf_2
XFILLER_40_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0786__A _0786_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput223 la_iena_mprj[67] vssd vssd vccd vccd _0741_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput234 la_iena_mprj[77] vssd vssd vccd vccd _0761_/B sky130_fd_sc_hd__buf_2
XFILLER_2_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput245 la_iena_mprj[87] vssd vssd vccd vccd _0781_/B sky130_fd_sc_hd__buf_4
XFILLER_40_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput256 la_iena_mprj[97] vssd vssd vccd vccd _0801_/B sky130_fd_sc_hd__clkbuf_1
Xinput267 la_oenb_mprj[106] vssd vssd vccd vccd _1487_/A sky130_fd_sc_hd__buf_4
XANTENNA_input323_A la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1063__A_N _1319_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput278 la_oenb_mprj[116] vssd vssd vccd vccd _1507_/A sky130_fd_sc_hd__buf_2
XFILLER_5_1141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput289 la_oenb_mprj[126] vssd vssd vccd vccd _1527_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input17_A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1113__C _1113_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_82 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2142 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1410__A _1410_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput708 _0535_/Y vssd vssd vccd vccd la_data_in_mprj[90] sky130_fd_sc_hd__buf_12
Xoutput719 _1276_/X vssd vssd vccd vccd la_oenb_core[0] sky130_fd_sc_hd__buf_12
X_0511_ _0511_/A vssd vssd vccd vccd _0511_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1491_ _1491_/A _1491_/B vssd vssd vccd vccd _1492_/A sky130_fd_sc_hd__and2_1
XFILLER_25_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output807_A _1404_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] _0716_/X vssd vssd vccd vccd _0499_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_48_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1023__C _1023_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1320__A _1320_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0709_ _0709_/A _0709_/B vssd vssd vccd vccd _0710_/A sky130_fd_sc_hd__and2_1
XFILLER_47_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1610 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1230__A _1230_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input273_A la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input440_A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1405__A _1405_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0963__B _0963_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1140__A _1140_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output492_A _1272_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0991_ _0991_/A _0991_/B vssd vssd vccd vccd _0992_/A sky130_fd_sc_hd__and2_4
XFILLER_31_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output757_A _1314_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput505 _1064_/X vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__buf_12
Xoutput516 _1084_/X vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__buf_12
Xoutput527 _1104_/X vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__buf_12
XFILLER_9_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput538 _1124_/X vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__buf_12
XANTENNA_output924_A _0958_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1543_ _1543_/A vssd vssd vccd vccd _1543_/Y sky130_fd_sc_hd__inv_2
Xoutput549 _1144_/X vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__buf_12
XFILLER_29_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1474_ _1474_/A vssd vssd vccd vccd _1474_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3830 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1315__A _1315_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3896 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0873__B input1/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1050__A _1050_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1209__B _1209_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3616 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__0783__B _0783_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1101__A_N _1357_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_546 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input390_A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1251__A_N _1507_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input84_A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1190_ _1190_/A vssd vssd vccd vccd _1190_/X sky130_fd_sc_hd__buf_2
Xinput9 la_data_out_mprj[104] vssd vssd vccd vccd input9/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0974__A _0974_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output505_A _1064_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0693__B _0693_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output874_A _0900_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] _0642_/X vssd vssd vccd vccd _0462_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_20_549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0974_ _0974_/A vssd vssd vccd vccd _0974_/X sky130_fd_sc_hd__buf_6
XFILLER_9_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1029__B _1029_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1526_ _1526_/A vssd vssd vccd vccd _1526_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1457_ _1457_/A _1457_/B vssd vssd vccd vccd _1458_/A sky130_fd_sc_hd__and2_2
XFILLER_29_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[26\]_A mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1388_ _1388_/A vssd vssd vccd vccd _1388_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0884__A _0884_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput880 _0878_/X vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__buf_12
Xoutput891 _0595_/Y vssd vssd vccd vccd mprj_dat_i_core[19] sky130_fd_sc_hd__buf_12
XFILLER_43_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[17\]_A mprj_dat_i_user[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input236_A la_iena_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0794__A _0794_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input403_A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1121__C _1121_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0690_ _0690_/A vssd vssd vccd vccd _0690_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0969__A _0969_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1139 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1311_ _1311_/A _1311_/B vssd vssd vccd vccd _1312_/A sky130_fd_sc_hd__and2_4
XFILLER_46_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1147__A_N _1403_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1242_ _1242_/A vssd vssd vccd vccd _1242_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1173_ _1429_/A _1173_/B _1173_/C vssd vssd vccd vccd _1174_/A sky130_fd_sc_hd__and3b_2
XTAP_4190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1031__C _1031_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0957_ _0957_/A _0957_/B vssd vssd vccd vccd _0958_/A sky130_fd_sc_hd__and2_1
XFILLER_9_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0888_ _0888_/A vssd vssd vccd vccd _0888_/X sky130_fd_sc_hd__buf_8
XFILLER_44_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0879__A _0879_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1509_ _1509_/A _1509_/B vssd vssd vccd vccd _1510_/A sky130_fd_sc_hd__and2_1
XFILLER_26_3891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1503__A _1503_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input186_A la_iena_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0789__A _0789_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input353_A la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2943 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input47_A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1413__A _1413_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0971__B _0971_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0811_ _0811_/A _0811_/B vssd vssd vccd vccd _0812_/A sky130_fd_sc_hd__and2_4
XFILLER_35_1082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output572_A _1186_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput12 la_data_out_mprj[107] vssd vssd vccd vccd _1233_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_30_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput23 la_data_out_mprj[117] vssd vssd vccd vccd _1253_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 la_data_out_mprj[127] vssd vssd vccd vccd _1273_/C sky130_fd_sc_hd__clkbuf_2
Xinput45 la_data_out_mprj[21] vssd vssd vccd vccd _1061_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_0742_ _0742_/A vssd vssd vccd vccd _0742_/X sky130_fd_sc_hd__clkbuf_1
Xinput56 la_data_out_mprj[31] vssd vssd vccd vccd _1081_/C sky130_fd_sc_hd__clkbuf_1
Xinput67 la_data_out_mprj[41] vssd vssd vccd vccd _1101_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_10_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput78 la_data_out_mprj[51] vssd vssd vccd vccd _1121_/C sky130_fd_sc_hd__clkbuf_2
Xinput89 la_data_out_mprj[61] vssd vssd vccd vccd _1141_/C sky130_fd_sc_hd__buf_2
XANTENNA__0699__A _0699_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0673_ _0673_/A _0673_/B vssd vssd vccd vccd _0674_/A sky130_fd_sc_hd__and2_1
XFILLER_48_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] _0776_/X vssd vssd vccd vccd _0529_/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA__1307__B _1307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1225_ _1481_/A _1225_/B input8/X vssd vssd vccd vccd _1226_/A sky130_fd_sc_hd__and3b_4
XFILLER_38_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1323__A _1323_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1156_ _1156_/A vssd vssd vccd vccd _1156_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1087_ _1343_/A _1087_/B _1087_/C vssd vssd vccd vccd _1088_/A sky130_fd_sc_hd__and3b_1
XFILLER_41_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0881__B _0881_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1217__B _1217_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput405 mprj_adr_o_core[25] vssd vssd vccd vccd _0941_/B sky130_fd_sc_hd__buf_8
XFILLER_2_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput416 mprj_adr_o_core[6] vssd vssd vccd vccd _0903_/B sky130_fd_sc_hd__buf_6
XFILLER_22_3541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput427 mprj_dat_o_core[15] vssd vssd vccd vccd _0985_/B sky130_fd_sc_hd__buf_4
XFILLER_6_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput438 mprj_dat_o_core[25] vssd vssd vccd vccd _1005_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput449 mprj_dat_o_core[6] vssd vssd vccd vccd _0967_/B sky130_fd_sc_hd__buf_4
XFILLER_2_2901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4046 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input101_A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1408__A _1408_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1127__B _1127_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1010_ _1010_/A vssd vssd vccd vccd _1010_/X sky130_fd_sc_hd__buf_6
XFILLER_40_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0982__A _0982_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output954_A output954/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[12\] mprj_dat_i_user[12] _0870_/X vssd vssd vccd vccd _0588_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_8_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0725_ _0725_/A _0725_/B vssd vssd vccd vccd _0726_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1318__A _1318_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0656_ _0656_/A vssd vssd vccd vccd _0656_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1037__B _1037_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0587_ _0587_/A vssd vssd vccd vccd _0587_/Y sky130_fd_sc_hd__inv_2
XTAP_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2294 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] _0828_/X vssd vssd vccd vccd _0555_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_27_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1208_ _1208_/A vssd vssd vccd vccd _1208_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1139_ _1395_/A _1139_/B _1139_/C vssd vssd vccd vccd _1140_/A sky130_fd_sc_hd__and3b_4
XFILLER_26_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_A mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput202 la_iena_mprj[48] vssd vssd vccd vccd _0703_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_4072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput213 la_iena_mprj[58] vssd vssd vccd vccd _0723_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput224 la_iena_mprj[68] vssd vssd vccd vccd _0743_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_49_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input149_A la_iena_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput235 la_iena_mprj[78] vssd vssd vccd vccd _0763_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput246 la_iena_mprj[88] vssd vssd vccd vccd _0783_/B sky130_fd_sc_hd__clkbuf_1
Xinput257 la_iena_mprj[98] vssd vssd vccd vccd _0803_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput268 la_oenb_mprj[107] vssd vssd vccd vccd _1489_/A sky130_fd_sc_hd__clkbuf_4
Xinput279 la_oenb_mprj[117] vssd vssd vccd vccd _1509_/A sky130_fd_sc_hd__buf_2
XFILLER_40_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input316_A la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_94 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput709 _0536_/Y vssd vssd vccd vccd la_data_in_mprj[91] sky130_fd_sc_hd__buf_12
XFILLER_29_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1138__A _1138_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0510_ _0510_/A vssd vssd vccd vccd _0510_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1490_ _1490_/A vssd vssd vccd vccd _1490_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output535_A _1028_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0977__A _0977_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2478 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] _0702_/X vssd vssd vccd vccd _0492_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_47_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1048__A _1048_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0708_ _0708_/A vssd vssd vccd vccd _0708_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_3934 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] _0626_/X vssd vssd vccd vccd _1542_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_28_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0887__A _0887_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0639_ _0639_/A _0639_/B vssd vssd vccd vccd _0640_/A sky130_fd_sc_hd__and2_1
XFILLER_28_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1511__A _1511_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input266_A la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0797__A _0797_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input433_A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1405__B _1405_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1421__A _1421_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0990_ _0990_/A vssd vssd vccd vccd _0990_/X sky130_fd_sc_hd__buf_6
XFILLER_53_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput506 _1066_/X vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__buf_12
Xoutput517 _1086_/X vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__buf_12
Xoutput528 _1106_/X vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__buf_12
Xoutput539 _1126_/X vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__buf_12
X_1542_ _1542_/A vssd vssd vccd vccd _1542_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1473_ _1473_/A _1473_/B vssd vssd vccd vccd _1474_/A sky130_fd_sc_hd__and2_1
XFILLER_29_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output917_A _0982_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1315__B _1315_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1331__A _1331_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1968 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1053__A_N _1309_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1225__B _1225_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_558 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input383_A la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input77_A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_779 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2190 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1416__A _1416_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1135__B _1135_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0990__A _0990_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output867_A _0946_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0973_ _0973_/A _0973_/B vssd vssd vccd vccd _0974_/A sky130_fd_sc_hd__and2_2
XFILLER_31_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1525_ _1525_/A _1525_/B vssd vssd vccd vccd _1526_/A sky130_fd_sc_hd__and2_1
XFILLER_9_1811 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1326__A _1326_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3926 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1456_ _1456_/A vssd vssd vccd vccd _1456_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1045__B _1045_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1387_ _1387_/A _1387_/B vssd vssd vccd vccd _1388_/A sky130_fd_sc_hd__and2_2
XANTENNA_user_wb_dat_gates\[26\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_716 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput870 _0896_/X vssd vssd vccd vccd mprj_adr_o_user[2] sky130_fd_sc_hd__buf_12
XANTENNA__1236__A _1236_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput881 _0576_/Y vssd vssd vccd vccd mprj_dat_i_core[0] sky130_fd_sc_hd__buf_12
Xoutput892 _0577_/Y vssd vssd vccd vccd mprj_dat_i_core[1] sky130_fd_sc_hd__buf_12
XFILLER_21_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[17\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input131_A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input229_A la_iena_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1099__A_N _1355_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0969__B _0969_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1146__A _1146_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1310_ _1310_/A vssd vssd vccd vccd _1310_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1241_ _1497_/A _1241_/B _1241_/C vssd vssd vccd vccd _1242_/A sky130_fd_sc_hd__and3b_1
XANTENNA__0985__A _0985_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_gates\[2\]_A user_irq_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output615_A _0566_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1172_ _1172_/A vssd vssd vccd vccd _1172_/X sky130_fd_sc_hd__buf_2
XFILLER_37_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0956_ _0956_/A vssd vssd vccd vccd _0956_/X sky130_fd_sc_hd__buf_6
XFILLER_50_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0887_ _0887_/A _0887_/B vssd vssd vccd vccd _0888_/A sky130_fd_sc_hd__and2_4
XFILLER_31_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0879__B _0879_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1056__A _1056_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1508_ _1508_/A vssd vssd vccd vccd _1508_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0895__A _0895_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1439_ _1439_/A _1439_/B vssd vssd vccd vccd _1440_/A sky130_fd_sc_hd__and2_2
XFILLER_22_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1241__A_N _1497_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1503__B _1503_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input179_A la_iena_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input346_A la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1413__B _1413_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0810_ _0810_/A vssd vssd vccd vccd _0810_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput13 la_data_out_mprj[108] vssd vssd vccd vccd _1235_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput24 la_data_out_mprj[118] vssd vssd vccd vccd _1255_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput35 la_data_out_mprj[12] vssd vssd vccd vccd _1043_/C sky130_fd_sc_hd__clkbuf_1
Xinput46 la_data_out_mprj[22] vssd vssd vccd vccd _1063_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_0741_ _0741_/A _0741_/B vssd vssd vccd vccd _0742_/A sky130_fd_sc_hd__and2_1
XANTENNA_output565_A _1174_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput57 la_data_out_mprj[32] vssd vssd vccd vccd _1083_/C sky130_fd_sc_hd__clkbuf_1
Xinput68 la_data_out_mprj[42] vssd vssd vccd vccd _1103_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_6_340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput79 la_data_out_mprj[52] vssd vssd vccd vccd _1123_/C sky130_fd_sc_hd__buf_2
X_0672_ _0672_/A vssd vssd vccd vccd _0672_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0699__B _0699_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output732_A _1498_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] _0762_/X vssd vssd vccd vccd _0522_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_38_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1224_ _1224_/A vssd vssd vccd vccd _1224_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1323__B _1323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1155_ _1411_/A _1155_/B _1155_/C vssd vssd vccd vccd _1156_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1086_ _1086_/A vssd vssd vccd vccd _1086_/X sky130_fd_sc_hd__buf_4
XFILLER_0_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_166 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0939_ _0939_/A _0939_/B vssd vssd vccd vccd _0940_/A sky130_fd_sc_hd__and2_2
XFILLER_28_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput406 mprj_adr_o_core[26] vssd vssd vccd vccd _0943_/B sky130_fd_sc_hd__buf_8
Xinput417 mprj_adr_o_core[7] vssd vssd vccd vccd _0905_/B sky130_fd_sc_hd__clkbuf_16
Xinput428 mprj_dat_o_core[16] vssd vssd vccd vccd _0987_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput439 mprj_dat_o_core[26] vssd vssd vccd vccd _1007_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1514__A _1514_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1233__B _1233_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1137__A_N _1393_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input296_A la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_51 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1127__C _1127_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2774 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1143__B _1143_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output947_A _0888_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0503__A _0503_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0724_ _0724_/A vssd vssd vccd vccd _0724_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0655_ _0655_/A _0655_/B vssd vssd vccd vccd _0656_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1037__C _1037_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0586_ _0586_/A vssd vssd vccd vccd _0586_/Y sky130_fd_sc_hd__inv_2
XTAP_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1334__A _1334_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1414 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1053__B _1053_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1207_ _1463_/A _1207_/B _1207_/C vssd vssd vccd vccd _1208_/A sky130_fd_sc_hd__and3b_4
XFILLER_39_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] _0814_/X vssd vssd vccd vccd _0548_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_25_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1138_ _1138_/A vssd vssd vccd vccd _1138_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_3644 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1069_ _1325_/A _1069_/B _1069_/C vssd vssd vccd vccd _1070_/A sky130_fd_sc_hd__and3b_4
XFILLER_41_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1509__A _1509_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3030 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput203 la_iena_mprj[49] vssd vssd vccd vccd _0705_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_44_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput214 la_iena_mprj[59] vssd vssd vccd vccd _0725_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_2947 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput225 la_iena_mprj[69] vssd vssd vccd vccd _0745_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_27_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput236 la_iena_mprj[79] vssd vssd vccd vccd _0765_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1244__A _1244_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput247 la_iena_mprj[89] vssd vssd vccd vccd _0785_/B sky130_fd_sc_hd__clkbuf_1
Xinput258 la_iena_mprj[99] vssd vssd vccd vccd _0805_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput269 la_oenb_mprj[108] vssd vssd vccd vccd _1491_/A sky130_fd_sc_hd__buf_2
XFILLER_2_2721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input211_A la_iena_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input309_A la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1419__A _1419_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0977__B _0977_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1154__A _1154_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0993__A _0993_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1329__A _1329_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0707_ _0707_/A _0707_/B vssd vssd vccd vccd _0708_/A sky130_fd_sc_hd__and2_1
XFILLER_45_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0887__B _0887_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0638_ _0638_/A vssd vssd vccd vccd _0638_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0569_ _0569_/A vssd vssd vccd vccd _0569_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__1064__A _1064_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1511__B _1511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4006 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1638 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1682 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input161_A la_iena_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input259_A la_iena_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input426_A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input22_A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1421__B _1421_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3850 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output478_A _1246_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput507 _1068_/X vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__buf_12
XFILLER_9_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput518 _1088_/X vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__buf_12
X_1541_ _1541_/A vssd vssd vccd vccd _1541_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__0988__A _0988_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput529 _1108_/X vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__buf_12
XANTENNA_output645_A _0478_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1472_ _1472_/A vssd vssd vccd vccd _1472_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_3080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3854 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1331__B _1331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0898__A _0898_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1225__C input8/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1241__B _1241_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input376_A la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1135__C _1135_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1151__B _1151_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0972_ _0972_/A vssd vssd vccd vccd _0972_/X sky130_fd_sc_hd__buf_6
XFILLER_35_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0511__A _0511_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1524_ _1524_/A vssd vssd vccd vccd _1524_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1823 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1455_ _1455_/A _1455_/B vssd vssd vccd vccd _1456_/A sky130_fd_sc_hd__and2_4
XFILLER_22_3938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1045__C _1045_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1386_ _1386_/A vssd vssd vccd vccd _1386_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1342__A _1342_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1061__B _1061_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1517__A _1517_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput860 _0932_/X vssd vssd vccd vccd mprj_adr_o_user[20] sky130_fd_sc_hd__buf_12
Xoutput871 _0952_/X vssd vssd vccd vccd mprj_adr_o_user[30] sky130_fd_sc_hd__buf_12
XFILLER_5_3623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput882 _0586_/Y vssd vssd vccd vccd mprj_dat_i_core[10] sky130_fd_sc_hd__buf_12
XFILLER_25_3562 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput893 _0596_/Y vssd vssd vccd vccd mprj_dat_i_core[20] sky130_fd_sc_hd__buf_12
XFILLER_5_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1252__A _1252_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input124_A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3366 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[5\] mprj_dat_i_user[5] _0870_/X vssd vssd vccd vccd _0581_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1427__A _1427_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1240_ _1240_/A vssd vssd vccd vccd _1240_/X sky130_fd_sc_hd__buf_2
XANTENNA__0985__B _0985_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output510_A _1074_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1171_ _1427_/A _1171_/B _1171_/C vssd vssd vccd vccd _1172_/A sky130_fd_sc_hd__and3b_1
XANTENNA_output608_A _0560_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1162__A _1162_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1043__A_N _1299_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] _0652_/X vssd vssd vccd vccd _0467_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_21_816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1193__A_N _1449_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0506__A _0506_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0955_ _0955_/A _0955_/B vssd vssd vccd vccd _0956_/A sky130_fd_sc_hd__and2_1
XFILLER_31_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0886_ _0886_/A vssd vssd vccd vccd _0886_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_12_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1507_ _1507_/A _1507_/B vssd vssd vccd vccd _1508_/A sky130_fd_sc_hd__and2_1
XFILLER_9_1631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1438_ _1438_/A vssd vssd vccd vccd _1438_/X sky130_fd_sc_hd__buf_2
XFILLER_9_1675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0895__B _0895_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1369_ _1369_/A _1369_/B vssd vssd vccd vccd _1370_/A sky130_fd_sc_hd__and2_2
XFILLER_20_3470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1072__A _1072_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2202 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput690 _0519_/Y vssd vssd vccd vccd la_data_in_mprj[74] sky130_fd_sc_hd__buf_12
XFILLER_40_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input241_A la_iena_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input339_A la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput14 la_data_out_mprj[109] vssd vssd vccd vccd _1237_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_32_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput25 la_data_out_mprj[119] vssd vssd vccd vccd _1257_/C sky130_fd_sc_hd__clkbuf_1
Xinput36 la_data_out_mprj[13] vssd vssd vccd vccd _1045_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_0740_ _0740_/A vssd vssd vccd vccd _0740_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput47 la_data_out_mprj[23] vssd vssd vccd vccd _1065_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_10_381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput58 la_data_out_mprj[33] vssd vssd vccd vccd _1085_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_48_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput69 la_data_out_mprj[43] vssd vssd vccd vccd _1105_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_7_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0671_ _0671_/A _0671_/B vssd vssd vccd vccd _0672_/A sky130_fd_sc_hd__and2_2
XFILLER_13_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0996__A _0996_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1223_ _1479_/A _1223_/B input7/X vssd vssd vccd vccd _1224_/A sky130_fd_sc_hd__and3b_2
XFILLER_38_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1154_ _1154_/A vssd vssd vccd vccd _1154_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1085_ _1341_/A _1085_/B _1085_/C vssd vssd vccd vccd _1086_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0938_ _0938_/A vssd vssd vccd vccd _0938_/X sky130_fd_sc_hd__buf_4
XFILLER_31_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0869_ _0869_/A _0869_/B vssd vssd vccd vccd _0870_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1089__A_N _1345_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput407 mprj_adr_o_core[27] vssd vssd vccd vccd _0945_/B sky130_fd_sc_hd__buf_8
XFILLER_6_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput418 mprj_adr_o_core[8] vssd vssd vccd vccd _0907_/B sky130_fd_sc_hd__buf_8
Xinput429 mprj_dat_o_core[17] vssd vssd vccd vccd _0989_/B sky130_fd_sc_hd__buf_2
XFILLER_44_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input191_A la_iena_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input289_A la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_63 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input456_A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input52_A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2330 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3086 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1143__C _1143_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1440__A _1440_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1231__A_N _1487_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0723_ _0723_/A _0723_/B vssd vssd vccd vccd _0724_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0654_ _0654_/A vssd vssd vccd vccd _0654_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0585_ _0585_/A vssd vssd vccd vccd _0585_/Y sky130_fd_sc_hd__inv_2
XTAP_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3902 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1206_ _1206_/A vssd vssd vccd vccd _1206_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1137_ _1393_/A _1137_/B _1137_/C vssd vssd vccd vccd _1138_/A sky130_fd_sc_hd__and3b_4
XANTENNA__1350__A _1350_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1068_ _1068_/A vssd vssd vccd vccd _1068_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_3656 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1509__B _1509_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1525__A _1525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput204 la_iena_mprj[4] vssd vssd vccd vccd _0615_/B sky130_fd_sc_hd__clkbuf_1
Xinput215 la_iena_mprj[5] vssd vssd vccd vccd _0617_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput226 la_iena_mprj[6] vssd vssd vccd vccd _0619_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_2959 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput237 la_iena_mprj[7] vssd vssd vccd vccd _0621_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput248 la_iena_mprj[8] vssd vssd vccd vccd _0623_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput259 la_iena_mprj[9] vssd vssd vccd vccd _0625_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1260__A _1260_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input204_A la_iena_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1419__B _1419_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1435__A _1435_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3990 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0993__B _0993_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output792_A _1376_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0514__A _0514_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1329__B _1329_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0706_ _0706_/A vssd vssd vccd vccd _0706_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0637_ _0637_/A _0637_/B vssd vssd vccd vccd _0638_/A sky130_fd_sc_hd__and2_1
XFILLER_48_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1345__A _1345_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0568_ _0568_/A vssd vssd vccd vccd _0568_/Y sky130_fd_sc_hd__inv_2
XTAP_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1127__A_N _1383_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0499_ _0499_/A vssd vssd vccd vccd _0499_/Y sky130_fd_sc_hd__clkinv_2
XTAP_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1080__A _1080_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1239__B _1239_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input154_A la_iena_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input321_A la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input419_A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input15_A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1149__B _1149_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput508 _1070_/X vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__buf_12
XFILLER_5_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1540_ _1540_/A vssd vssd vccd vccd _1540_/Y sky130_fd_sc_hd__clkinv_2
Xoutput519 _1090_/X vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__buf_12
XFILLER_5_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1471_ _1471_/A _1471_/B vssd vssd vccd vccd _1472_/A sky130_fd_sc_hd__and2_1
XFILLER_46_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output638_A _0472_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_ack_gate mprj_ack_i_user _0870_/X vssd vssd vccd vccd _0608_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3866 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] _0712_/X vssd vssd vccd vccd _0497_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_36_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_847 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1059__B _1059_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3952 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[29\]_A mprj_dat_i_user[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input7_A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3490 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1241__C _1241_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input271_A la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input369_A la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2818 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_954 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output490_A _1268_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0971_ _0971_/A _0971_/B vssd vssd vccd vccd _0972_/A sky130_fd_sc_hd__and2_1
XFILLER_31_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output588_A _1216_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0999__A _0999_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3755 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output922_A _0992_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1523_ _1523_/A _1523_/B vssd vssd vccd vccd _1524_/A sky130_fd_sc_hd__and2_1
XFILLER_25_3029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1454_ _1454_/A vssd vssd vccd vccd _1454_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_2569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1879 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1385_ _1385_/A _1385_/B vssd vssd vccd vccd _1386_/A sky130_fd_sc_hd__and2_4
XFILLER_3_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3674 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1061__C _1061_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_699 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1517__B _1517_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput850 _0914_/X vssd vssd vccd vccd mprj_adr_o_user[11] sky130_fd_sc_hd__buf_12
XFILLER_47_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput861 _0934_/X vssd vssd vccd vccd mprj_adr_o_user[21] sky130_fd_sc_hd__buf_12
Xoutput872 _0954_/X vssd vssd vccd vccd mprj_adr_o_user[31] sky130_fd_sc_hd__buf_12
XFILLER_5_3635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput883 _0587_/Y vssd vssd vccd vccd mprj_dat_i_core[11] sky130_fd_sc_hd__buf_12
Xoutput894 _0597_/Y vssd vssd vccd vccd mprj_dat_i_core[21] sky130_fd_sc_hd__buf_12
XFILLER_25_3574 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input117_A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input82_A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1427__B _1427_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1443__A _1443_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1170_ _1170_/A vssd vssd vccd vccd _1170_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output503_A _1060_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output872_A _0954_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[28\] mprj_dat_i_user[28] _0870_/X vssd vssd vccd vccd _0604_/A
+ sky130_fd_sc_hd__nand2_1
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] _0638_/X vssd vssd vccd vccd _1548_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_31_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0954_ _0954_/A vssd vssd vccd vccd _0954_/X sky130_fd_sc_hd__buf_4
XFILLER_50_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0885_ _0885_/A _0885_/B vssd vssd vccd vccd _0886_/A sky130_fd_sc_hd__and2_4
XANTENNA__0522__A _0522_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1337__B _1337_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1506_ _1506_/A vssd vssd vccd vccd _1506_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1437_ _1437_/A _1437_/B vssd vssd vccd vccd _1438_/A sky130_fd_sc_hd__and2_1
XFILLER_29_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] _0860_/X vssd vssd vccd vccd _0571_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_9_1687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1368_ _1368_/A vssd vssd vccd vccd _1368_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1299_ _1299_/A _1299_/B vssd vssd vccd vccd _1300_/A sky130_fd_sc_hd__and2_2
XFILLER_3_1253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2719 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1528__A _1528_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1247__B _1247_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4050 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2214 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput680 _0510_/Y vssd vssd vccd vccd la_data_in_mprj[65] sky130_fd_sc_hd__buf_12
Xoutput691 _0520_/Y vssd vssd vccd vccd la_data_in_mprj[75] sky130_fd_sc_hd__buf_12
XFILLER_43_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input234_A la_iena_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input401_A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput15 la_data_out_mprj[10] vssd vssd vccd vccd _1039_/C sky130_fd_sc_hd__clkbuf_2
Xinput26 la_data_out_mprj[11] vssd vssd vccd vccd _1041_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_32_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput37 la_data_out_mprj[14] vssd vssd vccd vccd _1047_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_6_320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1438__A _1438_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput48 la_data_out_mprj[24] vssd vssd vccd vccd _1067_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_7_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput59 la_data_out_mprj[34] vssd vssd vccd vccd _1087_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_10_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0670_ _0670_/A vssd vssd vccd vccd _0670_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1157__B _1157_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output620_A _0571_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output718_A _1542_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1222_ _1222_/A vssd vssd vccd vccd _1222_/X sky130_fd_sc_hd__buf_2
XFILLER_42_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1153_ _1409_/A _1153_/B _1153_/C vssd vssd vccd vccd _1154_/A sky130_fd_sc_hd__and3b_1
XFILLER_42_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1084_ _1084_/A vssd vssd vccd vccd _1084_/X sky130_fd_sc_hd__buf_4
XFILLER_20_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0517__A _0517_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0937_ _0937_/A _0937_/B vssd vssd vccd vccd _0938_/A sky130_fd_sc_hd__and2_1
XFILLER_48_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1348__A _1348_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0868_ _0868_/A vssd vssd vccd vccd _0868_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1067__B _1067_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0799_ _0799_/A _0799_/B vssd vssd vccd vccd _0800_/A sky130_fd_sc_hd__and2_4
XFILLER_28_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput408 mprj_adr_o_core[28] vssd vssd vccd vccd _0947_/B sky130_fd_sc_hd__buf_8
XFILLER_44_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput419 mprj_adr_o_core[9] vssd vssd vccd vccd _0909_/B sky130_fd_sc_hd__buf_4
XFILLER_9_1451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4016 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1258__A _1258_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input184_A la_iena_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1033__A_N _1289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input351_A la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input449_A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input45_A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1183__A_N _1439_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3098 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2386 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_430 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_474 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output570_A _1182_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output668_A _0499_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1168__A _1168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0722_ _0722_/A vssd vssd vccd vccd _0722_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0653_ _0653_/A _0653_/B vssd vssd vccd vccd _0654_/A sky130_fd_sc_hd__and2_1
XFILLER_45_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0800__A _0800_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0584_ _0584_/A vssd vssd vccd vccd _0584_/Y sky130_fd_sc_hd__clkinv_2
XTAP_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] _0772_/X vssd vssd vccd vccd _0527_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1205_ _1461_/A _1205_/B _1205_/C vssd vssd vccd vccd _1206_/A sky130_fd_sc_hd__and3b_4
XFILLER_4_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1136_ _1136_/A vssd vssd vccd vccd _1136_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1067_ _1323_/A _1067_/B _1067_/C vssd vssd vccd vccd _1068_/A sky130_fd_sc_hd__and3b_4
XFILLER_41_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1078__A _1078_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0710__A _0710_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1525__B _1525_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput205 la_iena_mprj[50] vssd vssd vccd vccd _0707_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput216 la_iena_mprj[60] vssd vssd vccd vccd _0727_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_41_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput227 la_iena_mprj[70] vssd vssd vccd vccd _0747_/B sky130_fd_sc_hd__buf_2
XFILLER_6_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput238 la_iena_mprj[80] vssd vssd vccd vccd _0767_/B sky130_fd_sc_hd__buf_4
XFILLER_5_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput249 la_iena_mprj[90] vssd vssd vccd vccd _0787_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input399_A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1435__B _1435_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1451__A _1451_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1079__A_N _1335_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output785_A _1364_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output952_A output952/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[10\] mprj_dat_i_user[10] _0870_/X vssd vssd vccd vccd _0586_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_30_1729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0705_ _0705_/A _0705_/B vssd vssd vccd vccd _0706_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0530__A _0530_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0636_ _0636_/A vssd vssd vccd vccd _0636_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1345__B _1345_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0567_ _0567_/A vssd vssd vccd vccd _0567_/Y sky130_fd_sc_hd__inv_2
XTAP_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0498_ _0498_/A vssd vssd vccd vccd _0498_/Y sky130_fd_sc_hd__clkinv_2
XTAP_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1361__A _1361_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ _1375_/A _1119_/B _1119_/C vssd vssd vccd vccd _1120_/A sky130_fd_sc_hd__and3b_2
XTAP_1919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0705__A _0705_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1239__C _1239_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1536__A _1536_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1255__B _1255_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input147_A la_iena_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input314_A la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1221__A_N _1477_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0615__A _0615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput509 _1072_/X vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__buf_12
XFILLER_29_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1446__A _1446_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1470_ _1470_/A vssd vssd vccd vccd _1470_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1165__B _1165_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output533_A _1116_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3878 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] _0698_/X vssd vssd vccd vccd _0490_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_47_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3616 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0525__A _0525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1059__C _1059_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1356__A _1356_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] _0622_/X vssd vssd vccd vccd _1540_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__1075__B _1075_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0619_ _0619_/A _0619_/B vssd vssd vccd vccd _0620_/A sky130_fd_sc_hd__and2_1
XANTENNA_user_wb_dat_gates\[29\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2884 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1266__A _1266_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input264_A la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input431_A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2314 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0970_ _0970_/A vssd vssd vccd vccd _0970_/X sky130_fd_sc_hd__buf_6
XFILLER_13_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output483_A _1256_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1117__A_N _1373_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0999__B _0999_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output650_A _0483_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1176__A _1176_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1522_ _1522_/A vssd vssd vccd vccd _1522_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_4045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1267__A_N _1523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_270 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output915_A _0978_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1453_ _1453_/A _1453_/B vssd vssd vccd vccd _1454_/A sky130_fd_sc_hd__and2_2
XFILLER_29_1753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1384_ _1384_/A vssd vssd vccd vccd _1384_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3090 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3686 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1086__A _1086_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput840 _1464_/X vssd vssd vccd vccd la_oenb_core[94] sky130_fd_sc_hd__buf_12
XFILLER_47_1820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput851 _0916_/X vssd vssd vccd vccd mprj_adr_o_user[12] sky130_fd_sc_hd__buf_12
XFILLER_43_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput862 _0936_/X vssd vssd vccd vccd mprj_adr_o_user[22] sky130_fd_sc_hd__buf_12
Xoutput873 _0898_/X vssd vssd vccd vccd mprj_adr_o_user[3] sky130_fd_sc_hd__buf_12
Xoutput884 _0588_/Y vssd vssd vccd vccd mprj_dat_i_core[12] sky130_fd_sc_hd__buf_12
Xoutput895 _0598_/Y vssd vssd vccd vccd mprj_dat_i_core[22] sky130_fd_sc_hd__buf_12
XFILLER_43_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2863 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input381_A la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input75_A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1443__B _1443_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output865_A _0942_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0953_ _0953_/A _0953_/B vssd vssd vccd vccd _0954_/A sky130_fd_sc_hd__and2_1
XFILLER_35_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0803__A _0803_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0884_ _0884_/A vssd vssd vccd vccd _0884_/X sky130_fd_sc_hd__buf_8
XFILLER_12_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1505_ _1505_/A _1505_/B vssd vssd vccd vccd _1506_/A sky130_fd_sc_hd__and2_1
XFILLER_47_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1436_ _1436_/A vssd vssd vccd vccd _1436_/X sky130_fd_sc_hd__buf_2
XFILLER_9_1655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1353__B _1353_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1699 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1367_ _1367_/A _1367_/B vssd vssd vccd vccd _1368_/A sky130_fd_sc_hd__and2_2
XFILLER_20_3450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] _0846_/X vssd vssd vccd vccd _0564_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_3_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1298_ _1298_/A vssd vssd vccd vccd _1298_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0713__A _0713_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1247__C _1247_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2226 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput670 _0501_/Y vssd vssd vccd vccd la_data_in_mprj[56] sky130_fd_sc_hd__buf_12
XFILLER_25_4095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput681 _0511_/Y vssd vssd vccd vccd la_data_in_mprj[66] sky130_fd_sc_hd__buf_12
XFILLER_47_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput692 _0521_/Y vssd vssd vccd vccd la_data_in_mprj[76] sky130_fd_sc_hd__buf_12
XFILLER_40_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1263__B _1263_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input227_A la_iena_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput16 la_data_out_mprj[110] vssd vssd vccd vccd _1239_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__0623__A _0623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput27 la_data_out_mprj[120] vssd vssd vccd vccd _1259_/C sky130_fd_sc_hd__clkbuf_2
Xinput38 la_data_out_mprj[15] vssd vssd vccd vccd _1049_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_32_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput49 la_data_out_mprj[25] vssd vssd vccd vccd _1069_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1157__C _1157_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1454__A _1454_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1173__B _1173_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1221_ _1477_/A _1221_/B input6/X vssd vssd vccd vccd _1222_/A sky130_fd_sc_hd__and3b_4
XFILLER_43_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1152_ _1152_/A vssd vssd vccd vccd _1152_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1083_ _1339_/A _1083_/B _1083_/C vssd vssd vccd vccd _1084_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1104 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0533__A _0533_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0936_ _0936_/A vssd vssd vccd vccd _0936_/X sky130_fd_sc_hd__buf_6
XFILLER_9_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0867_ _0867_/A _0867_/B vssd vssd vccd vccd _0868_/A sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
X_0798_ _0798_/A vssd vssd vccd vccd _0798_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1364__A _1364_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput409 mprj_adr_o_core[29] vssd vssd vccd vccd _0949_/B sky130_fd_sc_hd__buf_8
XFILLER_44_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1083__B _1083_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1419_ _1419_/A _1419_/B vssd vssd vccd vccd _1420_/A sky130_fd_sc_hd__and2_1
XFILLER_29_704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input177_A la_iena_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1274__A _1274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input344_A la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input38_A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1449__A _1449_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0721_ _0721_/A _0721_/B vssd vssd vccd vccd _0722_/A sky130_fd_sc_hd__and2_1
XANTENNA_output563_A _1170_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0652_ _0652_/A vssd vssd vccd vccd _0652_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output828_A _1442_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0583_ _0583_/A vssd vssd vccd vccd _0583_/Y sky130_fd_sc_hd__inv_2
XTAP_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] _0758_/X vssd vssd vccd vccd _0520_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1204_ _1204_/A vssd vssd vccd vccd _1204_/X sky130_fd_sc_hd__buf_2
XFILLER_39_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_718 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0528__A _0528_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1135_ _1391_/A _1135_/B _1135_/C vssd vssd vccd vccd _1136_/A sky130_fd_sc_hd__and3b_4
XFILLER_0_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1066_ _1066_/A vssd vssd vccd vccd _1066_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1359__A _1359_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0919_ _0919_/A _0919_/B vssd vssd vccd vccd _0920_/A sky130_fd_sc_hd__and2_2
XFILLER_11_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1094__A _1094_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput206 la_iena_mprj[51] vssd vssd vccd vccd _0709_/B sky130_fd_sc_hd__clkbuf_2
Xinput217 la_iena_mprj[61] vssd vssd vccd vccd _0729_/B sky130_fd_sc_hd__clkbuf_2
Xinput228 la_iena_mprj[71] vssd vssd vccd vccd _0749_/B sky130_fd_sc_hd__buf_2
XFILLER_48_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput239 la_iena_mprj[81] vssd vssd vccd vccd _0769_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_206 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input294_A la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input461_A user_irq_ena[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__0901__A _0901_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1451__B _1451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_294 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output945_A _0884_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0811__A _0811_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0704_ _0704_/A vssd vssd vccd vccd _0704_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0635_ _0635_/A _0635_/B vssd vssd vccd vccd _0636_/A sky130_fd_sc_hd__and2_1
XFILLER_25_3927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0566_ _0566_/A vssd vssd vccd vccd _0566_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0497_ _0497_/A vssd vssd vccd vccd _0497_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_39_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1361__B _1361_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] _0810_/X vssd vssd vccd vccd _0546_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA__1023__A_N _1279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1118_ _1118_/A vssd vssd vccd vccd _1118_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1049_ _1305_/A _1049_/B _1049_/C vssd vssd vccd vccd _1050_/A sky130_fd_sc_hd__and3b_4
XFILLER_41_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1173__A_N _1429_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0721__A _0721_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1255__C _1255_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1271__B _1271_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input307_A la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0631__A _0631_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1165__C _1165_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1462__A _1462_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1181__B _1181_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] _0684_/X vssd vssd vccd vccd _0483_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_36_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0806__A _0806_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0541__A _0541_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1075__C _1075_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0618_ _0618_/A vssd vssd vccd vccd _0618_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0549_ _0549_/A vssd vssd vccd vccd _0549_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__1372__A _1372_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1091__B _1091_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_802 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1069__A_N _1325_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input257_A la_iena_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1282__A _1282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input424_A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1915 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input20_A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output476_A _1242_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1457__A _1457_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[71\]_B _0750_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1521_ _1521_/A _1521_/B vssd vssd vccd vccd _1522_/A sky130_fd_sc_hd__and2_1
XANTENNA_output643_A _0476_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1452_ _1452_/A vssd vssd vccd vccd _1452_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_42_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output810_A _1410_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output908_A _0581_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1383_ _1383_/A _1383_/B vssd vssd vccd vccd _1384_/A sky130_fd_sc_hd__and2_1
XANTENNA__1192__A _1192_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0536__A _0536_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1102 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1367__A _1367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1211__A_N _1467_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput830 _1446_/X vssd vssd vccd vccd la_oenb_core[85] sky130_fd_sc_hd__buf_12
Xoutput841 _1466_/X vssd vssd vccd vccd la_oenb_core[95] sky130_fd_sc_hd__buf_12
XFILLER_25_3532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput852 _0918_/X vssd vssd vccd vccd mprj_adr_o_user[13] sky130_fd_sc_hd__buf_12
XFILLER_47_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput863 _0938_/X vssd vssd vccd vccd mprj_adr_o_user[23] sky130_fd_sc_hd__buf_12
XFILLER_5_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput874 _0900_/X vssd vssd vccd vccd mprj_adr_o_user[4] sky130_fd_sc_hd__buf_12
XFILLER_8_2037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput885 _0589_/Y vssd vssd vccd vccd mprj_dat_i_core[13] sky130_fd_sc_hd__buf_12
XFILLER_8_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput896 _0599_/Y vssd vssd vccd vccd mprj_dat_i_core[23] sky130_fd_sc_hd__buf_12
XFILLER_25_2831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1277__A _1277_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input374_A la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input68_A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_142 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0952_ _0952_/A vssd vssd vccd vccd _0952_/X sky130_fd_sc_hd__buf_4
XFILLER_31_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0883_ _0883_/A _0883_/B vssd vssd vccd vccd _0884_/A sky130_fd_sc_hd__and2_4
XFILLER_35_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output858_A _0930_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3830 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1504_ _1504_/A vssd vssd vccd vccd _1504_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1435_ _1435_/A _1435_/B vssd vssd vccd vccd _1436_/A sky130_fd_sc_hd__and2_1
XFILLER_9_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1366_ _1366_/A vssd vssd vccd vccd _1366_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1297_ _1297_/A _1297_/B vssd vssd vccd vccd _1298_/A sky130_fd_sc_hd__and2_2
XFILLER_3_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0713__B _0713_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4074 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput660 _0492_/Y vssd vssd vccd vccd la_data_in_mprj[47] sky130_fd_sc_hd__buf_12
XFILLER_40_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput671 _0502_/Y vssd vssd vccd vccd la_data_in_mprj[57] sky130_fd_sc_hd__buf_12
XFILLER_9_3592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput682 _0512_/Y vssd vssd vccd vccd la_data_in_mprj[67] sky130_fd_sc_hd__buf_12
XFILLER_21_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput693 _0522_/Y vssd vssd vccd vccd la_data_in_mprj[77] sky130_fd_sc_hd__buf_12
XFILLER_8_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input122_A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1257__A_N _1513_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0904__A _0904_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0623__B _0623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput17 la_data_out_mprj[111] vssd vssd vccd vccd _1241_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_32_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput28 la_data_out_mprj[121] vssd vssd vccd vccd _1261_/C sky130_fd_sc_hd__clkbuf_2
Xinput39 la_data_out_mprj[16] vssd vssd vccd vccd _1051_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_49_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[3\] mprj_dat_i_user[3] _0870_/X vssd vssd vccd vccd _0579_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_1363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1220_ _1220_/A vssd vssd vccd vccd _1220_/X sky130_fd_sc_hd__buf_2
XANTENNA__1173__C _1173_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1151_ _1407_/A _1151_/B _1151_/C vssd vssd vccd vccd _1152_/A sky130_fd_sc_hd__and3b_2
XFILLER_42_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output606_A _0558_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1470__A _1470_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1082_ _1082_/A vssd vssd vccd vccd _1082_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] _0648_/X vssd vssd vccd vccd _0465_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_15_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0814__A _0814_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0935_ _0935_/A _0935_/B vssd vssd vccd vccd _0936_/A sky130_fd_sc_hd__and2_1
XFILLER_31_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0866_ _0866_/A vssd vssd vccd vccd _0866_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[101\]_B _0810_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0797_ _0797_/A _0797_/B vssd vssd vccd vccd _0798_/A sky130_fd_sc_hd__and2_4
XFILLER_48_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1083__C _1083_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1418_ _1418_/A vssd vssd vccd vccd _1418_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1475 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1349_ _1349_/A _1349_/B vssd vssd vccd vccd _1350_/A sky130_fd_sc_hd__and2_2
XANTENNA__1380__A _1380_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[10\]_A mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput490 _1268_/X vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__buf_12
XFILLER_43_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input337_A la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1290__A _1290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1449__B _1449_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0720_ _0720_/A vssd vssd vccd vccd _0720_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0651_ _0651_/A _0651_/B vssd vssd vccd vccd _0652_/A sky130_fd_sc_hd__and2_1
XANTENNA_output556_A _1158_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1465__A _1465_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0582_ _0582_/A vssd vssd vccd vccd _0582_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output723_A _1482_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1203_ _1459_/A _1203_/B _1203_/C vssd vssd vccd vccd _1204_/A sky130_fd_sc_hd__and3b_4
XFILLER_38_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] _0744_/X vssd vssd vccd vccd _0513_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__0809__A _0809_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1134_ _1134_/A vssd vssd vccd vccd _1134_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1065_ _1321_/A _1065_/B _1065_/C vssd vssd vccd vccd _1066_/A sky130_fd_sc_hd__and3b_2
XFILLER_52_3539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0544__A _0544_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1359__B _1359_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0918_ _0918_/A vssd vssd vccd vccd _0918_/X sky130_fd_sc_hd__buf_4
XFILLER_50_1894 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0849_ _0849_/A _0849_/B vssd vssd vccd vccd _0850_/A sky130_fd_sc_hd__and2_1
XFILLER_11_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1375__A _1375_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput207 la_iena_mprj[52] vssd vssd vccd vccd _0711_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput218 la_iena_mprj[62] vssd vssd vccd vccd _0731_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput229 la_iena_mprj[72] vssd vssd vccd vccd _0751_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0719__A _0719_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1269__B _1269_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input287_A la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0901__B _0901_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1285__A _1285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input454_A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input50_A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0629__A _0629_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1179__B _1179_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1266 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0703_ _0703_/A _0703_/B vssd vssd vccd vccd _0704_/A sky130_fd_sc_hd__and2_1
XANTENNA__0811__B _0811_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output938_A _0962_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0634_ _0634_/A vssd vssd vccd vccd _0634_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0565_ _0565_/A vssd vssd vccd vccd _0565_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_28_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0496_ _0496_/A vssd vssd vccd vccd _0496_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0539__A _0539_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1117_ _1373_/A _1117_/B _1117_/C vssd vssd vccd vccd _1118_/A sky130_fd_sc_hd__and3b_2
XFILLER_1_2791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1048_ _1048_/A vssd vssd vccd vccd _1048_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_2023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1089__B _1089_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0721__B _0721_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1271__C _1271_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input202_A la_iena_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input98_A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0912__A _0912_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1947 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3814 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output519_A _1090_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1181__C _1181_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output790_A _1374_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0617_ _0617_/A _0617_/B vssd vssd vccd vccd _0618_/A sky130_fd_sc_hd__and2_1
XFILLER_9_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[2\]_A mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0548_ _0548_/A vssd vssd vccd vccd _0548_/Y sky130_fd_sc_hd__inv_2
XTAP_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0479_ _0479_/A vssd vssd vccd vccd _0479_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_814 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input152_A la_iena_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input417_A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0907__A _0907_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_891 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1457__B _1457_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output469_A _1230_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1520_ _1520_/A vssd vssd vccd vccd _1520_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1451_ _1451_/A _1451_/B vssd vssd vccd vccd _1452_/A sky130_fd_sc_hd__and2_1
XFILLER_45_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output636_A _0470_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1473__A _1473_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1382_ _1382_/A vssd vssd vccd vccd _1382_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output803_A _1396_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1163__A_N _1419_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput390 mprj_adr_o_core[11] vssd vssd vccd vccd _0913_/B sky130_fd_sc_hd__clkbuf_4
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] _0708_/X vssd vssd vccd vccd _0495_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__0817__A _0817_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0552__A _0552_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1367__B _1367_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput820 _1428_/X vssd vssd vccd vccd la_oenb_core[76] sky130_fd_sc_hd__buf_12
XFILLER_47_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput831 _1448_/X vssd vssd vccd vccd la_oenb_core[86] sky130_fd_sc_hd__buf_12
XFILLER_9_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput842 _1468_/X vssd vssd vccd vccd la_oenb_core[96] sky130_fd_sc_hd__buf_12
Xoutput853 _0920_/X vssd vssd vccd vccd mprj_adr_o_user[14] sky130_fd_sc_hd__buf_12
Xoutput864 _0940_/X vssd vssd vccd vccd mprj_adr_o_user[24] sky130_fd_sc_hd__buf_12
XFILLER_43_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1383__A _1383_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput875 _0902_/X vssd vssd vccd vccd mprj_adr_o_user[5] sky130_fd_sc_hd__buf_12
XFILLER_9_3796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput886 _0590_/Y vssd vssd vccd vccd mprj_dat_i_core[14] sky130_fd_sc_hd__buf_12
Xoutput897 _0600_/Y vssd vssd vccd vccd mprj_dat_i_core[24] sky130_fd_sc_hd__buf_12
XFILLER_5_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input5_A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0727__A _0727_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1277__B _1277_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input367_A la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_irq_gates\[2\] user_irq_core[2] _0868_/X vssd vssd vccd vccd _0575_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1293__A _1293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0637__A _0637_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0951_ _0951_/A _0951_/B vssd vssd vccd vccd _0952_/A sky130_fd_sc_hd__and2_1
XANTENNA_output586_A _1212_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0882_ _0882_/A vssd vssd vccd vccd _0882_/X sky130_fd_sc_hd__buf_8
XFILLER_31_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1187__B _1187_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output920_A _0988_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] _0804_/X vssd vssd vccd vccd _0543_/A
+ sky130_fd_sc_hd__nand2_4
X_1503_ _1503_/A _1503_/B vssd vssd vccd vccd _1504_/A sky130_fd_sc_hd__and2_1
XFILLER_29_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1434_ _1434_/A vssd vssd vccd vccd _1434_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1365_ _1365_/A _1365_/B vssd vssd vccd vccd _1366_/A sky130_fd_sc_hd__and2_1
XFILLER_29_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1296_ _1296_/A vssd vssd vccd vccd _1296_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0547__A _0547_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1059__A_N _1315_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1378__A _1378_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1097__B _1097_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput650 _0483_/Y vssd vssd vccd vccd la_data_in_mprj[38] sky130_fd_sc_hd__buf_12
XFILLER_44_3964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput661 _0493_/Y vssd vssd vccd vccd la_data_in_mprj[48] sky130_fd_sc_hd__buf_12
XFILLER_9_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput672 _0503_/Y vssd vssd vccd vccd la_data_in_mprj[58] sky130_fd_sc_hd__buf_12
Xoutput683 _0513_/Y vssd vssd vccd vccd la_data_in_mprj[68] sky130_fd_sc_hd__buf_12
XFILLER_40_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput694 _0523_/Y vssd vssd vccd vccd la_data_in_mprj[78] sky130_fd_sc_hd__buf_12
XFILLER_8_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_986 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input115_A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1288__A _1288_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput18 la_data_out_mprj[112] vssd vssd vccd vccd _1243_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input80_A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput29 la_data_out_mprj[122] vssd vssd vccd vccd _1263_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_10_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3654 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0920__A _0920_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1162 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1150_ _1150_/A vssd vssd vccd vccd _1150_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output501_A _1058_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1081_ _1337_/A _1081_/B _1081_/C vssd vssd vccd vccd _1082_/A sky130_fd_sc_hd__and3b_1
XFILLER_37_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1201__A_N _1457_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output870_A _0896_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] _0634_/X vssd vssd vccd vccd _1546_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__1198__A _1198_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[26\] mprj_dat_i_user[26] _0870_/X vssd vssd vccd vccd _0602_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_31_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0934_ _0934_/A vssd vssd vccd vccd _0934_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0865_ _0865_/A _0865_/B vssd vssd vccd vccd _0866_/A sky130_fd_sc_hd__and2_1
XFILLER_48_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0796_ _0796_/A vssd vssd vccd vccd _0796_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1417_ _1417_/A _1417_/B vssd vssd vccd vccd _1418_/A sky130_fd_sc_hd__and2_1
XFILLER_0_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] _0856_/X vssd vssd vccd vccd _0569_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_42_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1348_ _1348_/A vssd vssd vccd vccd _1348_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1279_ _1279_/A _1279_/B vssd vssd vccd vccd _1280_/A sky130_fd_sc_hd__and2_2
XFILLER_0_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_934 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[10\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_67 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_89 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput480 _1250_/X vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__buf_12
Xoutput491 _1270_/X vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__buf_12
XFILLER_40_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input232_A la_iena_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1751 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0650_ _0650_/A vssd vssd vccd vccd _0650_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1465__B _1465_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0581_ _0581_/A vssd vssd vccd vccd _0581_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_49_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1481__A _1481_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1202_ _1202_/A vssd vssd vccd vccd _1202_/X sky130_fd_sc_hd__buf_2
XFILLER_1_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0809__B _0809_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1133_ _1389_/A _1133_/B _1133_/C vssd vssd vccd vccd _1134_/A sky130_fd_sc_hd__and3b_4
XFILLER_19_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1064_ _1064_/A vssd vssd vccd vccd _1064_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0825__A _0825_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1050 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0917_ _0917_/A _0917_/B vssd vssd vccd vccd _0918_/A sky130_fd_sc_hd__and2_1
X_0848_ _0848_/A vssd vssd vccd vccd _0848_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1375__B _1375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0779_ _0779_/A _0779_/B vssd vssd vccd vccd _0780_/A sky130_fd_sc_hd__and2_4
XFILLER_44_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1247__A_N _1503_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2919 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput208 la_iena_mprj[53] vssd vssd vccd vccd _0713_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_4078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput219 la_iena_mprj[63] vssd vssd vccd vccd _0733_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1251 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1391__A _1391_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0719__B _0719_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2654 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0735__A _0735_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1269__C _1269_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input182_A la_iena_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1285__B _1285_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input447_A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input43_A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0629__B _0629_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0645__A _0645_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1179__C _1179_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output666_A _0497_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0702_ _0702_/A vssd vssd vccd vccd _0702_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1195__B _1195_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output833_A _1452_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0633_ _0633_/A _0633_/B vssd vssd vccd vccd _0634_/A sky130_fd_sc_hd__and2_1
XFILLER_25_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0564_ _0564_/A vssd vssd vccd vccd _0564_/Y sky130_fd_sc_hd__clkinv_2
XTAP_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] _0768_/X vssd vssd vccd vccd _0525_/A
+ sky130_fd_sc_hd__nand2_8
XTAP_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1330 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0495_ _0495_/A vssd vssd vccd vccd _0495_/Y sky130_fd_sc_hd__clkinv_2
XTAP_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1116_ _1116_/A vssd vssd vccd vccd _1116_/X sky130_fd_sc_hd__buf_2
XFILLER_17_3402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0555__A _0555_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1047_ _1303_/A _1047_/B _1047_/C vssd vssd vccd vccd _1048_/A sky130_fd_sc_hd__and3b_4
XFILLER_39_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1089__C _1089_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1386__A _1386_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input397_A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1296__A _1296_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3744 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output783_A _1360_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output950_A _0882_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0616_ _0616_/A vssd vssd vccd vccd _0616_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[2\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0547_ _0547_/A vssd vssd vccd vccd _0547_/Y sky130_fd_sc_hd__inv_2
XTAP_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0478_ _0478_/A vssd vssd vccd vccd _0478_/Y sky130_fd_sc_hd__inv_2
XTAP_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_826 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input145_A la_iena_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input312_A la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0907__B _0907_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0923__A _0923_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1450_ _1450_/A vssd vssd vccd vccd _1450_/X sky130_fd_sc_hd__buf_2
XFILLER_42_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1473__B _1473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output531_A _1112_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1381_ _1381_/A _1381_/B vssd vssd vccd vccd _1382_/A sky130_fd_sc_hd__and2_4
XANTENNA_output629_A _0464_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput380 la_oenb_mprj[93] vssd vssd vccd vccd _1461_/A sky130_fd_sc_hd__buf_2
XFILLER_36_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput391 mprj_adr_o_core[12] vssd vssd vccd vccd _0915_/B sky130_fd_sc_hd__buf_6
XFILLER_23_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] _0694_/X vssd vssd vccd vccd _0488_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_18_3530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0833__A _0833_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput810 _1410_/X vssd vssd vccd vccd la_oenb_core[67] sky130_fd_sc_hd__buf_12
Xoutput821 _1430_/X vssd vssd vccd vccd la_oenb_core[77] sky130_fd_sc_hd__buf_12
Xoutput832 _1450_/X vssd vssd vccd vccd la_oenb_core[87] sky130_fd_sc_hd__buf_12
XFILLER_47_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput843 _1470_/X vssd vssd vccd vccd la_oenb_core[97] sky130_fd_sc_hd__buf_12
XFILLER_9_3764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput854 _0922_/X vssd vssd vccd vccd mprj_adr_o_user[15] sky130_fd_sc_hd__buf_12
Xoutput865 _0942_/X vssd vssd vccd vccd mprj_adr_o_user[25] sky130_fd_sc_hd__buf_12
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] _0618_/X vssd vssd vccd vccd _1538_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput876 _0904_/X vssd vssd vccd vccd mprj_adr_o_user[6] sky130_fd_sc_hd__buf_12
XFILLER_8_2039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1383__B _1383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput887 _0591_/Y vssd vssd vccd vccd mprj_dat_i_core[15] sky130_fd_sc_hd__buf_12
XFILLER_28_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput898 _0601_/Y vssd vssd vccd vccd mprj_dat_i_core[25] sky130_fd_sc_hd__buf_12
XTAP_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0727__B _0727_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_41_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input262_A la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1293__B _1293_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0918__A _0918_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0637__B _0637_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0653__A _0653_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0950_ _0950_/A vssd vssd vccd vccd _0950_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output481_A _1252_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0881_ _0881_/A _0881_/B vssd vssd vccd vccd _0882_/A sky130_fd_sc_hd__and2_2
XANTENNA_output579_A _1036_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1187__C _1187_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1502_ _1502_/A vssd vssd vccd vccd _1502_/X sky130_fd_sc_hd__buf_2
XFILLER_47_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output913_A _0956_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1433_ _1433_/A _1433_/B vssd vssd vccd vccd _1434_/A sky130_fd_sc_hd__and2_1
X_1364_ _1364_/A vssd vssd vccd vccd _1364_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0828__A _0828_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1295_ _1295_/A _1295_/B vssd vssd vccd vccd _1296_/A sky130_fd_sc_hd__and2_4
XFILLER_0_3547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1394__A _1394_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput640 _0474_/Y vssd vssd vccd vccd la_data_in_mprj[29] sky130_fd_sc_hd__buf_12
XFILLER_47_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput651 _0484_/Y vssd vssd vccd vccd la_data_in_mprj[39] sky130_fd_sc_hd__buf_12
Xoutput662 _0494_/Y vssd vssd vccd vccd la_data_in_mprj[49] sky130_fd_sc_hd__buf_12
Xoutput673 _0504_/Y vssd vssd vccd vccd la_data_in_mprj[59] sky130_fd_sc_hd__buf_12
Xoutput684 _0514_/Y vssd vssd vccd vccd la_data_in_mprj[69] sky130_fd_sc_hd__buf_12
Xoutput695 _0524_/Y vssd vssd vccd vccd la_data_in_mprj[79] sky130_fd_sc_hd__buf_12
XFILLER_40_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2674 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input108_A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1153__A_N _1409_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput19 la_data_out_mprj[113] vssd vssd vccd vccd _1245_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_32_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input73_A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3139 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1080_ _1080_/A vssd vssd vccd vccd _1080_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output696_A _1540_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1479__A _1479_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0933_ _0933_/A _0933_/B vssd vssd vccd vccd _0934_/A sky130_fd_sc_hd__and2_1
XANTENNA_output863_A _0938_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[19\] mprj_dat_i_user[19] _0870_/X vssd vssd vccd vccd _0595_/A
+ sky130_fd_sc_hd__nand2_2
X_0864_ _0864_/A vssd vssd vccd vccd _0864_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0795_ _0795_/A _0795_/B vssd vssd vccd vccd _0796_/A sky130_fd_sc_hd__and2_4
XFILLER_28_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1416_ _1416_/A vssd vssd vccd vccd _1416_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1347_ _1347_/A _1347_/B vssd vssd vccd vccd _1348_/A sky130_fd_sc_hd__and2_2
XFILLER_29_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] _0842_/X vssd vssd vccd vccd _0562_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_3_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1278_ _1278_/A vssd vssd vccd vccd _1278_/X sky130_fd_sc_hd__buf_2
XFILLER_25_902 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1389__A _1389_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3931 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput470 _1232_/X vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__buf_12
XFILLER_44_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput481 _1252_/X vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__buf_12
Xoutput492 _1272_/X vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__buf_12
XFILLER_40_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input225_A la_iena_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0915__B _0915_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1299__A _1299_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0931__A _0931_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0580_ _0580_/A vssd vssd vccd vccd _0580_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1049__A_N _1305_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1481__B _1481_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1201_ _1457_/A _1201_/B _1201_/C vssd vssd vccd vccd _1202_/A sky130_fd_sc_hd__and3b_4
XANTENNA_output611_A _0563_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output709_A _0536_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1132_ _1132_/A vssd vssd vccd vccd _1132_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_1122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1199__A_N _1455_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1063_ _1319_/A _1063_/B _1063_/C vssd vssd vccd vccd _1064_/A sky130_fd_sc_hd__and3b_4
XFILLER_17_3606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0825__B _0825_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4064 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1002__A _1002_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0841__A _0841_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0916_ _0916_/A vssd vssd vccd vccd _0916_/X sky130_fd_sc_hd__buf_4
XFILLER_50_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0847_ _0847_/A _0847_/B vssd vssd vccd vccd _0848_/A sky130_fd_sc_hd__and2_1
XFILLER_44_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0778_ _0778_/A vssd vssd vccd vccd _0778_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput209 la_iena_mprj[54] vssd vssd vccd vccd _0715_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1391__B _1391_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0735__B _0735_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0751__A _0751_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input175_A la_iena_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input342_A la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input36_A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0926__A _0926_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0645__B _0645_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0661__A _0661_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0701_ _0701_/A _0701_/B vssd vssd vccd vccd _0702_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output659_A _0491_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0632_ _0632_/A vssd vssd vccd vccd _0632_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1195__C _1195_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0563_ _0563_/A vssd vssd vccd vccd _0563_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output826_A _1438_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0494_ _0494_/A vssd vssd vccd vccd _0494_/Y sky130_fd_sc_hd__inv_2
XTAP_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1342 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] _0754_/X vssd vssd vccd vccd _0518_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1115_ _1371_/A _1115_/B _1115_/C vssd vssd vccd vccd _1116_/A sky130_fd_sc_hd__and3b_2
XANTENNA__0836__A _0836_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1046_ _1046_/A vssd vssd vccd vccd _1046_/X sky130_fd_sc_hd__buf_2
XFILLER_22_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1758 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2430 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0746__A _0746_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__0481__A _0481_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input292_A la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_978 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3756 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1237__A_N _1493_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output776_A _1348_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1487__A _1487_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output943_A _0972_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0615_ _0615_/A _0615_/B vssd vssd vccd vccd _0616_/A sky130_fd_sc_hd__and2_1
XFILLER_41_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0546_ _0546_/A vssd vssd vccd vccd _0546_/Y sky130_fd_sc_hd__inv_2
XTAP_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0477_ _0477_/A vssd vssd vccd vccd _0477_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_1029_ _1285_/A _1029_/B _1029_/C vssd vssd vccd vccd _1030_/A sky130_fd_sc_hd__and3b_1
XFILLER_41_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1397__A _1397_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3478 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1294 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input138_A la_iena_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0476__A _0476_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input305_A la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0923__B _0923_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_B _0720_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1100__A _1100_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_90 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1380_ _1380_/A vssd vssd vccd vccd _1380_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_3602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output524_A _1026_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput370 la_oenb_mprj[84] vssd vssd vccd vccd _1443_/A sky130_fd_sc_hd__buf_4
XFILLER_3_1417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput381 la_oenb_mprj[94] vssd vssd vccd vccd _1463_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput392 mprj_adr_o_core[13] vssd vssd vccd vccd _0917_/B sky130_fd_sc_hd__buf_6
XFILLER_36_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] _0680_/X vssd vssd vccd vccd _0481_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0833__B _0833_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1010__A _1010_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput800 _1392_/X vssd vssd vccd vccd la_oenb_core[58] sky130_fd_sc_hd__buf_12
Xoutput811 _1412_/X vssd vssd vccd vccd la_oenb_core[68] sky130_fd_sc_hd__buf_12
Xoutput822 _1432_/X vssd vssd vccd vccd la_oenb_core[78] sky130_fd_sc_hd__buf_12
Xoutput833 _1452_/X vssd vssd vccd vccd la_oenb_core[88] sky130_fd_sc_hd__buf_12
Xoutput844 _1472_/X vssd vssd vccd vccd la_oenb_core[98] sky130_fd_sc_hd__buf_12
XFILLER_8_2007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput855 _0924_/X vssd vssd vccd vccd mprj_adr_o_user[16] sky130_fd_sc_hd__buf_12
XFILLER_47_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput866 _0944_/X vssd vssd vccd vccd mprj_adr_o_user[26] sky130_fd_sc_hd__buf_12
XFILLER_29_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput877 _0906_/X vssd vssd vccd vccd mprj_adr_o_user[7] sky130_fd_sc_hd__buf_12
XFILLER_5_3629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput888 _0592_/Y vssd vssd vccd vccd mprj_dat_i_core[16] sky130_fd_sc_hd__buf_12
XFILLER_28_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput899 _0602_/Y vssd vssd vccd vccd mprj_dat_i_core[26] sky130_fd_sc_hd__buf_12
XTAP_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0529_ _0529_/A vssd vssd vccd vccd _0529_/Y sky130_fd_sc_hd__inv_2
XTAP_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2146 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0743__B _0743_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input255_A la_iena_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input422_A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[31\]_A mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0934__A _0934_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0653__B _0653_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0880_ _0880_/A vssd vssd vccd vccd _0880_/X sky130_fd_sc_hd__buf_8
XFILLER_16_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output474_A _1040_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1501_ _1501_/A _1501_/B vssd vssd vccd vccd _1502_/A sky130_fd_sc_hd__and2_1
XFILLER_42_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output739_A _1512_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1432_ _1432_/A vssd vssd vccd vccd _1432_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1363_ _1363_/A _1363_/B vssd vssd vccd vccd _1364_/A sky130_fd_sc_hd__and2_2
XANTENNA_output906_A _0579_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1294_ _1294_/A vssd vssd vccd vccd _1294_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_3695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1142 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1005__A _1005_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_A mprj_dat_i_user[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0844__A _0844_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3258 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[104\]_B _0816_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput630 _1534_/Y vssd vssd vccd vccd la_data_in_mprj[1] sky130_fd_sc_hd__buf_12
Xoutput641 _1535_/Y vssd vssd vccd vccd la_data_in_mprj[2] sky130_fd_sc_hd__buf_12
XFILLER_5_3404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput652 _1536_/Y vssd vssd vccd vccd la_data_in_mprj[3] sky130_fd_sc_hd__buf_12
XFILLER_47_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput663 _1537_/Y vssd vssd vccd vccd la_data_in_mprj[4] sky130_fd_sc_hd__buf_12
XFILLER_9_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput674 _1538_/Y vssd vssd vccd vccd la_data_in_mprj[5] sky130_fd_sc_hd__buf_12
XFILLER_28_1020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput685 _1539_/Y vssd vssd vccd vccd la_data_in_mprj[6] sky130_fd_sc_hd__buf_12
Xoutput696 _1540_/Y vssd vssd vccd vccd la_data_in_mprj[7] sky130_fd_sc_hd__buf_12
XFILLER_5_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1242 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[13\]_A mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1770 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0754__A _0754_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input372_A la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input66_A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0929__A _0929_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1479__B _1479_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output689_A _0518_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0932_ _0932_/A vssd vssd vccd vccd _0932_/X sky130_fd_sc_hd__buf_4
XFILLER_53_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output856_A _0926_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0863_ _0863_/A _0863_/B vssd vssd vccd vccd _0864_/A sky130_fd_sc_hd__and2_1
XANTENNA__1495__A _1495_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0794_ _0794_/A vssd vssd vccd vccd _0794_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1415_ _1415_/A _1415_/B vssd vssd vccd vccd _1416_/A sky130_fd_sc_hd__and2_1
XFILLER_6_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0839__A _0839_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1346_ _1346_/A vssd vssd vccd vccd _1346_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_1259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1277_ _1277_/A _1277_/B vssd vssd vccd vccd _1278_/A sky130_fd_sc_hd__and2_2
XFILLER_37_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1389__B _1389_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput471 _1234_/X vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__buf_12
Xoutput482 _1254_/X vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__buf_12
Xoutput493 _1274_/X vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__buf_12
XFILLER_5_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0749__A _0749_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input120_A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input218_A la_iena_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0484__A _0484_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1299__B _1299_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0931__B _0931_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[1\] mprj_dat_i_user[1] _0870_/X vssd vssd vccd vccd _0577_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0659__A _0659_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1200_ _1200_/A vssd vssd vccd vccd _1200_/X sky130_fd_sc_hd__buf_2
X_1131_ _1387_/A _1131_/B _1131_/C vssd vssd vccd vccd _1132_/A sky130_fd_sc_hd__and3b_4
XANTENNA_output604_A _0556_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1062_ _1062_/A vssd vssd vccd vccd _1062_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[31\] mprj_dat_i_user[31] _0870_/X vssd vssd vccd vccd _0607_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_15_980 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1074 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0915_ _0915_/A _0915_/B vssd vssd vccd vccd _0916_/A sky130_fd_sc_hd__and2_1
XFILLER_11_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0841__B _0841_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0846_ _0846_/A vssd vssd vccd vccd _0846_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0777_ _0777_/A _0777_/B vssd vssd vccd vccd _0778_/A sky130_fd_sc_hd__and2_4
XFILLER_48_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1143__A_N _1399_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1329_ _1329_/A _1329_/B vssd vssd vccd vccd _1330_/A sky130_fd_sc_hd__and2_2
XFILLER_39_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_744 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0751__B _0751_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input168_A la_iena_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0479__A _0479_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input335_A la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input29_A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0942__A _0942_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0661__B _0661_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0700_ _0700_/A vssd vssd vccd vccd _0700_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0631_ _0631_/A _0631_/B vssd vssd vccd vccd _0632_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output554_A _1154_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0562_ _0562_/A vssd vssd vccd vccd _0562_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output721_A _1478_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0493_ _0493_/A vssd vssd vccd vccd _0493_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1354 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] _0740_/X vssd vssd vccd vccd _0511_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_39_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1114_ _1114_/A vssd vssd vccd vccd _1114_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_2750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1045_ _1301_/A _1045_/B _1045_/C vssd vssd vccd vccd _1046_/A sky130_fd_sc_hd__and3b_2
XFILLER_52_3317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1013__A _1013_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0829_ _0829_/A _0829_/B vssd vssd vccd vccd _0830_/A sky130_fd_sc_hd__and2_1
XANTENNA_user_wb_dat_gates\[5\]_A mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1083 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0762__A _0762_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1039__A_N _1295_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input285_A la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1870 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1189__A_N _1445_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input452_A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1863 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0672__A _0672_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1487__B _1487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output671_A _0502_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output769_A _1280_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output936_A _1016_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0614_ _0614_/A vssd vssd vccd vccd _0614_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0545_ _0545_/A vssd vssd vccd vccd _0545_/Y sky130_fd_sc_hd__inv_2
XTAP_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1008__A _1008_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0476_ _0476_/A vssd vssd vccd vccd _0476_/Y sky130_fd_sc_hd__clkinv_2
XTAP_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0847__A _0847_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1028_ _1028_/A vssd vssd vccd vccd _1028_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1397__B _1397_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0757__A _0757_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input200_A la_iena_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0492__A _0492_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input96_A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0667__A _0667_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output517_A _1086_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput360 la_oenb_mprj[75] vssd vssd vccd vccd _1425_/A sky130_fd_sc_hd__clkbuf_4
Xinput371 la_oenb_mprj[85] vssd vssd vccd vccd _1445_/A sky130_fd_sc_hd__buf_4
XFILLER_23_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput382 la_oenb_mprj[95] vssd vssd vccd vccd _1465_/A sky130_fd_sc_hd__buf_2
XFILLER_2_3590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput393 mprj_adr_o_core[14] vssd vssd vccd vccd _0919_/B sky130_fd_sc_hd__buf_4
XFILLER_36_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] _0666_/X vssd vssd vccd vccd _0474_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_31_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput801 _1394_/X vssd vssd vccd vccd la_oenb_core[59] sky130_fd_sc_hd__buf_12
Xoutput812 _1414_/X vssd vssd vccd vccd la_oenb_core[69] sky130_fd_sc_hd__buf_12
Xoutput823 _1434_/X vssd vssd vccd vccd la_oenb_core[79] sky130_fd_sc_hd__buf_12
Xoutput834 _1454_/X vssd vssd vccd vccd la_oenb_core[89] sky130_fd_sc_hd__buf_12
XFILLER_47_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput845 _1474_/X vssd vssd vccd vccd la_oenb_core[99] sky130_fd_sc_hd__buf_12
Xoutput856 _0926_/X vssd vssd vccd vccd mprj_adr_o_user[17] sky130_fd_sc_hd__buf_12
XFILLER_8_2019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput867 _0946_/X vssd vssd vccd vccd mprj_adr_o_user[27] sky130_fd_sc_hd__buf_12
Xoutput878 _0908_/X vssd vssd vccd vccd mprj_adr_o_user[8] sky130_fd_sc_hd__buf_12
XFILLER_29_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput889 _0593_/Y vssd vssd vccd vccd mprj_dat_i_core[17] sky130_fd_sc_hd__buf_12
XFILLER_3_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0528_ _0528_/A vssd vssd vccd vccd _0528_/Y sky130_fd_sc_hd__inv_2
XTAP_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0871__A_N input3/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3772 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input150_A la_iena_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1227__A_N _1483_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input248_A la_iena_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0487__A _0487_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input415_A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input11_A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[31\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output467_A _1226_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1500_ _1500_/A vssd vssd vccd vccd _1500_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1431_ _1431_/A _1431_/B vssd vssd vccd vccd _1432_/A sky130_fd_sc_hd__and2_1
XANTENNA_output634_A _0468_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1362_ _1362_/A vssd vssd vccd vccd _1362_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1293_ _1293_/A _1293_/B vssd vssd vccd vccd _1294_/A sky130_fd_sc_hd__and2_4
XFILLER_23_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput190 la_iena_mprj[37] vssd vssd vccd vccd _0681_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1005__B _1005_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput620 _0571_/Y vssd vssd vccd vccd la_data_in_mprj[126] sky130_fd_sc_hd__buf_12
XFILLER_47_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput631 _0465_/Y vssd vssd vccd vccd la_data_in_mprj[20] sky130_fd_sc_hd__buf_12
XFILLER_9_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2919 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput642 _0475_/Y vssd vssd vccd vccd la_data_in_mprj[30] sky130_fd_sc_hd__buf_12
Xoutput653 _0485_/Y vssd vssd vccd vccd la_data_in_mprj[40] sky130_fd_sc_hd__buf_12
XFILLER_47_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput664 _0495_/Y vssd vssd vccd vccd la_data_in_mprj[50] sky130_fd_sc_hd__buf_12
XFILLER_44_3978 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput675 _0505_/Y vssd vssd vccd vccd la_data_in_mprj[60] sky130_fd_sc_hd__buf_12
XFILLER_9_3596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput686 _0515_/Y vssd vssd vccd vccd la_data_in_mprj[70] sky130_fd_sc_hd__buf_12
Xoutput697 _0525_/Y vssd vssd vccd vccd la_data_in_mprj[80] sky130_fd_sc_hd__buf_12
XFILLER_28_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input3_A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[13\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0770__A _0770_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input198_A la_iena_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input365_A la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_irq_gates\[0\] user_irq_core[0] _0864_/X vssd vssd vccd vccd _0573_/A sky130_fd_sc_hd__nand2_1
XANTENNA_input59_A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0929__B _0929_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1671 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1106__A _1106_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0945__A _0945_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1835 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ _0931_/A _0931_/B vssd vssd vccd vccd _0932_/A sky130_fd_sc_hd__and2_1
XANTENNA_output584_A _1208_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0680__A _0680_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0862_ _0862_/A vssd vssd vccd vccd _0862_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1495__B _1495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output849_A _0912_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0793_ _0793_/A _0793_/B vssd vssd vccd vccd _0794_/A sky130_fd_sc_hd__and2_4
XFILLER_44_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] _0800_/X vssd vssd vccd vccd _0541_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_6_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1414_ _1414_/A vssd vssd vccd vccd _1414_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0839__B _0839_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1345_ _1345_/A _1345_/B vssd vssd vccd vccd _1346_/A sky130_fd_sc_hd__and2_1
XANTENNA__1016__A _1016_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1276_ _1276_/A vssd vssd vccd vccd _1276_/X sky130_fd_sc_hd__buf_2
XFILLER_20_2540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0855__A _0855_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput472 _1236_/X vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__buf_12
XFILLER_47_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput483 _1256_/X vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__buf_12
Xoutput494 _1044_/X vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__buf_12
XFILLER_5_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2670 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0749__B _0749_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0765__A _0765_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input113_A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3708 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0659__B _0659_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1130_ _1130_/A vssd vssd vccd vccd _1130_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1061_ _1317_/A _1061_/B _1061_/C vssd vssd vccd vccd _1062_/A sky130_fd_sc_hd__and3b_4
XANTENNA__0675__A _0675_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1095__A_N _1351_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] _0630_/X vssd vssd vccd vccd _1544_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_50_2533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[24\] mprj_dat_i_user[24] _0870_/X vssd vssd vccd vccd _0600_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_15_3398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0914_ _0914_/A vssd vssd vccd vccd _0914_/X sky130_fd_sc_hd__buf_6
XFILLER_50_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0845_ _0845_/A _0845_/B vssd vssd vccd vccd _0846_/A sky130_fd_sc_hd__and2_1
XFILLER_11_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0776_ _0776_/A vssd vssd vccd vccd _0776_/X sky130_fd_sc_hd__buf_2
XFILLER_22_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1046 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] _0852_/X vssd vssd vccd vccd _0567_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_29_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1328_ _1328_/A vssd vssd vccd vccd _1328_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1259_ _1515_/A _1259_/B _1259_/C vssd vssd vccd vccd _1260_/A sky130_fd_sc_hd__and3b_2
XFILLER_37_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input230_A la_iena_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input328_A la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0495__A _0495_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1103__B _1103_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0630_ _0630_/A vssd vssd vccd vccd _0630_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0561_ _0561_/A vssd vssd vccd vccd _0561_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_49_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0492_ _0492_/A vssd vssd vccd vccd _0492_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_2128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1113_ _1369_/A _1113_/B _1113_/C vssd vssd vccd vccd _1114_/A sky130_fd_sc_hd__and3b_4
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] _0726_/X vssd vssd vccd vccd _0504_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1044_ _1044_/A vssd vssd vccd vccd _1044_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1013__B _1013_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_726 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0828_ _0828_/A vssd vssd vccd vccd _0828_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_wb_dat_gates\[5\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0759_ _0759_/A _0759_/B vssd vssd vccd vccd _0760_/A sky130_fd_sc_hd__and2_4
XFILLER_46_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1204__A _1204_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_770 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1882 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input180_A la_iena_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input278_A la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input445_A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input41_A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3998 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0937__B _0937_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1114__A _1114_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_4036 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output664_A _0495_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1133__A_N _1389_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3926 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0613_ _0613_/A _0613_/B vssd vssd vccd vccd _0614_/A sky130_fd_sc_hd__and2_1
XANTENNA_output831_A _1448_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output929_A _1004_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0544_ _0544_/A vssd vssd vccd vccd _0544_/Y sky130_fd_sc_hd__inv_2
XTAP_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0475_ _0475_/A vssd vssd vccd vccd _0475_/Y sky130_fd_sc_hd__inv_2
XTAP_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0847__B _0847_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1024__A _1024_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1027_ _1283_/A _1027_/B _1027_/C vssd vssd vccd vccd _1028_/A sky130_fd_sc_hd__and3b_1
XANTENNA__0863__A _0863_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0757__B _0757_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_840 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0773__A _0773_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_9_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input395_A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input89_A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0667__B _0667_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput350 la_oenb_mprj[66] vssd vssd vccd vccd _1407_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput361 la_oenb_mprj[76] vssd vssd vccd vccd _1427_/A sky130_fd_sc_hd__buf_4
Xinput372 la_oenb_mprj[86] vssd vssd vccd vccd _1447_/A sky130_fd_sc_hd__clkbuf_8
Xinput383 la_oenb_mprj[96] vssd vssd vccd vccd _1467_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput394 mprj_adr_o_core[15] vssd vssd vccd vccd _0921_/B sky130_fd_sc_hd__buf_8
XFILLER_23_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0683__A _0683_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output879_A _0910_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1410 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput802 _1286_/X vssd vssd vccd vccd la_oenb_core[5] sky130_fd_sc_hd__buf_12
XFILLER_9_3723 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput813 _1288_/X vssd vssd vccd vccd la_oenb_core[6] sky130_fd_sc_hd__buf_12
Xoutput824 _1290_/X vssd vssd vccd vccd la_oenb_core[7] sky130_fd_sc_hd__buf_12
Xoutput835 _1292_/X vssd vssd vccd vccd la_oenb_core[8] sky130_fd_sc_hd__buf_12
XFILLER_6_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput846 _1294_/X vssd vssd vccd vccd la_oenb_core[9] sky130_fd_sc_hd__buf_12
XFILLER_29_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput857 _0928_/X vssd vssd vccd vccd mprj_adr_o_user[18] sky130_fd_sc_hd__buf_12
XFILLER_9_3778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput868 _0948_/X vssd vssd vccd vccd mprj_adr_o_user[28] sky130_fd_sc_hd__buf_12
XFILLER_3_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput879 _0910_/X vssd vssd vccd vccd mprj_adr_o_user[9] sky130_fd_sc_hd__buf_12
XFILLER_25_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0527_ _0527_/A vssd vssd vccd vccd _0527_/Y sky130_fd_sc_hd__inv_2
XTAP_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0858__A _0858_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1029__A_N _1285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1179__A_N _1435_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0593__A _0593_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__1201__B _1201_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3784 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0768__A _0768_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input143_A la_iena_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input310_A la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input408_A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1111__B _1111_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1430_ _1430_/A vssd vssd vccd vccd _1430_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3879 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1361_ _1361_/A _1361_/B vssd vssd vccd vccd _1362_/A sky130_fd_sc_hd__and2_1
XFILLER_29_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1292_ _1292_/A vssd vssd vccd vccd _1292_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput180 la_iena_mprj[28] vssd vssd vccd vccd _0663_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_23_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput191 la_iena_mprj[38] vssd vssd vccd vccd _0683_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_40_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_4042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] _0690_/X vssd vssd vccd vccd _0486_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_53_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1302__A _1302_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1021__B _1021_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput610 _0562_/Y vssd vssd vccd vccd la_data_in_mprj[117] sky130_fd_sc_hd__buf_12
Xoutput621 _0572_/Y vssd vssd vccd vccd la_data_in_mprj[127] sky130_fd_sc_hd__buf_12
Xoutput632 _0466_/Y vssd vssd vccd vccd la_data_in_mprj[21] sky130_fd_sc_hd__buf_12
XFILLER_47_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput643 _0476_/Y vssd vssd vccd vccd la_data_in_mprj[31] sky130_fd_sc_hd__buf_12
XFILLER_9_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput654 _0486_/Y vssd vssd vccd vccd la_data_in_mprj[41] sky130_fd_sc_hd__buf_12
XFILLER_5_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput665 _0496_/Y vssd vssd vccd vccd la_data_in_mprj[51] sky130_fd_sc_hd__buf_12
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] _0614_/X vssd vssd vccd vccd _1536_/A
+ sky130_fd_sc_hd__nand2_2
Xoutput676 _0506_/Y vssd vssd vccd vccd la_data_in_mprj[61] sky130_fd_sc_hd__buf_12
XFILLER_25_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput687 _0516_/Y vssd vssd vccd vccd la_data_in_mprj[71] sky130_fd_sc_hd__buf_12
Xoutput698 _0526_/Y vssd vssd vccd vccd la_data_in_mprj[81] sky130_fd_sc_hd__buf_12
XFILLER_42_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1212__A _1212_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input260_A la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input358_A la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0945__B _0945_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1122__A _1122_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0930_ _0930_/A vssd vssd vccd vccd _0930_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0861_ _0861_/A _0861_/B vssd vssd vccd vccd _0862_/A sky130_fd_sc_hd__and2_2
XFILLER_31_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0792_ _0792_/A vssd vssd vccd vccd _0792_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output744_A _1520_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] _0786_/X vssd vssd vccd vccd _0534_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA_output911_A _0584_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1413_ _1413_/A _1413_/B vssd vssd vccd vccd _1414_/A sky130_fd_sc_hd__and2_1
XFILLER_26_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1386 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1344_ _1344_/A vssd vssd vccd vccd _1344_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1275_ _1275_/A _1275_/B vssd vssd vccd vccd _1276_/A sky130_fd_sc_hd__and2_1
XFILLER_4_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0855__B _0855_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1217__A_N _1473_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput473 _1238_/X vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__buf_12
XFILLER_5_3225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput484 _1258_/X vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__buf_12
XFILLER_43_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput495 _1046_/X vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__buf_12
XFILLER_5_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0765__B _0765_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0781__A _0781_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_658 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input71_A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1060_ _1060_/A vssd vssd vccd vccd _1060_/X sky130_fd_sc_hd__buf_2
XFILLER_4_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0675__B _0675_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0691__A _0691_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output861_A _0934_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0913_ _0913_/A _0913_/B vssd vssd vccd vccd _0914_/A sky130_fd_sc_hd__and2_2
XFILLER_32_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[17\] mprj_dat_i_user[17] _0870_/X vssd vssd vccd vccd _0593_/A
+ sky130_fd_sc_hd__nand2_2
X_0844_ _0844_/A vssd vssd vccd vccd _0844_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3006 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0775_ _0775_/A _0775_/B vssd vssd vccd vccd _0776_/A sky130_fd_sc_hd__and2_4
XFILLER_28_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1327_ _1327_/A _1327_/B vssd vssd vccd vccd _1328_/A sky130_fd_sc_hd__and2_1
XFILLER_39_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] _0838_/X vssd vssd vccd vccd _0560_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1258_ _1258_/A vssd vssd vccd vccd _1258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1189_ _1445_/A _1189_/B _1189_/C vssd vssd vccd vccd _1190_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_2498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0776__A _0776_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input223_A la_iena_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1103__C _1103_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1400__A _1400_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2887 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0560_ _0560_/A vssd vssd vccd vccd _0560_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0491_ _0491_/A vssd vssd vccd vccd _0491_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output707_A _1541_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1112_ _1112_/A vssd vssd vccd vccd _1112_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1043_ _1299_/A _1043_/B _1043_/C vssd vssd vccd vccd _1044_/A sky130_fd_sc_hd__and3b_1
XFILLER_17_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1310__A _1310_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0827_ _0827_/A _0827_/B vssd vssd vccd vccd _0828_/A sky130_fd_sc_hd__and2_2
XFILLER_11_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0758_ _0758_/A vssd vssd vccd vccd _0758_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_0689_ _0689_/A _0689_/B vssd vssd vccd vccd _0690_/A sky130_fd_sc_hd__and2_1
XFILLER_44_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0596__A _0596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3826 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1220__A _1220_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input173_A la_iena_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input340_A la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1085__A_N _1341_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input438_A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input34_A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0953__B _0953_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_576 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[59\]_B _0726_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1130__A _1130_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output657_A _0489_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0612_ _0612_/A vssd vssd vccd vccd _0612_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_3938 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0543_ _0543_/A vssd vssd vccd vccd _0543_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0474_ _0474_/A vssd vssd vccd vccd _0474_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] _0750_/X vssd vssd vccd vccd _0516_/A
+ sky130_fd_sc_hd__nand2_2
XTAP_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1305__A _1305_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1026_ _1026_/A vssd vssd vccd vccd _1026_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0863__B _0863_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1040__A _1040_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_852 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input290_A la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input388_A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1109__B _1109_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput340 la_oenb_mprj[57] vssd vssd vccd vccd _1389_/A sky130_fd_sc_hd__buf_4
XFILLER_48_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput351 la_oenb_mprj[67] vssd vssd vccd vccd _1409_/A sky130_fd_sc_hd__buf_2
Xinput362 la_oenb_mprj[77] vssd vssd vccd vccd _1429_/A sky130_fd_sc_hd__buf_4
XFILLER_49_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput373 la_oenb_mprj[87] vssd vssd vccd vccd _1449_/A sky130_fd_sc_hd__buf_6
Xinput384 la_oenb_mprj[97] vssd vssd vccd vccd _1469_/A sky130_fd_sc_hd__clkbuf_4
Xinput395 mprj_adr_o_core[16] vssd vssd vccd vccd _0923_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_40_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0683__B _0683_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output941_A _0968_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3702 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput803 _1396_/X vssd vssd vccd vccd la_oenb_core[60] sky130_fd_sc_hd__buf_12
Xoutput814 _1416_/X vssd vssd vccd vccd la_oenb_core[70] sky130_fd_sc_hd__buf_12
XFILLER_9_3735 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput825 _1436_/X vssd vssd vccd vccd la_oenb_core[80] sky130_fd_sc_hd__buf_12
XFILLER_47_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput836 _1456_/X vssd vssd vccd vccd la_oenb_core[90] sky130_fd_sc_hd__buf_12
XANTENNA__1019__B _1019_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput847 _0608_/Y vssd vssd vccd vccd mprj_ack_i_core sky130_fd_sc_hd__buf_12
Xoutput858 _0930_/X vssd vssd vccd vccd mprj_adr_o_user[19] sky130_fd_sc_hd__buf_12
Xoutput869 _0950_/X vssd vssd vccd vccd mprj_adr_o_user[29] sky130_fd_sc_hd__buf_12
XFILLER_47_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0526_ _0526_/A vssd vssd vccd vccd _0526_/Y sky130_fd_sc_hd__inv_2
XTAP_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[25\]_A mprj_dat_i_user[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0874__A _0874_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1009_ _1009_/A _1009_/B vssd vssd vccd vccd _1010_/A sky130_fd_sc_hd__and2_4
XFILLER_22_343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[16\]_A mprj_dat_i_user[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input136_A la_iena_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0784__A _0784_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1123__A_N _1379_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input303_A la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1273__A_N _1529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0959__A _0959_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1360_ _1360_/A vssd vssd vccd vccd _1360_/X sky130_fd_sc_hd__buf_2
XFILLER_4_3621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output522_A _1096_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1291_ _1291_/A _1291_/B vssd vssd vccd vccd _1292_/A sky130_fd_sc_hd__and2_4
XFILLER_49_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput170 la_iena_mprj[19] vssd vssd vccd vccd _0645_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput181 la_iena_mprj[29] vssd vssd vccd vccd _0665_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_4_2986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput192 la_iena_mprj[39] vssd vssd vccd vccd _0685_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] _0676_/X vssd vssd vccd vccd _0479_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_18_3364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_170 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1021__C _1021_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput600 _0553_/Y vssd vssd vccd vccd la_data_in_mprj[108] sky130_fd_sc_hd__buf_12
Xoutput611 _0563_/Y vssd vssd vccd vccd la_data_in_mprj[118] sky130_fd_sc_hd__buf_12
Xoutput622 _1545_/Y vssd vssd vccd vccd la_data_in_mprj[12] sky130_fd_sc_hd__buf_12
XFILLER_29_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput633 _0467_/Y vssd vssd vccd vccd la_data_in_mprj[22] sky130_fd_sc_hd__buf_12
XFILLER_44_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0869__A _0869_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput644 _0477_/Y vssd vssd vccd vccd la_data_in_mprj[32] sky130_fd_sc_hd__buf_12
XFILLER_28_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput655 _0487_/Y vssd vssd vccd vccd la_data_in_mprj[42] sky130_fd_sc_hd__buf_12
XFILLER_9_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput666 _0497_/Y vssd vssd vccd vccd la_data_in_mprj[52] sky130_fd_sc_hd__buf_12
Xoutput677 _0507_/Y vssd vssd vccd vccd la_data_in_mprj[62] sky130_fd_sc_hd__buf_12
XFILLER_29_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput688 _0517_/Y vssd vssd vccd vccd la_data_in_mprj[72] sky130_fd_sc_hd__buf_12
XFILLER_25_3379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput699 _0527_/Y vssd vssd vccd vccd la_data_in_mprj[82] sky130_fd_sc_hd__buf_12
X_0509_ _0509_/A vssd vssd vccd vccd _0509_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1489_ _1489_/A _1489_/B vssd vssd vccd vccd _1490_/A sky130_fd_sc_hd__and2_1
XFILLER_41_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0779__A _0779_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input253_A la_iena_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input420_A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1403__A _1403_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0961__B _0961_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1019__A_N _1275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0860_ _0860_/A vssd vssd vccd vccd _0860_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output472_A _1236_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0791_ _0791_/A _0791_/B vssd vssd vccd vccd _0792_/A sky130_fd_sc_hd__and2_4
XFILLER_31_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0689__A _0689_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1169__A_N _1425_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output737_A _1508_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1412_ _1412_/A vssd vssd vccd vccd _1412_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1343_ _1343_/A _1343_/B vssd vssd vccd vccd _1344_/A sky130_fd_sc_hd__and2_2
XFILLER_29_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1274_ _1274_/A vssd vssd vccd vccd _1274_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1313__A _1313_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0871__B _0871_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0989_ _0989_/A _0989_/B vssd vssd vccd vccd _0990_/A sky130_fd_sc_hd__and2_4
XFILLER_27_2707 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput463 _1020_/X vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__buf_12
Xoutput474 _1040_/X vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__buf_12
Xoutput485 _1042_/X vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__buf_12
XFILLER_5_3237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput496 _1048_/X vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__buf_12
XANTENNA__1207__B _1207_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0781__B _0781_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_622 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input370_A la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input64_A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1117__B _1117_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0972__A _0972_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0691__B _0691_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0912_ _0912_/A vssd vssd vccd vccd _0912_/X sky130_fd_sc_hd__buf_6
XFILLER_32_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output854_A _0922_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0843_ _0843_/A _0843_/B vssd vssd vccd vccd _0844_/A sky130_fd_sc_hd__and2_1
XFILLER_31_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0774_ _0774_/A vssd vssd vccd vccd _0774_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1308__A _1308_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1616 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1027__B _1027_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1326_ _1326_/A vssd vssd vccd vccd _1326_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1257_ _1513_/A _1257_/B _1257_/C vssd vssd vccd vccd _1258_/A sky130_fd_sc_hd__and3b_2
XFILLER_37_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] _0824_/X vssd vssd vccd vccd _0553_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_39_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1188_ _1188_/A vssd vssd vccd vccd _1188_/X sky130_fd_sc_hd__buf_2
XFILLER_37_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0882__A _0882_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[8\]_A mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_618 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1218__A _1218_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input216_A la_iena_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0792__A _0792_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1128__A _1128_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0490_ _0490_/A vssd vssd vccd vccd _0490_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_3783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3658 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0967__A _0967_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1207__A_N _1463_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1111_ _1367_/A _1111_/B _1111_/C vssd vssd vccd vccd _1112_/A sky130_fd_sc_hd__and3b_2
XFILLER_1_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output602_A _1543_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1042_ _1042_/A vssd vssd vccd vccd _1042_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0826_ _0826_/A vssd vssd vccd vccd _0826_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0757_ _0757_/A _0757_/B vssd vssd vccd vccd _0758_/A sky130_fd_sc_hd__and2_2
XFILLER_28_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1038__A _1038_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0688_ _0688_/A vssd vssd vccd vccd _0688_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1309_ _1309_/A _1309_/B vssd vssd vccd vccd _1310_/A sky130_fd_sc_hd__and2_4
XFILLER_29_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1501__A _1501_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3838 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3912 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input166_A la_iena_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0787__A _0787_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input333_A la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input27_A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1411__A _1411_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1751 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0611_ _0611_/A _0611_/B vssd vssd vccd vccd _0612_/A sky130_fd_sc_hd__and2_1
XANTENNA_output552_A _1150_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0542_ _0542_/A vssd vssd vccd vccd _0542_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0697__A _0697_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output817_A _1422_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0473_ _0473_/A vssd vssd vccd vccd _0473_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1305__B _1305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] _0736_/X vssd vssd vccd vccd _0509_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_22_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1025_ _1281_/A _1025_/B _1025_/C vssd vssd vccd vccd _1026_/A sky130_fd_sc_hd__and3b_1
XFILLER_35_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1321__A _1321_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0809_ _0809_/A _0809_/B vssd vssd vccd vccd _0810_/A sky130_fd_sc_hd__and2_4
XFILLER_28_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1215__B _1215_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input283_A la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input450_A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1109__C _1109_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1406__A _1406_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput330 la_oenb_mprj[48] vssd vssd vccd vccd _1371_/A sky130_fd_sc_hd__buf_6
XFILLER_4_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput341 la_oenb_mprj[58] vssd vssd vccd vccd _1391_/A sky130_fd_sc_hd__buf_2
XANTENNA__1125__B _1125_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput352 la_oenb_mprj[68] vssd vssd vccd vccd _1411_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput363 la_oenb_mprj[78] vssd vssd vccd vccd _1431_/A sky130_fd_sc_hd__buf_4
Xinput374 la_oenb_mprj[88] vssd vssd vccd vccd _1451_/A sky130_fd_sc_hd__buf_4
XFILLER_29_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput385 la_oenb_mprj[98] vssd vssd vccd vccd _1471_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput396 mprj_adr_o_core[17] vssd vssd vccd vccd _0925_/B sky130_fd_sc_hd__buf_6
XFILLER_35_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0980__A _0980_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput804 _1398_/X vssd vssd vccd vccd la_oenb_core[61] sky130_fd_sc_hd__buf_12
XANTENNA_output934_A _1014_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput815 _1418_/X vssd vssd vccd vccd la_oenb_core[71] sky130_fd_sc_hd__buf_12
Xoutput826 _1438_/X vssd vssd vccd vccd la_oenb_core[81] sky130_fd_sc_hd__buf_12
XFILLER_9_3747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput837 _1458_/X vssd vssd vccd vccd la_oenb_core[91] sky130_fd_sc_hd__buf_12
XFILLER_6_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1019__C input4/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput848 _0892_/X vssd vssd vccd vccd mprj_adr_o_user[0] sky130_fd_sc_hd__buf_12
XFILLER_28_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput859 _0894_/X vssd vssd vccd vccd mprj_adr_o_user[1] sky130_fd_sc_hd__buf_12
XFILLER_25_2805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0525_ _0525_/A vssd vssd vccd vccd _0525_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1316__A _1316_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1035__B _1035_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[25\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1008_ _1008_/A vssd vssd vccd vccd _1008_/X sky130_fd_sc_hd__buf_6
XFILLER_52_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0890__A _0890_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1075__A_N _1331_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1226__A _1226_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[16\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input129_A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input94_A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0959__B _0959_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1136__A _1136_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1290_ _1290_/A vssd vssd vccd vccd _1290_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0975__A _0975_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output515_A _1082_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_irq_gates\[1\]_A user_irq_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput160 la_iena_mprj[125] vssd vssd vccd vccd _0857_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput171 la_iena_mprj[1] vssd vssd vccd vccd _0609_/B sky130_fd_sc_hd__clkbuf_1
Xinput182 la_iena_mprj[2] vssd vssd vccd vccd _0611_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_18_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput193 la_iena_mprj[3] vssd vssd vccd vccd _0613_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4066 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output884_A _0588_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_182 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] _0662_/X vssd vssd vccd vccd _0472_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_31_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput601 _0554_/Y vssd vssd vccd vccd la_data_in_mprj[109] sky130_fd_sc_hd__buf_12
XFILLER_25_4037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput612 _0564_/Y vssd vssd vccd vccd la_data_in_mprj[119] sky130_fd_sc_hd__buf_12
XFILLER_25_3303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput623 _1546_/Y vssd vssd vccd vccd la_data_in_mprj[13] sky130_fd_sc_hd__buf_12
Xoutput634 _0468_/Y vssd vssd vccd vccd la_data_in_mprj[23] sky130_fd_sc_hd__buf_12
Xoutput645 _0478_/Y vssd vssd vccd vccd la_data_in_mprj[33] sky130_fd_sc_hd__buf_12
XFILLER_47_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput656 _0488_/Y vssd vssd vccd vccd la_data_in_mprj[43] sky130_fd_sc_hd__buf_12
XFILLER_25_3347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput667 _0498_/Y vssd vssd vccd vccd la_data_in_mprj[53] sky130_fd_sc_hd__buf_12
Xoutput678 _0508_/Y vssd vssd vccd vccd la_data_in_mprj[63] sky130_fd_sc_hd__buf_12
Xoutput689 _0518_/Y vssd vssd vccd vccd la_data_in_mprj[73] sky130_fd_sc_hd__buf_12
XFILLER_29_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1046__A _1046_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0508_ _0508_/A vssd vssd vccd vccd _0508_/Y sky130_fd_sc_hd__inv_2
X_1488_ _1488_/A vssd vssd vccd vccd _1488_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0885__A _0885_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input246_A la_iena_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0795__A _0795_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input413_A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1403__B _1403_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0790_ _0790_/A vssd vssd vccd vccd _0790_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output465_A _1222_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0689__B _0689_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1411_ _1411_/A _1411_/B vssd vssd vccd vccd _1412_/A sky130_fd_sc_hd__and2_1
XANTENNA_output632_A _0466_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1342_ _1342_/A vssd vssd vccd vccd _1342_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_3430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1273_ _1529_/A _1273_/B _1273_/C vssd vssd vccd vccd _1274_/A sky130_fd_sc_hd__and3b_1
XFILLER_20_3244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1313__B _1313_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0988_ _0988_/A vssd vssd vccd vccd _0988_/X sky130_fd_sc_hd__buf_6
XANTENNA__1113__A_N _1369_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2719 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput464 _1220_/X vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__buf_12
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput475 _1240_/X vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__buf_12
XFILLER_47_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput486 _1260_/X vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__buf_12
Xoutput497 _1050_/X vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__buf_12
XFILLER_5_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1263__A_N _1519_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input1_A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1223__B _1223_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input196_A la_iena_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input363_A la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input57_A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1117__C _1117_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1414__A _1414_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1133__B _1133_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0911_ _0911_/A _0911_/B vssd vssd vccd vccd _0912_/A sky130_fd_sc_hd__and2_1
XANTENNA_output582_A _1204_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0842_ _0842_/A vssd vssd vccd vccd _0842_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0773_ _0773_/A _0773_/B vssd vssd vccd vccd _0774_/A sky130_fd_sc_hd__and2_4
XANTENNA_output847_A _0608_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] _0796_/X vssd vssd vccd vccd _0539_/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1628 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1325_ _1325_/A _1325_/B vssd vssd vccd vccd _1326_/A sky130_fd_sc_hd__and2_4
XFILLER_22_2627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1324__A _1324_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1256_ _1256_/A vssd vssd vccd vccd _1256_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1043__B _1043_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1187_ _1443_/A _1187_/B _1187_/C vssd vssd vccd vccd _1188_/A sky130_fd_sc_hd__and3b_1
XFILLER_25_715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[8\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3840 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1234__A _1234_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input111_A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input209_A la_iena_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__1159__A_N _1415_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1409__A _1409_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0967__B _0967_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1144__A _1144_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1110_ _1110_/A vssd vssd vccd vccd _1110_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_3455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1041_ _1297_/A _1041_/B _1041_/C vssd vssd vccd vccd _1042_/A sky130_fd_sc_hd__and3b_4
XFILLER_24_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0983__A _0983_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[22\] mprj_dat_i_user[22] _0870_/X vssd vssd vccd vccd _0598_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_15_2464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0825_ _0825_/A _0825_/B vssd vssd vccd vccd _0826_/A sky130_fd_sc_hd__and2_1
XANTENNA__1319__A _1319_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0756_ _0756_/A vssd vssd vccd vccd _0756_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0687_ _0687_/A _0687_/B vssd vssd vccd vccd _0688_/A sky130_fd_sc_hd__and2_1
XFILLER_6_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0877__B _0877_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] _0848_/X vssd vssd vccd vccd _0565_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__1054__A _1054_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_1308_ _1308_/A vssd vssd vccd vccd _1308_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_2479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1239_ _1495_/A _1239_/B _1239_/C vssd vssd vccd vccd _1240_/A sky130_fd_sc_hd__and3b_2
XANTENNA__0893__A _0893_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1501__B _1501_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input159_A la_iena_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input326_A la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1411__B _1411_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_887 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0610_ _0610_/A vssd vssd vccd vccd _0610_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0541_ _0541_/A vssd vssd vccd vccd _0541_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1671 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0978__A _0978_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0472_ _0472_/A vssd vssd vccd vccd _0472_/Y sky130_fd_sc_hd__clkinv_2
XTAP_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0697__B _0697_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] _0722_/X vssd vssd vccd vccd _0502_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_1_2540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1024_ _1024_/A vssd vssd vccd vccd _1024_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_35_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1321__B _1321_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0808_ _0808_/A vssd vssd vccd vccd _0808_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0888__A _0888_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0739_ _0739_/A _0739_/B vssd vssd vccd vccd _0740_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1215__C _1215_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1231__B _1231_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input276_A la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0798__A _0798_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input443_A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput320 la_oenb_mprj[39] vssd vssd vccd vccd _1353_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_48_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput331 la_oenb_mprj[49] vssd vssd vccd vccd _1373_/A sky130_fd_sc_hd__buf_2
Xinput342 la_oenb_mprj[59] vssd vssd vccd vccd _1393_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_7_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput353 la_oenb_mprj[69] vssd vssd vccd vccd _1413_/A sky130_fd_sc_hd__buf_2
XANTENNA__1125__C _1125_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput364 la_oenb_mprj[79] vssd vssd vccd vccd _1433_/A sky130_fd_sc_hd__buf_4
Xinput375 la_oenb_mprj[89] vssd vssd vccd vccd _1453_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput386 la_oenb_mprj[99] vssd vssd vccd vccd _1473_/A sky130_fd_sc_hd__clkbuf_4
Xinput397 mprj_adr_o_core[18] vssd vssd vccd vccd _0927_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_2_3594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1422__A _1422_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1141__B _1141_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output495_A _1046_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput805 _1400_/X vssd vssd vccd vccd la_oenb_core[62] sky130_fd_sc_hd__buf_12
XFILLER_47_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput816 _1420_/X vssd vssd vccd vccd la_oenb_core[72] sky130_fd_sc_hd__buf_12
Xoutput827 _1440_/X vssd vssd vccd vccd la_oenb_core[82] sky130_fd_sc_hd__buf_12
Xoutput838 _1460_/X vssd vssd vccd vccd la_oenb_core[92] sky130_fd_sc_hd__buf_12
Xoutput849 _0912_/X vssd vssd vccd vccd mprj_adr_o_user[10] sky130_fd_sc_hd__buf_12
XANTENNA_output927_A _1000_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0501__A _0501_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0524_ _0524_/A vssd vssd vccd vccd _0524_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1035__C _1035_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1332__A _1332_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1051__B _1051_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1007_ _1007_/A _1007_/B vssd vssd vccd vccd _1008_/A sky130_fd_sc_hd__and2_4
XFILLER_35_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1800 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1507__A _1507_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1242__A _1242_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input393_A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input87_A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1417__A _1417_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput150 la_iena_mprj[116] vssd vssd vccd vccd _0839_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_2883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0975__B _0975_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput161 la_iena_mprj[126] vssd vssd vccd vccd _0859_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput172 la_iena_mprj[20] vssd vssd vccd vccd _0647_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_48_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput183 la_iena_mprj[30] vssd vssd vccd vccd _0667_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_output508_A _1070_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput194 la_iena_mprj[40] vssd vssd vccd vccd _0687_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_18_4023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1152__A _1152_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0991__A _0991_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output877_A _0906_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput602 _1543_/Y vssd vssd vccd vccd la_data_in_mprj[10] sky130_fd_sc_hd__buf_12
Xoutput613 _1544_/Y vssd vssd vccd vccd la_data_in_mprj[11] sky130_fd_sc_hd__buf_12
Xoutput624 _1547_/Y vssd vssd vccd vccd la_data_in_mprj[14] sky130_fd_sc_hd__buf_12
XFILLER_29_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput635 _0469_/Y vssd vssd vccd vccd la_data_in_mprj[24] sky130_fd_sc_hd__buf_12
XANTENNA__1327__A _1327_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput646 _0479_/Y vssd vssd vccd vccd la_data_in_mprj[34] sky130_fd_sc_hd__buf_12
Xoutput657 _0489_/Y vssd vssd vccd vccd la_data_in_mprj[44] sky130_fd_sc_hd__buf_12
XFILLER_28_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput668 _0499_/Y vssd vssd vccd vccd la_data_in_mprj[54] sky130_fd_sc_hd__buf_12
Xoutput679 _0509_/Y vssd vssd vccd vccd la_data_in_mprj[64] sky130_fd_sc_hd__buf_12
XFILLER_25_3359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0507_ _0507_/A vssd vssd vccd vccd _0507_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1487_ _1487_/A _1487_/B vssd vssd vccd vccd _1488_/A sky130_fd_sc_hd__and2_1
XFILLER_23_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1062__A _1062_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input141_A la_iena_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input239_A la_iena_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input406_A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1410_ _1410_/A vssd vssd vccd vccd _1410_/X sky130_fd_sc_hd__buf_2
XFILLER_29_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1341_ _1341_/A _1341_/B vssd vssd vccd vccd _1342_/A sky130_fd_sc_hd__and2_2
XFILLER_25_1209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0986__A _0986_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output625_A _1548_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1065__A_N _1321_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1272_ _1272_/A vssd vssd vccd vccd _1272_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0987_ _0987_/A _0987_/B vssd vssd vccd vccd _0988_/A sky130_fd_sc_hd__and2_2
XFILLER_9_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] _0610_/X vssd vssd vccd vccd _1534_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput465 _1222_/X vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__buf_12
Xoutput476 _1242_/X vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__buf_12
XFILLER_44_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput487 _1262_/X vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__buf_12
Xoutput498 _1052_/X vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__buf_12
XANTENNA__0896__A _0896_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1539_ _1539_/A vssd vssd vccd vccd _1539_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_418 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1520__A _1520_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input189_A la_iena_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input356_A la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1133__C _1133_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_790 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1430__A _1430_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0910_ _0910_/A vssd vssd vccd vccd _0910_/X sky130_fd_sc_hd__buf_6
XFILLER_53_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0841_ _0841_/A _0841_/B vssd vssd vccd vccd _0842_/A sky130_fd_sc_hd__and2_1
XANTENNA_output575_A _1192_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0772_ _0772_/A vssd vssd vccd vccd _0772_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3908 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] _0782_/X vssd vssd vccd vccd _0532_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_2814 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1324_ _1324_/A vssd vssd vccd vccd _1324_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1255_ _1511_/A _1255_/B _1255_/C vssd vssd vccd vccd _1256_/A sky130_fd_sc_hd__and3b_2
XFILLER_0_3169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1043__C _1043_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1186_ _1186_/A vssd vssd vccd vccd _1186_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_25_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1340__A _1340_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1515__A _1515_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3852 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1250__A _1250_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input104_A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1409__B _1409_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1425__A _1425_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1662 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1040_ _1040_/A vssd vssd vccd vccd _1040_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0983__B _0983_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1103__A_N _1359_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1253__A_N _1509_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[15\] mprj_dat_i_user[15] _0870_/X vssd vssd vccd vccd _0591_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA__0504__A _0504_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0824_ _0824_/A vssd vssd vccd vccd _0824_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1319__B _1319_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0755_ _0755_/A _0755_/B vssd vssd vccd vccd _0756_/A sky130_fd_sc_hd__and2_1
XFILLER_6_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0686_ _0686_/A vssd vssd vccd vccd _0686_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1335__A _1335_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1307_ _1307_/A _1307_/B vssd vssd vccd vccd _1308_/A sky130_fd_sc_hd__and2_2
XFILLER_29_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] _0834_/X vssd vssd vccd vccd _0558_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_6_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__0893__B _0893_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1238_ _1238_/A vssd vssd vccd vccd _1238_/X sky130_fd_sc_hd__buf_2
XFILLER_39_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1169_ _1425_/A _1169_/B _1169_/C vssd vssd vccd vccd _1170_/A sky130_fd_sc_hd__and3b_1
XFILLER_25_535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1070__A _1070_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1229__B _1229_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input221_A la_iena_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input319_A la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_62 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1628 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1139__B _1139_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0540_ _0540_/A vssd vssd vccd vccd _0540_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0471_ _0471_/A vssd vssd vccd vccd _0471_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output538_A _1124_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0994__A _0994_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1023_ _1279_/A _1023_/B _1023_/C vssd vssd vccd vccd _1024_/A sky130_fd_sc_hd__and3b_1
XFILLER_35_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1049__B _1049_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0807_ _0807_/A _0807_/B vssd vssd vccd vccd _0808_/A sky130_fd_sc_hd__and2_4
XFILLER_11_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_0738_ _0738_/A vssd vssd vccd vccd _0738_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1149__A_N _1405_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_0669_ _0669_/A _0669_/B vssd vssd vccd vccd _0670_/A sky130_fd_sc_hd__and2_1
XFILLER_28_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[28\]_A mprj_dat_i_user[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1231__C _1231_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input171_A la_iena_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input269_A la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[19\]_A mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input436_A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput310 la_oenb_mprj[2] vssd vssd vccd vccd _1279_/A sky130_fd_sc_hd__buf_2
XFILLER_40_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput321 la_oenb_mprj[3] vssd vssd vccd vccd _1281_/A sky130_fd_sc_hd__buf_2
XFILLER_24_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input32_A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput332 la_oenb_mprj[4] vssd vssd vccd vccd _1283_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput343 la_oenb_mprj[5] vssd vssd vccd vccd _1285_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_3078 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput354 la_oenb_mprj[6] vssd vssd vccd vccd _1287_/A sky130_fd_sc_hd__clkbuf_2
Xinput365 la_oenb_mprj[7] vssd vssd vccd vccd _1289_/A sky130_fd_sc_hd__clkbuf_2
Xinput376 la_oenb_mprj[8] vssd vssd vccd vccd _1291_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput387 la_oenb_mprj[9] vssd vssd vccd vccd _1293_/A sky130_fd_sc_hd__clkbuf_2
Xinput398 mprj_adr_o_core[19] vssd vssd vccd vccd _0929_/B sky130_fd_sc_hd__buf_8
XFILLER_29_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1141__C _1141_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output488_A _1264_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0989__A _0989_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output655_A _0487_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput806 _1402_/X vssd vssd vccd vccd la_oenb_core[63] sky130_fd_sc_hd__buf_12
Xoutput817 _1422_/X vssd vssd vccd vccd la_oenb_core[73] sky130_fd_sc_hd__buf_12
XFILLER_6_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput828 _1442_/X vssd vssd vccd vccd la_oenb_core[83] sky130_fd_sc_hd__buf_12
XFILLER_29_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput839 _1462_/X vssd vssd vccd vccd la_oenb_core[93] sky130_fd_sc_hd__buf_12
XFILLER_45_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0523_ _0523_/A vssd vssd vccd vccd _0523_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1051__C _1051_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_1006_ _1006_/A vssd vssd vccd vccd _1006_/X sky130_fd_sc_hd__buf_6
XFILLER_1_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0899__A _0899_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1507__B _1507_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1523__A _1523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1996 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3868 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input386_A la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1417__B _1417_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput140 la_iena_mprj[107] vssd vssd vccd vccd _0821_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput151 la_iena_mprj[117] vssd vssd vccd vccd _0841_/B sky130_fd_sc_hd__buf_2
XANTENNA__1433__A _1433_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput162 la_iena_mprj[127] vssd vssd vccd vccd _0861_/B sky130_fd_sc_hd__clkbuf_1
Xinput173 la_iena_mprj[21] vssd vssd vccd vccd _0649_/B sky130_fd_sc_hd__clkbuf_1
Xinput184 la_iena_mprj[31] vssd vssd vccd vccd _0669_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_48_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput195 la_iena_mprj[41] vssd vssd vccd vccd _0689_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_490 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0991__B _0991_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput603 _0555_/Y vssd vssd vccd vccd la_data_in_mprj[110] sky130_fd_sc_hd__buf_12
XANTENNA__0512__A _0512_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput614 _0565_/Y vssd vssd vccd vccd la_data_in_mprj[120] sky130_fd_sc_hd__buf_12
XFILLER_25_4039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput625 _1548_/Y vssd vssd vccd vccd la_data_in_mprj[15] sky130_fd_sc_hd__buf_12
XFILLER_47_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput636 _0470_/Y vssd vssd vccd vccd la_data_in_mprj[25] sky130_fd_sc_hd__buf_12
XFILLER_29_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput647 _0480_/Y vssd vssd vccd vccd la_data_in_mprj[35] sky130_fd_sc_hd__buf_12
Xoutput658 _0490_/Y vssd vssd vccd vccd la_data_in_mprj[45] sky130_fd_sc_hd__buf_12
XFILLER_47_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput669 _0500_/Y vssd vssd vccd vccd la_data_in_mprj[55] sky130_fd_sc_hd__buf_12
XFILLER_28_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0506_ _0506_/A vssd vssd vccd vccd _0506_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1486_ _1486_/A vssd vssd vccd vccd _1486_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1518__A _1518_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1237__B _1237_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input134_A la_iena_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input301_A la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1428__A _1428_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1340_ _1340_/A vssd vssd vccd vccd _1340_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output520_A _1092_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1271_ _1527_/A _1271_/B _1271_/C vssd vssd vccd vccd _1272_/A sky130_fd_sc_hd__and3b_1
XFILLER_24_3393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output618_A _0569_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] _0672_/X vssd vssd vccd vccd _0477_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__0507__A _0507_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0986_ _0986_/A vssd vssd vccd vccd _0986_/X sky130_fd_sc_hd__buf_6
XFILLER_9_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1338__A _1338_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1057__B _1057_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput466 _1224_/X vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__buf_12
XFILLER_25_2401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput477 _1244_/X vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__buf_12
XFILLER_47_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput488 _1264_/X vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__buf_12
X_1538_ _1538_/A vssd vssd vccd vccd _1538_/Y sky130_fd_sc_hd__inv_2
Xoutput499 _1054_/X vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__buf_12
XFILLER_42_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_1469_ _1469_/A _1469_/B vssd vssd vccd vccd _1470_/A sky130_fd_sc_hd__and2_1
XFILLER_41_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1248__A _1248_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input251_A la_iena_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input349_A la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0840_ _0840_/A vssd vssd vccd vccd _0840_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output470_A _1232_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0771_ _0771_/A _0771_/B vssd vssd vccd vccd _0772_/A sky130_fd_sc_hd__and2_4
XFILLER_10_3971 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output568_A _1034_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_662 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output735_A _1504_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0997__A _0997_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1323_ _1323_/A _1323_/B vssd vssd vccd vccd _1324_/A sky130_fd_sc_hd__and2_2
XFILLER_22_2618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1254_ _1254_/A vssd vssd vccd vccd _1254_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1185_ _1441_/A _1185_/B _1185_/C vssd vssd vccd vccd _1186_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0969_ _0969_/A _0969_/B vssd vssd vccd vccd _0970_/A sky130_fd_sc_hd__and2_2
XANTENNA__1068__A _1068_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1515__B _1515_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1531__A _1531_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1055__A_N _1311_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input299_A la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_426 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input62_A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1425__B _1425_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__1441__A _1441_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_0823_ _0823_/A _0823_/B vssd vssd vccd vccd _0824_/A sky130_fd_sc_hd__and2_2
XFILLER_31_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output852_A _0918_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0754_ _0754_/A vssd vssd vccd vccd _0754_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0685_ _0685_/A _0685_/B vssd vssd vccd vccd _0686_/A sky130_fd_sc_hd__and2_1
XFILLER_6_3313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__0520__A _0520_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__1335__B _1335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_1306_ _1306_/A vssd vssd vccd vccd _1306_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1237_ _1493_/A _1237_/B _1237_/C vssd vssd vccd vccd _1238_/A sky130_fd_sc_hd__and3b_4
XANTENNA__1351__A _1351_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] _0820_/X vssd vssd vccd vccd _0551_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_1168_ _1168_/A vssd vssd vccd vccd _1168_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1099_ _1355_/A _1099_/B _1099_/C vssd vssd vccd vccd _1100_/A sky130_fd_sc_hd__and3b_1
XFILLER_13_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1526__A _1526_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1245__B _1245_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input214_A la_iena_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1139__C _1139_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__1436__A _1436_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_0470_ _0470_/A vssd vssd vccd vccd _0470_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1155__B _1155_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output600_A _0553_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_1022_ _1022_/A vssd vssd vccd vccd _1022_/X sky130_fd_sc_hd__buf_4
XFILLER_1_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__0515__A _0515_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1049__C _1049_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0806_ _0806_/A vssd vssd vccd vccd _0806_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_0737_ _0737_/A _0737_/B vssd vssd vccd vccd _0738_/A sky130_fd_sc_hd__and2_1
XANTENNA__1346__A _1346_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_0668_ _0668_/A vssd vssd vccd vccd _0668_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__1065__B _1065_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[28\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_0599_ _0599_/A vssd vssd vccd vccd _0599_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1256__A _1256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input164_A la_iena_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[19\]_B _0870_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput300 la_oenb_mprj[20] vssd vssd vccd vccd _1315_/A sky130_fd_sc_hd__buf_2
Xinput311 la_oenb_mprj[30] vssd vssd vccd vccd _1335_/A sky130_fd_sc_hd__clkbuf_1
Xinput322 la_oenb_mprj[40] vssd vssd vccd vccd _1355_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input331_A la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput333 la_oenb_mprj[50] vssd vssd vccd vccd _1375_/A sky130_fd_sc_hd__buf_2
Xinput344 la_oenb_mprj[60] vssd vssd vccd vccd _1395_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1243__A_N _1499_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input429_A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput355 la_oenb_mprj[70] vssd vssd vccd vccd _1415_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput366 la_oenb_mprj[80] vssd vssd vccd vccd _1435_/A sky130_fd_sc_hd__buf_4
XANTENNA_input25_A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput377 la_oenb_mprj[90] vssd vssd vccd vccd _1455_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput388 mprj_adr_o_core[0] vssd vssd vccd vccd _0891_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_40_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput399 mprj_adr_o_core[1] vssd vssd vccd vccd _0893_/B sky130_fd_sc_hd__buf_6
XFILLER_21_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__0989__B _0989_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput807 _1404_/X vssd vssd vccd vccd la_oenb_core[64] sky130_fd_sc_hd__buf_12
XFILLER_49_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput818 _1424_/X vssd vssd vccd vccd la_oenb_core[74] sky130_fd_sc_hd__buf_12
XANTENNA_output550_A _1146_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput829 _1444_/X vssd vssd vccd vccd la_oenb_core[84] sky130_fd_sc_hd__buf_12
XANTENNA_output648_A _0481_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__1166__A _1166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0522_ _0522_/A vssd vssd vccd vccd _0522_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] _0732_/X vssd vssd vccd vccd _0507_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_39_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_1005_ _1005_/A _1005_/B vssd vssd vccd vccd _1006_/A sky130_fd_sc_hd__and2_4
XFILLER_35_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__0899__B _0899_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1076__A _1076_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1523__B _1523_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input281_A la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input379_A la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3807 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput130 la_data_out_mprj[99] vssd vssd vccd vccd _1217_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_24_2863 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput141 la_iena_mprj[108] vssd vssd vccd vccd _0823_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput152 la_iena_mprj[118] vssd vssd vccd vccd _0843_/B sky130_fd_sc_hd__buf_2
XFILLER_4_2957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__1433__B _1433_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput163 la_iena_mprj[12] vssd vssd vccd vccd _0631_/B sky130_fd_sc_hd__clkbuf_1
Xinput174 la_iena_mprj[22] vssd vssd vccd vccd _0651_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput185 la_iena_mprj[32] vssd vssd vccd vccd _0671_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput196 la_iena_mprj[42] vssd vssd vccd vccd _0691_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output598_A _0551_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__1139__A_N _1395_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output932_A _1010_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput604 _0556_/Y vssd vssd vccd vccd la_data_in_mprj[111] sky130_fd_sc_hd__buf_12
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput615 _0566_/Y vssd vssd vccd vccd la_data_in_mprj[121] sky130_fd_sc_hd__buf_12
XFILLER_44_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput626 _1549_/Y vssd vssd vccd vccd la_data_in_mprj[16] sky130_fd_sc_hd__buf_12
XFILLER_47_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput637 _0471_/Y vssd vssd vccd vccd la_data_in_mprj[26] sky130_fd_sc_hd__buf_12
Xoutput648 _0481_/Y vssd vssd vccd vccd la_data_in_mprj[36] sky130_fd_sc_hd__buf_12
XFILLER_29_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput659 _0491_/Y vssd vssd vccd vccd la_data_in_mprj[46] sky130_fd_sc_hd__buf_12
XFILLER_45_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_0505_ _0505_/A vssd vssd vccd vccd _0505_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_1485_ _1485_/A _1485_/B vssd vssd vccd vccd _1486_/A sky130_fd_sc_hd__and2_1
XFILLER_42_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
.ends

