magic
tech sky130A
magscale 1 2
timestamp 1659794613
<< viali >>
rect 3801 11305 3835 11339
rect 8033 11305 8067 11339
rect 9229 11305 9263 11339
rect 6929 11169 6963 11203
rect 7297 11169 7331 11203
rect 7573 11169 7607 11203
rect 8309 11169 8343 11203
rect 8493 11169 8527 11203
rect 9413 11169 9447 11203
rect 3065 11101 3099 11135
rect 4077 11101 4111 11135
rect 4353 11101 4387 11135
rect 5181 11101 5215 11135
rect 6009 11101 6043 11135
rect 6653 11101 6687 11135
rect 7941 11101 7975 11135
rect 8861 11101 8895 11135
rect 3341 11033 3375 11067
rect 3617 11033 3651 11067
rect 4261 11033 4295 11067
rect 4813 11033 4847 11067
rect 2973 10965 3007 10999
rect 4629 10965 4663 10999
rect 5917 10965 5951 10999
rect 6193 10965 6227 10999
rect 6377 10965 6411 10999
rect 7849 10965 7883 10999
rect 9045 10965 9079 10999
rect 5365 10693 5399 10727
rect 7941 10693 7975 10727
rect 2789 10625 2823 10659
rect 4629 10625 4663 10659
rect 5549 10625 5583 10659
rect 5825 10625 5859 10659
rect 6285 10625 6319 10659
rect 6837 10625 6871 10659
rect 7021 10625 7055 10659
rect 7481 10625 7515 10659
rect 7665 10625 7699 10659
rect 2053 10557 2087 10591
rect 3157 10557 3191 10591
rect 6561 10557 6595 10591
rect 5733 10489 5767 10523
rect 2697 10421 2731 10455
rect 5189 10421 5223 10455
rect 5917 10421 5951 10455
rect 6377 10421 6411 10455
rect 7113 10421 7147 10455
rect 7389 10421 7423 10455
rect 9413 10421 9447 10455
rect 4721 10217 4755 10251
rect 5273 10149 5307 10183
rect 1869 10081 1903 10115
rect 3341 10081 3375 10115
rect 4169 10081 4203 10115
rect 4813 10081 4847 10115
rect 5457 10081 5491 10115
rect 1593 10013 1627 10047
rect 4537 10013 4571 10047
rect 5089 10013 5123 10047
rect 5825 10013 5859 10047
rect 7297 10013 7331 10047
rect 8125 10013 8159 10047
rect 8493 10013 8527 10047
rect 8953 10013 8987 10047
rect 9137 10013 9171 10047
rect 8309 9945 8343 9979
rect 8769 9945 8803 9979
rect 9229 9945 9263 9979
rect 9413 9945 9447 9979
rect 3617 9877 3651 9911
rect 4445 9877 4479 9911
rect 7861 9877 7895 9911
rect 5917 9673 5951 9707
rect 5745 9605 5779 9639
rect 3249 9537 3283 9571
rect 3341 9537 3375 9571
rect 5181 9537 5215 9571
rect 7021 9537 7055 9571
rect 8861 9537 8895 9571
rect 1501 9469 1535 9503
rect 2973 9469 3007 9503
rect 3709 9469 3743 9503
rect 6193 9469 6227 9503
rect 6745 9469 6779 9503
rect 7389 9469 7423 9503
rect 9425 9333 9459 9367
rect 2329 9129 2363 9163
rect 2789 9129 2823 9163
rect 4629 9129 4663 9163
rect 8217 9129 8251 9163
rect 9505 9129 9539 9163
rect 3433 9061 3467 9095
rect 8493 9061 8527 9095
rect 6377 8993 6411 9027
rect 6469 8993 6503 9027
rect 8861 8925 8895 8959
rect 3065 8857 3099 8891
rect 3249 8857 3283 8891
rect 3801 8857 3835 8891
rect 3985 8857 4019 8891
rect 4169 8857 4203 8891
rect 4261 8857 4295 8891
rect 6101 8857 6135 8891
rect 6745 8857 6779 8891
rect 2605 8789 2639 8823
rect 2973 8789 3007 8823
rect 3709 8789 3743 8823
rect 9045 8789 9079 8823
rect 9321 8789 9355 8823
rect 8033 8585 8067 8619
rect 1777 8517 1811 8551
rect 6193 8517 6227 8551
rect 8953 8517 8987 8551
rect 6009 8449 6043 8483
rect 8585 8449 8619 8483
rect 9137 8449 9171 8483
rect 9229 8449 9263 8483
rect 1501 8381 1535 8415
rect 3249 8381 3283 8415
rect 3985 8381 4019 8415
rect 4721 8313 4755 8347
rect 7481 8313 7515 8347
rect 8769 8313 8803 8347
rect 9413 8313 9447 8347
rect 3433 8245 3467 8279
rect 2789 8041 2823 8075
rect 4721 8041 4755 8075
rect 9413 8041 9447 8075
rect 3709 7973 3743 8007
rect 9045 7973 9079 8007
rect 6101 7905 6135 7939
rect 9321 7905 9355 7939
rect 3065 7837 3099 7871
rect 3617 7837 3651 7871
rect 4077 7837 4111 7871
rect 6469 7837 6503 7871
rect 7941 7837 7975 7871
rect 3249 7769 3283 7803
rect 6009 7769 6043 7803
rect 8505 7769 8539 7803
rect 2973 7701 3007 7735
rect 3433 7701 3467 7735
rect 8861 7701 8895 7735
rect 2513 7497 2547 7531
rect 9413 7497 9447 7531
rect 6193 7429 6227 7463
rect 7941 7429 7975 7463
rect 9045 7429 9079 7463
rect 2789 7361 2823 7395
rect 3157 7361 3191 7395
rect 4629 7361 4663 7395
rect 5549 7361 5583 7395
rect 9229 7361 9263 7395
rect 5825 7293 5859 7327
rect 8585 7293 8619 7327
rect 8953 7293 8987 7327
rect 5193 7225 5227 7259
rect 2697 7157 2731 7191
rect 5917 7157 5951 7191
rect 8033 7157 8067 7191
rect 1764 6953 1798 6987
rect 7489 6953 7523 6987
rect 9505 6885 9539 6919
rect 3249 6817 3283 6851
rect 4169 6817 4203 6851
rect 8953 6817 8987 6851
rect 1501 6749 1535 6783
rect 4353 6749 4387 6783
rect 4813 6749 4847 6783
rect 5089 6749 5123 6783
rect 5457 6749 5491 6783
rect 6929 6749 6963 6783
rect 7849 6749 7883 6783
rect 8125 6749 8159 6783
rect 8585 6749 8619 6783
rect 4629 6681 4663 6715
rect 7757 6681 7791 6715
rect 8309 6681 8343 6715
rect 9045 6681 9079 6715
rect 3617 6613 3651 6647
rect 9137 6613 9171 6647
rect 2237 6409 2271 6443
rect 8125 6409 8159 6443
rect 8953 6409 8987 6443
rect 9045 6409 9079 6443
rect 2053 6341 2087 6375
rect 2421 6341 2455 6375
rect 5365 6341 5399 6375
rect 6469 6341 6503 6375
rect 8309 6341 8343 6375
rect 8769 6341 8803 6375
rect 9137 6341 9171 6375
rect 2697 6273 2731 6307
rect 4629 6273 4663 6307
rect 6193 6273 6227 6307
rect 8493 6273 8527 6307
rect 8677 6273 8711 6307
rect 2605 6205 2639 6239
rect 2789 6205 2823 6239
rect 3157 6205 3191 6239
rect 5917 6205 5951 6239
rect 7941 6205 7975 6239
rect 9321 6137 9355 6171
rect 5193 6069 5227 6103
rect 9413 6069 9447 6103
rect 1856 5865 1890 5899
rect 3985 5865 4019 5899
rect 5917 5865 5951 5899
rect 8493 5865 8527 5899
rect 8401 5797 8435 5831
rect 1593 5729 1627 5763
rect 4445 5729 4479 5763
rect 6193 5729 6227 5763
rect 6469 5729 6503 5763
rect 7941 5729 7975 5763
rect 8861 5729 8895 5763
rect 4169 5661 4203 5695
rect 1501 5593 1535 5627
rect 3709 5593 3743 5627
rect 3893 5593 3927 5627
rect 8953 5593 8987 5627
rect 9505 5593 9539 5627
rect 3341 5525 3375 5559
rect 8217 5525 8251 5559
rect 8309 5321 8343 5355
rect 8125 5253 8159 5287
rect 6009 5185 6043 5219
rect 9045 5185 9079 5219
rect 9229 5185 9263 5219
rect 3341 5117 3375 5151
rect 3617 5117 3651 5151
rect 5273 5117 5307 5151
rect 5825 5117 5859 5151
rect 6285 5117 6319 5151
rect 7757 5117 7791 5151
rect 8861 5117 8895 5151
rect 5089 4981 5123 5015
rect 9321 4981 9355 5015
rect 5089 4777 5123 4811
rect 9413 4777 9447 4811
rect 5365 4641 5399 4675
rect 5733 4641 5767 4675
rect 6285 4641 6319 4675
rect 3341 4573 3375 4607
rect 5457 4573 5491 4607
rect 6561 4573 6595 4607
rect 6929 4573 6963 4607
rect 8401 4573 8435 4607
rect 9321 4573 9355 4607
rect 3617 4505 3651 4539
rect 8965 4505 8999 4539
rect 9229 4437 9263 4471
rect 6377 4233 6411 4267
rect 3341 4097 3375 4131
rect 3525 4097 3559 4131
rect 5365 4097 5399 4131
rect 6285 4097 6319 4131
rect 8125 4097 8159 4131
rect 9413 4097 9447 4131
rect 3893 4029 3927 4063
rect 6561 4029 6595 4063
rect 8309 4029 8343 4063
rect 8861 4029 8895 4063
rect 6101 3961 6135 3995
rect 8033 3961 8067 3995
rect 5925 3893 5959 3927
rect 9137 3893 9171 3927
rect 9229 3893 9263 3927
rect 5457 3689 5491 3723
rect 5825 3689 5859 3723
rect 3433 3553 3467 3587
rect 7205 3553 7239 3587
rect 5089 3485 5123 3519
rect 5733 3485 5767 3519
rect 6193 3485 6227 3519
rect 6745 3485 6779 3519
rect 6837 3485 6871 3519
rect 8677 3485 8711 3519
rect 5181 3417 5215 3451
rect 5365 3417 5399 3451
rect 6377 3417 6411 3451
rect 6561 3417 6595 3451
rect 9241 3417 9275 3451
rect 8861 3349 8895 3383
rect 9413 3349 9447 3383
rect 4169 3145 4203 3179
rect 8125 3145 8159 3179
rect 8401 3145 8435 3179
rect 8953 3145 8987 3179
rect 9413 3145 9447 3179
rect 3433 3077 3467 3111
rect 7481 3077 7515 3111
rect 8493 3077 8527 3111
rect 3525 3009 3559 3043
rect 4445 3009 4479 3043
rect 6469 3009 6503 3043
rect 7297 3009 7331 3043
rect 9045 3009 9079 3043
rect 4629 2941 4663 2975
rect 4997 2941 5031 2975
rect 7033 2941 7067 2975
rect 7573 2941 7607 2975
rect 7941 2941 7975 2975
rect 8861 2941 8895 2975
rect 4353 2805 4387 2839
rect 4813 2601 4847 2635
rect 5181 2601 5215 2635
rect 6101 2601 6135 2635
rect 6561 2601 6595 2635
rect 7021 2601 7055 2635
rect 7941 2601 7975 2635
rect 9045 2601 9079 2635
rect 9229 2601 9263 2635
rect 5273 2533 5307 2567
rect 5457 2533 5491 2567
rect 6377 2533 6411 2567
rect 6745 2533 6779 2567
rect 7205 2533 7239 2567
rect 8493 2533 8527 2567
rect 3985 2465 4019 2499
rect 9505 2465 9539 2499
rect 3433 2397 3467 2431
rect 3617 2397 3651 2431
rect 4077 2397 4111 2431
rect 4353 2397 4387 2431
rect 4905 2397 4939 2431
rect 5917 2397 5951 2431
rect 6193 2397 6227 2431
rect 6929 2397 6963 2431
rect 7573 2397 7607 2431
rect 7849 2397 7883 2431
rect 8125 2397 8159 2431
rect 8677 2397 8711 2431
rect 4169 2329 4203 2363
rect 4537 2329 4571 2363
rect 8309 2329 8343 2363
rect 9091 2329 9125 2363
rect 5741 2057 5775 2091
rect 6009 2057 6043 2091
rect 8309 2057 8343 2091
rect 8585 2057 8619 2091
rect 8769 2057 8803 2091
rect 9321 2057 9355 2091
rect 7297 1989 7331 2023
rect 7941 1989 7975 2023
rect 9413 1989 9447 2023
rect 3341 1921 3375 1955
rect 5181 1921 5215 1955
rect 3709 1853 3743 1887
rect 9137 1853 9171 1887
rect 8953 1785 8987 1819
rect 5365 1513 5399 1547
rect 9413 1513 9447 1547
rect 5273 1445 5307 1479
rect 5089 1309 5123 1343
rect 3801 1173 3835 1207
<< obsli1 >>
rect 0 12986 853 13014
rect 0 12969 9963 12986
rect 0 11481 33962 12969
rect 0 6005 853 11481
rect 0 5899 3359 6005
rect 0 5865 1856 5899
rect 1890 5865 3359 5899
rect 0 5763 3359 5865
rect 0 5729 1593 5763
rect 1627 5729 3359 5763
rect 0 5627 3359 5729
rect 0 5593 1501 5627
rect 1535 5593 3359 5627
rect 0 5559 3359 5593
rect 0 5525 3341 5559
rect 0 5151 3359 5525
rect 0 5117 3341 5151
rect 0 4607 3359 5117
rect 0 4573 3341 4607
rect 0 4131 3359 4573
rect 0 4097 3341 4131
rect 0 1955 3359 4097
rect 0 1921 3341 1955
rect 0 0 3359 1921
rect 9800 1048 33962 11481
rect 3366 0 33962 1048
<< metal1 >>
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 7566 11450
rect 7618 11398 7630 11450
rect 7682 11398 7694 11450
rect 7746 11398 7758 11450
rect 7810 11398 7822 11450
rect 7874 11398 9844 11450
rect 920 11376 9844 11398
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 1820 11308 3801 11336
rect 1820 11296 1826 11308
rect 3789 11305 3801 11308
rect 3835 11336 3847 11339
rect 4338 11336 4344 11348
rect 3835 11308 4344 11336
rect 3835 11305 3847 11308
rect 3789 11299 3847 11305
rect 4338 11296 4344 11308
rect 4396 11296 4402 11348
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 8021 11339 8079 11345
rect 8021 11336 8033 11339
rect 6972 11308 8033 11336
rect 6972 11296 6978 11308
rect 8021 11305 8033 11308
rect 8067 11336 8079 11339
rect 8110 11336 8116 11348
rect 8067 11308 8116 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8110 11296 8116 11308
rect 8168 11336 8174 11348
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 8168 11308 9229 11336
rect 8168 11296 8174 11308
rect 9217 11305 9229 11308
rect 9263 11305 9275 11339
rect 9217 11299 9275 11305
rect 4798 11200 4804 11212
rect 3068 11172 4804 11200
rect 3068 11141 3096 11172
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 6362 11160 6368 11212
rect 6420 11200 6426 11212
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 6420 11172 6929 11200
rect 6420 11160 6426 11172
rect 6917 11169 6929 11172
rect 6963 11200 6975 11203
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 6963 11172 7297 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 7285 11169 7297 11172
rect 7331 11200 7343 11203
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7331 11172 7573 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 7561 11169 7573 11172
rect 7607 11200 7619 11203
rect 8018 11200 8024 11212
rect 7607 11172 8024 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 8018 11160 8024 11172
rect 8076 11200 8082 11212
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 8076 11172 8309 11200
rect 8076 11160 8082 11172
rect 8297 11169 8309 11172
rect 8343 11200 8355 11203
rect 8481 11203 8539 11209
rect 8481 11200 8493 11203
rect 8343 11172 8493 11200
rect 8343 11169 8355 11172
rect 8297 11163 8355 11169
rect 8481 11169 8493 11172
rect 8527 11200 8539 11203
rect 9401 11203 9459 11209
rect 9401 11200 9413 11203
rect 8527 11172 9413 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 9401 11169 9413 11172
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 3053 11095 3111 11101
rect 3620 11104 4077 11132
rect 3142 11024 3148 11076
rect 3200 11064 3206 11076
rect 3620 11073 3648 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4338 11132 4344 11144
rect 4299 11104 4344 11132
rect 4065 11095 4123 11101
rect 3329 11067 3387 11073
rect 3329 11064 3341 11067
rect 3200 11036 3341 11064
rect 3200 11024 3206 11036
rect 3329 11033 3341 11036
rect 3375 11064 3387 11067
rect 3605 11067 3663 11073
rect 3605 11064 3617 11067
rect 3375 11036 3617 11064
rect 3375 11033 3387 11036
rect 3329 11027 3387 11033
rect 3605 11033 3617 11036
rect 3651 11033 3663 11067
rect 3605 11027 3663 11033
rect 2958 10996 2964 11008
rect 2919 10968 2964 10996
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 4080 10996 4108 11095
rect 4338 11092 4344 11104
rect 4396 11132 4402 11144
rect 5169 11135 5227 11141
rect 5169 11132 5181 11135
rect 4396 11104 5181 11132
rect 4396 11092 4402 11104
rect 5169 11101 5181 11104
rect 5215 11132 5227 11135
rect 5350 11132 5356 11144
rect 5215 11104 5356 11132
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 5350 11092 5356 11104
rect 5408 11092 5414 11144
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 4246 11064 4252 11076
rect 4207 11036 4252 11064
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 4801 11067 4859 11073
rect 4801 11064 4813 11067
rect 4356 11036 4813 11064
rect 4356 10996 4384 11036
rect 4801 11033 4813 11036
rect 4847 11033 4859 11067
rect 6012 11064 6040 11095
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 6641 11135 6699 11141
rect 6641 11132 6653 11135
rect 6144 11104 6653 11132
rect 6144 11092 6150 11104
rect 6641 11101 6653 11104
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 6880 11104 7941 11132
rect 6880 11092 6886 11104
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 8849 11135 8907 11141
rect 8849 11101 8861 11135
rect 8895 11101 8907 11135
rect 8849 11095 8907 11101
rect 7006 11064 7012 11076
rect 6012 11036 7012 11064
rect 4801 11027 4859 11033
rect 7006 11024 7012 11036
rect 7064 11064 7070 11076
rect 8864 11064 8892 11095
rect 16574 11064 16580 11076
rect 7064 11036 8892 11064
rect 9048 11036 16580 11064
rect 7064 11024 7070 11036
rect 4080 10968 4384 10996
rect 4430 10956 4436 11008
rect 4488 10996 4494 11008
rect 4617 10999 4675 11005
rect 4617 10996 4629 10999
rect 4488 10968 4629 10996
rect 4488 10956 4494 10968
rect 4617 10965 4629 10968
rect 4663 10965 4675 10999
rect 4617 10959 4675 10965
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 5905 10999 5963 11005
rect 5905 10996 5917 10999
rect 5592 10968 5917 10996
rect 5592 10956 5598 10968
rect 5905 10965 5917 10968
rect 5951 10965 5963 10999
rect 5905 10959 5963 10965
rect 6086 10956 6092 11008
rect 6144 10996 6150 11008
rect 6181 10999 6239 11005
rect 6181 10996 6193 10999
rect 6144 10968 6193 10996
rect 6144 10956 6150 10968
rect 6181 10965 6193 10968
rect 6227 10965 6239 10999
rect 6362 10996 6368 11008
rect 6323 10968 6368 10996
rect 6181 10959 6239 10965
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 9048 11005 9076 11036
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 7837 10999 7895 11005
rect 7837 10996 7849 10999
rect 7708 10968 7849 10996
rect 7708 10956 7714 10968
rect 7837 10965 7849 10968
rect 7883 10965 7895 10999
rect 7837 10959 7895 10965
rect 9033 10999 9091 11005
rect 9033 10965 9045 10999
rect 9079 10965 9091 10999
rect 9033 10959 9091 10965
rect 920 10906 9844 10928
rect 920 10854 3816 10906
rect 3868 10854 3880 10906
rect 3932 10854 3944 10906
rect 3996 10854 4008 10906
rect 4060 10854 4072 10906
rect 4124 10854 8816 10906
rect 8868 10854 8880 10906
rect 8932 10854 8944 10906
rect 8996 10854 9008 10906
rect 9060 10854 9072 10906
rect 9124 10854 9844 10906
rect 920 10832 9844 10854
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 7006 10792 7012 10804
rect 4856 10764 7012 10792
rect 4856 10752 4862 10764
rect 4706 10724 4712 10736
rect 4278 10696 4712 10724
rect 4706 10684 4712 10696
rect 4764 10684 4770 10736
rect 5350 10724 5356 10736
rect 5311 10696 5356 10724
rect 5350 10684 5356 10696
rect 5408 10684 5414 10736
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 2958 10656 2964 10668
rect 2823 10628 2964 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 4617 10659 4675 10665
rect 4617 10656 4629 10659
rect 4396 10628 4629 10656
rect 4396 10616 4402 10628
rect 4617 10625 4629 10628
rect 4663 10625 4675 10659
rect 4617 10619 4675 10625
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 5537 10659 5595 10665
rect 5537 10656 5549 10659
rect 5316 10628 5549 10656
rect 5316 10616 5322 10628
rect 5537 10625 5549 10628
rect 5583 10625 5595 10659
rect 5736 10658 5764 10764
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 8018 10752 8024 10804
rect 8076 10792 8082 10804
rect 8076 10764 8340 10792
rect 8076 10752 8082 10764
rect 7024 10724 7052 10752
rect 7929 10727 7987 10733
rect 7024 10696 7512 10724
rect 5813 10659 5871 10665
rect 5813 10658 5825 10659
rect 5736 10630 5825 10658
rect 5537 10619 5595 10625
rect 5813 10625 5825 10630
rect 5859 10625 5871 10659
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 5813 10619 5871 10625
rect 5920 10628 6285 10656
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 2041 10591 2099 10597
rect 2041 10588 2053 10591
rect 1636 10560 2053 10588
rect 1636 10548 1642 10560
rect 2041 10557 2053 10560
rect 2087 10557 2099 10591
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 2041 10551 2099 10557
rect 2700 10560 3157 10588
rect 1762 10412 1768 10464
rect 1820 10452 1826 10464
rect 2700 10461 2728 10560
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 5552 10588 5580 10619
rect 5920 10588 5948 10628
rect 6273 10625 6285 10628
rect 6319 10656 6331 10659
rect 6362 10656 6368 10668
rect 6319 10628 6368 10656
rect 6319 10625 6331 10628
rect 6273 10619 6331 10625
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 7484 10665 7512 10696
rect 7929 10693 7941 10727
rect 7975 10724 7987 10727
rect 8202 10724 8208 10736
rect 7975 10696 8208 10724
rect 7975 10693 7987 10696
rect 7929 10687 7987 10693
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 8312 10724 8340 10764
rect 8312 10696 8418 10724
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6748 10628 6837 10656
rect 5552 10560 5948 10588
rect 3145 10551 3203 10557
rect 5718 10520 5724 10532
rect 5679 10492 5724 10520
rect 5718 10480 5724 10492
rect 5776 10480 5782 10532
rect 5920 10520 5948 10560
rect 6086 10548 6092 10600
rect 6144 10588 6150 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 6144 10560 6561 10588
rect 6144 10548 6150 10560
rect 6549 10557 6561 10560
rect 6595 10588 6607 10591
rect 6748 10588 6776 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10625 7527 10659
rect 7650 10656 7656 10668
rect 7611 10628 7656 10656
rect 7469 10619 7527 10625
rect 6595 10560 6776 10588
rect 6595 10557 6607 10560
rect 6549 10551 6607 10557
rect 7024 10520 7052 10619
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 7466 10520 7472 10532
rect 5920 10492 7472 10520
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 2685 10455 2743 10461
rect 2685 10452 2697 10455
rect 1820 10424 2697 10452
rect 1820 10412 1826 10424
rect 2685 10421 2697 10424
rect 2731 10421 2743 10455
rect 5166 10452 5172 10464
rect 5224 10461 5230 10464
rect 5135 10424 5172 10452
rect 2685 10415 2743 10421
rect 5166 10412 5172 10424
rect 5224 10415 5235 10461
rect 5902 10452 5908 10464
rect 5863 10424 5908 10452
rect 5224 10412 5230 10415
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 6362 10452 6368 10464
rect 6323 10424 6368 10452
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 7098 10452 7104 10464
rect 7059 10424 7104 10452
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 7190 10412 7196 10464
rect 7248 10452 7254 10464
rect 7377 10455 7435 10461
rect 7377 10452 7389 10455
rect 7248 10424 7389 10452
rect 7248 10412 7254 10424
rect 7377 10421 7389 10424
rect 7423 10421 7435 10455
rect 7377 10415 7435 10421
rect 9401 10455 9459 10461
rect 9401 10421 9413 10455
rect 9447 10452 9459 10455
rect 16574 10452 16580 10464
rect 9447 10424 16580 10452
rect 9447 10421 9459 10424
rect 9401 10415 9459 10421
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 7566 10362
rect 7618 10310 7630 10362
rect 7682 10310 7694 10362
rect 7746 10310 7758 10362
rect 7810 10310 7822 10362
rect 7874 10310 9844 10362
rect 920 10288 9844 10310
rect 4706 10248 4712 10260
rect 4667 10220 4712 10248
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8168 10220 9168 10248
rect 8168 10208 8174 10220
rect 3142 10140 3148 10192
rect 3200 10180 3206 10192
rect 5258 10180 5264 10192
rect 3200 10152 5264 10180
rect 3200 10140 3206 10152
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10112 1915 10115
rect 3329 10115 3387 10121
rect 1903 10084 3280 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 1486 10004 1492 10056
rect 1544 10044 1550 10056
rect 1581 10047 1639 10053
rect 1581 10044 1593 10047
rect 1544 10016 1593 10044
rect 1544 10004 1550 10016
rect 1581 10013 1593 10016
rect 1627 10013 1639 10047
rect 3142 10044 3148 10056
rect 2990 10016 3148 10044
rect 1581 10007 1639 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3252 9976 3280 10084
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 4157 10115 4215 10121
rect 4157 10112 4169 10115
rect 3375 10084 4169 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 4157 10081 4169 10084
rect 4203 10081 4215 10115
rect 4157 10075 4215 10081
rect 4430 10072 4436 10124
rect 4488 10112 4494 10124
rect 4801 10115 4859 10121
rect 4801 10112 4813 10115
rect 4488 10084 4813 10112
rect 4488 10072 4494 10084
rect 4801 10081 4813 10084
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 4706 10044 4712 10056
rect 4571 10016 4712 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 5092 10053 5120 10152
rect 5258 10140 5264 10152
rect 5316 10140 5322 10192
rect 5445 10115 5503 10121
rect 5445 10081 5457 10115
rect 5491 10112 5503 10115
rect 5534 10112 5540 10124
rect 5491 10084 5540 10112
rect 5491 10081 5503 10084
rect 5445 10075 5503 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 8018 10072 8024 10124
rect 8076 10112 8082 10124
rect 8076 10084 8340 10112
rect 8076 10072 8082 10084
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10013 5135 10047
rect 5810 10044 5816 10056
rect 5077 10007 5135 10013
rect 5184 10016 5816 10044
rect 5184 9976 5212 10016
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 7098 10004 7104 10056
rect 7156 10044 7162 10056
rect 7285 10047 7343 10053
rect 7285 10044 7297 10047
rect 7156 10016 7297 10044
rect 7156 10004 7162 10016
rect 7285 10013 7297 10016
rect 7331 10013 7343 10047
rect 8110 10044 8116 10056
rect 8071 10016 8116 10044
rect 7285 10007 7343 10013
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 8312 10044 8340 10084
rect 9140 10053 9168 10220
rect 8481 10047 8539 10053
rect 8481 10044 8493 10047
rect 8312 10016 8493 10044
rect 8481 10013 8493 10016
rect 8527 10044 8539 10047
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8527 10016 8953 10044
rect 8527 10013 8539 10016
rect 8481 10007 8539 10013
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 3252 9948 5212 9976
rect 6362 9936 6368 9988
rect 6420 9936 6426 9988
rect 8294 9976 8300 9988
rect 8255 9948 8300 9976
rect 8294 9936 8300 9948
rect 8352 9936 8358 9988
rect 8662 9936 8668 9988
rect 8720 9976 8726 9988
rect 8757 9979 8815 9985
rect 8757 9976 8769 9979
rect 8720 9948 8769 9976
rect 8720 9936 8726 9948
rect 8757 9945 8769 9948
rect 8803 9945 8815 9979
rect 8956 9976 8984 10007
rect 9217 9979 9275 9985
rect 9217 9976 9229 9979
rect 8956 9948 9229 9976
rect 8757 9939 8815 9945
rect 9217 9945 9229 9948
rect 9263 9976 9275 9979
rect 9401 9979 9459 9985
rect 9401 9976 9413 9979
rect 9263 9948 9413 9976
rect 9263 9945 9275 9948
rect 9217 9939 9275 9945
rect 9401 9945 9413 9948
rect 9447 9945 9459 9979
rect 9401 9939 9459 9945
rect 3605 9911 3663 9917
rect 3605 9877 3617 9911
rect 3651 9908 3663 9911
rect 3694 9908 3700 9920
rect 3651 9880 3700 9908
rect 3651 9877 3663 9880
rect 3605 9871 3663 9877
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 4433 9911 4491 9917
rect 4433 9908 4445 9911
rect 4212 9880 4445 9908
rect 4212 9868 4218 9880
rect 4433 9877 4445 9880
rect 4479 9877 4491 9911
rect 4433 9871 4491 9877
rect 7849 9911 7907 9917
rect 7849 9877 7861 9911
rect 7895 9908 7907 9911
rect 8570 9908 8576 9920
rect 7895 9880 8576 9908
rect 7895 9877 7907 9880
rect 7849 9871 7907 9877
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 920 9818 9844 9840
rect 920 9766 3816 9818
rect 3868 9766 3880 9818
rect 3932 9766 3944 9818
rect 3996 9766 4008 9818
rect 4060 9766 4072 9818
rect 4124 9766 8816 9818
rect 8868 9766 8880 9818
rect 8932 9766 8944 9818
rect 8996 9766 9008 9818
rect 9060 9766 9072 9818
rect 9124 9766 9844 9818
rect 920 9744 9844 9766
rect 1486 9664 1492 9716
rect 1544 9704 1550 9716
rect 1544 9676 2728 9704
rect 1544 9664 1550 9676
rect 2314 9596 2320 9648
rect 2372 9596 2378 9648
rect 2700 9636 2728 9676
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 5905 9707 5963 9713
rect 5905 9704 5917 9707
rect 5316 9676 5917 9704
rect 5316 9664 5322 9676
rect 5905 9673 5917 9676
rect 5951 9673 5963 9707
rect 5905 9667 5963 9673
rect 7466 9664 7472 9716
rect 7524 9704 7530 9716
rect 8110 9704 8116 9716
rect 7524 9676 8116 9704
rect 7524 9664 7530 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 2700 9608 3280 9636
rect 3252 9577 3280 9608
rect 4246 9596 4252 9648
rect 4304 9596 4310 9648
rect 5733 9639 5791 9645
rect 5733 9605 5745 9639
rect 5779 9636 5791 9639
rect 5779 9608 6914 9636
rect 5779 9605 5791 9608
rect 5733 9599 5791 9605
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 3329 9571 3387 9577
rect 3329 9537 3341 9571
rect 3375 9568 3387 9571
rect 5169 9571 5227 9577
rect 3375 9540 3832 9568
rect 3375 9537 3387 9540
rect 3329 9531 3387 9537
rect 1489 9503 1547 9509
rect 1489 9469 1501 9503
rect 1535 9500 1547 9503
rect 1578 9500 1584 9512
rect 1535 9472 1584 9500
rect 1535 9469 1547 9472
rect 1489 9463 1547 9469
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9500 3019 9503
rect 3694 9500 3700 9512
rect 3007 9472 3700 9500
rect 3007 9469 3019 9472
rect 2961 9463 3019 9469
rect 3694 9460 3700 9472
rect 3752 9460 3758 9512
rect 3804 9500 3832 9540
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5215 9540 5764 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5736 9512 5764 9540
rect 4154 9500 4160 9512
rect 3804 9472 4160 9500
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 5718 9460 5724 9512
rect 5776 9460 5782 9512
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 6181 9503 6239 9509
rect 6181 9500 6193 9503
rect 5868 9472 6193 9500
rect 5868 9460 5874 9472
rect 6181 9469 6193 9472
rect 6227 9469 6239 9503
rect 6730 9500 6736 9512
rect 6691 9472 6736 9500
rect 6181 9463 6239 9469
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 6086 9432 6092 9444
rect 5828 9404 6092 9432
rect 934 9324 940 9376
rect 992 9364 998 9376
rect 5828 9364 5856 9404
rect 6086 9392 6092 9404
rect 6144 9392 6150 9444
rect 992 9336 5856 9364
rect 6886 9364 6914 9608
rect 8294 9596 8300 9648
rect 8352 9596 8358 9648
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9568 7067 9571
rect 7190 9568 7196 9580
rect 7055 9540 7196 9568
rect 7055 9537 7067 9540
rect 7009 9531 7067 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8720 9540 8861 9568
rect 8720 9528 8726 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 7377 9503 7435 9509
rect 7377 9469 7389 9503
rect 7423 9500 7435 9503
rect 8018 9500 8024 9512
rect 7423 9472 8024 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8478 9364 8484 9376
rect 6886 9336 8484 9364
rect 992 9324 998 9336
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 9413 9367 9471 9373
rect 9413 9333 9425 9367
rect 9459 9364 9471 9367
rect 9582 9364 9588 9376
rect 9459 9336 9588 9364
rect 9459 9333 9471 9336
rect 9413 9327 9471 9333
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 7566 9274
rect 7618 9222 7630 9274
rect 7682 9222 7694 9274
rect 7746 9222 7758 9274
rect 7810 9222 7822 9274
rect 7874 9222 9844 9274
rect 920 9200 9844 9222
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 2317 9163 2375 9169
rect 2317 9160 2329 9163
rect 2004 9132 2329 9160
rect 2004 9120 2010 9132
rect 2317 9129 2329 9132
rect 2363 9129 2375 9163
rect 2317 9123 2375 9129
rect 2332 8888 2360 9123
rect 2406 9120 2412 9172
rect 2464 9160 2470 9172
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2464 9132 2789 9160
rect 2464 9120 2470 9132
rect 2777 9129 2789 9132
rect 2823 9160 2835 9163
rect 2958 9160 2964 9172
rect 2823 9132 2964 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 4617 9163 4675 9169
rect 4617 9129 4629 9163
rect 4663 9160 4675 9163
rect 6730 9160 6736 9172
rect 4663 9132 6736 9160
rect 4663 9129 4675 9132
rect 4617 9123 4675 9129
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 8202 9160 8208 9172
rect 8163 9132 8208 9160
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 9490 9160 9496 9172
rect 9451 9132 9496 9160
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 3421 9095 3479 9101
rect 3421 9061 3433 9095
rect 3467 9092 3479 9095
rect 4338 9092 4344 9104
rect 3467 9064 4344 9092
rect 3467 9061 3479 9064
rect 3421 9055 3479 9061
rect 4338 9052 4344 9064
rect 4396 9052 4402 9104
rect 8481 9095 8539 9101
rect 8481 9061 8493 9095
rect 8527 9092 8539 9095
rect 8527 9064 16574 9092
rect 8527 9061 8539 9064
rect 8481 9055 8539 9061
rect 4430 9024 4436 9036
rect 2884 8996 4436 9024
rect 2884 8888 2912 8996
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 6365 9027 6423 9033
rect 6365 8993 6377 9027
rect 6411 9024 6423 9027
rect 6457 9027 6515 9033
rect 6457 9024 6469 9027
rect 6411 8996 6469 9024
rect 6411 8993 6423 8996
rect 6365 8987 6423 8993
rect 6457 8993 6469 8996
rect 6503 9024 6515 9027
rect 6822 9024 6828 9036
rect 6503 8996 6828 9024
rect 6503 8993 6515 8996
rect 6457 8987 6515 8993
rect 6822 8984 6828 8996
rect 6880 9024 6886 9036
rect 6880 8996 8892 9024
rect 6880 8984 6886 8996
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 3016 8928 3372 8956
rect 3016 8916 3022 8928
rect 3053 8891 3111 8897
rect 3053 8888 3065 8891
rect 2332 8860 3065 8888
rect 3053 8857 3065 8860
rect 3099 8857 3111 8891
rect 3053 8851 3111 8857
rect 3237 8891 3295 8897
rect 3237 8857 3249 8891
rect 3283 8857 3295 8891
rect 3344 8888 3372 8928
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 4338 8956 4344 8968
rect 3660 8928 4344 8956
rect 3660 8916 3666 8928
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 4982 8956 4988 8968
rect 4448 8928 4988 8956
rect 3789 8891 3847 8897
rect 3789 8888 3801 8891
rect 3344 8860 3801 8888
rect 3237 8851 3295 8857
rect 3789 8857 3801 8860
rect 3835 8857 3847 8891
rect 3789 8851 3847 8857
rect 3973 8891 4031 8897
rect 3973 8857 3985 8891
rect 4019 8857 4031 8891
rect 4154 8888 4160 8900
rect 4115 8860 4160 8888
rect 3973 8851 4031 8857
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 2593 8823 2651 8829
rect 2593 8820 2605 8823
rect 2372 8792 2605 8820
rect 2372 8780 2378 8792
rect 2593 8789 2605 8792
rect 2639 8820 2651 8823
rect 2774 8820 2780 8832
rect 2639 8792 2780 8820
rect 2639 8789 2651 8792
rect 2593 8783 2651 8789
rect 2774 8780 2780 8792
rect 2832 8820 2838 8832
rect 2961 8823 3019 8829
rect 2961 8820 2973 8823
rect 2832 8792 2973 8820
rect 2832 8780 2838 8792
rect 2961 8789 2973 8792
rect 3007 8820 3019 8823
rect 3252 8820 3280 8851
rect 3697 8823 3755 8829
rect 3697 8820 3709 8823
rect 3007 8792 3709 8820
rect 3007 8789 3019 8792
rect 2961 8783 3019 8789
rect 3697 8789 3709 8792
rect 3743 8820 3755 8823
rect 3988 8820 4016 8851
rect 4154 8848 4160 8860
rect 4212 8848 4218 8900
rect 4249 8891 4307 8897
rect 4249 8857 4261 8891
rect 4295 8888 4307 8891
rect 4448 8888 4476 8928
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 8864 8965 8892 8996
rect 8849 8959 8907 8965
rect 8849 8925 8861 8959
rect 8895 8925 8907 8959
rect 8849 8919 8907 8925
rect 4295 8860 4476 8888
rect 6089 8891 6147 8897
rect 4295 8857 4307 8860
rect 4249 8851 4307 8857
rect 6089 8857 6101 8891
rect 6135 8857 6147 8891
rect 6089 8851 6147 8857
rect 6733 8891 6791 8897
rect 6733 8857 6745 8891
rect 6779 8888 6791 8891
rect 7006 8888 7012 8900
rect 6779 8860 7012 8888
rect 6779 8857 6791 8860
rect 6733 8851 6791 8857
rect 4264 8820 4292 8851
rect 3743 8792 4292 8820
rect 6104 8820 6132 8851
rect 7006 8848 7012 8860
rect 7064 8848 7070 8900
rect 8110 8888 8116 8900
rect 7958 8860 8116 8888
rect 8110 8848 8116 8860
rect 8168 8888 8174 8900
rect 8662 8888 8668 8900
rect 8168 8860 8668 8888
rect 8168 8848 8174 8860
rect 8662 8848 8668 8860
rect 8720 8848 8726 8900
rect 8956 8820 8984 9064
rect 16546 9024 16574 9064
rect 16758 9024 16764 9036
rect 16546 8996 16764 9024
rect 16758 8984 16764 8996
rect 16816 8984 16822 9036
rect 9048 8860 16574 8888
rect 9048 8829 9076 8860
rect 16546 8832 16574 8860
rect 6104 8792 8984 8820
rect 9033 8823 9091 8829
rect 3743 8789 3755 8792
rect 3697 8783 3755 8789
rect 9033 8789 9045 8823
rect 9079 8789 9091 8823
rect 9306 8820 9312 8832
rect 9267 8792 9312 8820
rect 9033 8783 9091 8789
rect 9306 8780 9312 8792
rect 9364 8780 9370 8832
rect 16546 8792 16580 8832
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 920 8730 9844 8752
rect 920 8678 3816 8730
rect 3868 8678 3880 8730
rect 3932 8678 3944 8730
rect 3996 8678 4008 8730
rect 4060 8678 4072 8730
rect 4124 8678 8816 8730
rect 8868 8678 8880 8730
rect 8932 8678 8944 8730
rect 8996 8678 9008 8730
rect 9060 8678 9072 8730
rect 9124 8678 9844 8730
rect 920 8656 9844 8678
rect 4522 8576 4528 8628
rect 4580 8616 4586 8628
rect 5626 8616 5632 8628
rect 4580 8588 5632 8616
rect 4580 8576 4586 8588
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 8018 8616 8024 8628
rect 6052 8588 6914 8616
rect 7979 8588 8024 8616
rect 6052 8576 6058 8588
rect 1762 8548 1768 8560
rect 1723 8520 1768 8548
rect 1762 8508 1768 8520
rect 1820 8508 1826 8560
rect 2774 8508 2780 8560
rect 2832 8508 2838 8560
rect 4706 8508 4712 8560
rect 4764 8548 4770 8560
rect 6181 8551 6239 8557
rect 6181 8548 6193 8551
rect 4764 8520 6193 8548
rect 4764 8508 4770 8520
rect 6181 8517 6193 8520
rect 6227 8517 6239 8551
rect 6886 8548 6914 8588
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8386 8548 8392 8560
rect 6886 8520 8392 8548
rect 6181 8511 6239 8517
rect 8386 8508 8392 8520
rect 8444 8508 8450 8560
rect 8662 8508 8668 8560
rect 8720 8548 8726 8560
rect 8941 8551 8999 8557
rect 8941 8548 8953 8551
rect 8720 8520 8953 8548
rect 8720 8508 8726 8520
rect 8941 8517 8953 8520
rect 8987 8548 8999 8551
rect 8987 8520 9260 8548
rect 8987 8517 8999 8520
rect 8941 8511 8999 8517
rect 9232 8492 9260 8520
rect 4614 8440 4620 8492
rect 4672 8480 4678 8492
rect 5810 8480 5816 8492
rect 4672 8452 5816 8480
rect 4672 8440 4678 8452
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 5994 8480 6000 8492
rect 5955 8452 6000 8480
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 8573 8483 8631 8489
rect 8573 8480 8585 8483
rect 8260 8452 8585 8480
rect 8260 8440 8266 8452
rect 8573 8449 8585 8452
rect 8619 8449 8631 8483
rect 8573 8443 8631 8449
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 1486 8412 1492 8424
rect 1447 8384 1492 8412
rect 1486 8372 1492 8384
rect 1544 8372 1550 8424
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8412 3295 8415
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 3283 8384 3985 8412
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 3973 8381 3985 8384
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 5074 8372 5080 8424
rect 5132 8412 5138 8424
rect 9140 8412 9168 8443
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 9272 8452 9317 8480
rect 9272 8440 9278 8452
rect 9306 8412 9312 8424
rect 5132 8384 9312 8412
rect 5132 8372 5138 8384
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 4709 8347 4767 8353
rect 4709 8313 4721 8347
rect 4755 8344 4767 8347
rect 4798 8344 4804 8356
rect 4755 8316 4804 8344
rect 4755 8313 4767 8316
rect 4709 8307 4767 8313
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 6086 8304 6092 8356
rect 6144 8344 6150 8356
rect 6822 8344 6828 8356
rect 6144 8316 6828 8344
rect 6144 8304 6150 8316
rect 6822 8304 6828 8316
rect 6880 8344 6886 8356
rect 7469 8347 7527 8353
rect 7469 8344 7481 8347
rect 6880 8316 7481 8344
rect 6880 8304 6886 8316
rect 7469 8313 7481 8316
rect 7515 8313 7527 8347
rect 7469 8307 7527 8313
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 8757 8347 8815 8353
rect 8757 8344 8769 8347
rect 8352 8316 8769 8344
rect 8352 8304 8358 8316
rect 8757 8313 8769 8316
rect 8803 8313 8815 8347
rect 8757 8307 8815 8313
rect 9401 8347 9459 8353
rect 9401 8313 9413 8347
rect 9447 8344 9459 8347
rect 16574 8344 16580 8356
rect 9447 8316 16580 8344
rect 9447 8313 9459 8316
rect 9401 8307 9459 8313
rect 16574 8304 16580 8316
rect 16632 8304 16638 8356
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 3421 8279 3479 8285
rect 3421 8276 3433 8279
rect 3200 8248 3433 8276
rect 3200 8236 3206 8248
rect 3421 8245 3433 8248
rect 3467 8245 3479 8279
rect 3421 8239 3479 8245
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 7566 8186
rect 7618 8134 7630 8186
rect 7682 8134 7694 8186
rect 7746 8134 7758 8186
rect 7810 8134 7822 8186
rect 7874 8134 9844 8186
rect 920 8112 9844 8134
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 2958 8072 2964 8084
rect 2823 8044 2964 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 2958 8032 2964 8044
rect 3016 8072 3022 8084
rect 3602 8072 3608 8084
rect 3016 8044 3608 8072
rect 3016 8032 3022 8044
rect 3602 8032 3608 8044
rect 3660 8032 3666 8084
rect 4706 8072 4712 8084
rect 4667 8044 4712 8072
rect 4706 8032 4712 8044
rect 4764 8072 4770 8084
rect 5074 8072 5080 8084
rect 4764 8044 5080 8072
rect 4764 8032 4770 8044
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 9306 8032 9312 8084
rect 9364 8072 9370 8084
rect 9401 8075 9459 8081
rect 9401 8072 9413 8075
rect 9364 8044 9413 8072
rect 9364 8032 9370 8044
rect 9401 8041 9413 8044
rect 9447 8041 9459 8075
rect 9401 8035 9459 8041
rect 3694 8004 3700 8016
rect 3655 7976 3700 8004
rect 3694 7964 3700 7976
rect 3752 7964 3758 8016
rect 9033 8007 9091 8013
rect 9033 7973 9045 8007
rect 9079 8004 9091 8007
rect 9490 8004 9496 8016
rect 9079 7976 9496 8004
rect 9079 7973 9091 7976
rect 9033 7967 9091 7973
rect 9490 7964 9496 7976
rect 9548 7964 9554 8016
rect 4798 7936 4804 7948
rect 3068 7908 4804 7936
rect 3068 7877 3096 7908
rect 4798 7896 4804 7908
rect 4856 7896 4862 7948
rect 5902 7896 5908 7948
rect 5960 7936 5966 7948
rect 6089 7939 6147 7945
rect 6089 7936 6101 7939
rect 5960 7908 6101 7936
rect 5960 7896 5966 7908
rect 6089 7905 6101 7908
rect 6135 7905 6147 7939
rect 6089 7899 6147 7905
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 9309 7939 9367 7945
rect 9309 7936 9321 7939
rect 8628 7908 9321 7936
rect 8628 7896 8634 7908
rect 9309 7905 9321 7908
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7837 3111 7871
rect 3602 7868 3608 7880
rect 3563 7840 3608 7868
rect 3053 7831 3111 7837
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 3712 7840 4077 7868
rect 3237 7803 3295 7809
rect 3237 7769 3249 7803
rect 3283 7800 3295 7803
rect 3712 7800 3740 7840
rect 4065 7837 4077 7840
rect 4111 7868 4123 7871
rect 4522 7868 4528 7880
rect 4111 7840 4528 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4522 7828 4528 7840
rect 4580 7868 4586 7880
rect 4982 7868 4988 7880
rect 4580 7840 4988 7868
rect 4580 7828 4586 7840
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 6454 7868 6460 7880
rect 6415 7840 6460 7868
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8294 7868 8300 7880
rect 7975 7840 8300 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 8404 7840 16574 7868
rect 3283 7772 3740 7800
rect 5997 7803 6055 7809
rect 3283 7769 3295 7772
rect 3237 7763 3295 7769
rect 5997 7769 6009 7803
rect 6043 7769 6055 7803
rect 8110 7800 8116 7812
rect 7590 7772 8116 7800
rect 5997 7763 6055 7769
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 2961 7735 3019 7741
rect 2961 7732 2973 7735
rect 2832 7704 2973 7732
rect 2832 7692 2838 7704
rect 2961 7701 2973 7704
rect 3007 7701 3019 7735
rect 2961 7695 3019 7701
rect 3421 7735 3479 7741
rect 3421 7701 3433 7735
rect 3467 7732 3479 7735
rect 6012 7732 6040 7763
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 8404 7732 8432 7840
rect 8493 7803 8551 7809
rect 8493 7769 8505 7803
rect 8539 7800 8551 7803
rect 16546 7800 16574 7840
rect 16666 7800 16672 7812
rect 8539 7772 12572 7800
rect 16546 7772 16672 7800
rect 8539 7769 8551 7772
rect 8493 7763 8551 7769
rect 3467 7704 8432 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 8849 7735 8907 7741
rect 8849 7732 8861 7735
rect 8720 7704 8861 7732
rect 8720 7692 8726 7704
rect 8849 7701 8861 7704
rect 8895 7701 8907 7735
rect 12544 7732 12572 7772
rect 16666 7760 16672 7772
rect 16724 7760 16730 7812
rect 16574 7732 16580 7744
rect 12544 7704 16580 7732
rect 8849 7695 8907 7701
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 920 7642 9844 7664
rect 920 7590 3816 7642
rect 3868 7590 3880 7642
rect 3932 7590 3944 7642
rect 3996 7590 4008 7642
rect 4060 7590 4072 7642
rect 4124 7590 8816 7642
rect 8868 7590 8880 7642
rect 8932 7590 8944 7642
rect 8996 7590 9008 7642
rect 9060 7590 9072 7642
rect 9124 7590 9844 7642
rect 920 7568 9844 7590
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 3050 7528 3056 7540
rect 2547 7500 3056 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 9214 7488 9220 7540
rect 9272 7528 9278 7540
rect 9401 7531 9459 7537
rect 9401 7528 9413 7531
rect 9272 7500 9413 7528
rect 9272 7488 9278 7500
rect 9401 7497 9413 7500
rect 9447 7497 9459 7531
rect 9401 7491 9459 7497
rect 3694 7420 3700 7472
rect 3752 7420 3758 7472
rect 5994 7420 6000 7472
rect 6052 7460 6058 7472
rect 6178 7460 6184 7472
rect 6052 7432 6184 7460
rect 6052 7420 6058 7432
rect 6178 7420 6184 7432
rect 6236 7420 6242 7472
rect 7926 7460 7932 7472
rect 7887 7432 7932 7460
rect 7926 7420 7932 7432
rect 7984 7420 7990 7472
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 9033 7463 9091 7469
rect 9033 7460 9045 7463
rect 8168 7432 9045 7460
rect 8168 7420 8174 7432
rect 9033 7429 9045 7432
rect 9079 7429 9091 7463
rect 9033 7423 9091 7429
rect 2774 7392 2780 7404
rect 2735 7364 2780 7392
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 3142 7392 3148 7404
rect 3103 7364 3148 7392
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 4212 7364 4629 7392
rect 4212 7352 4218 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 4982 7352 4988 7404
rect 5040 7392 5046 7404
rect 9232 7401 9260 7488
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 5040 7364 5549 7392
rect 5040 7352 5046 7364
rect 5537 7361 5549 7364
rect 5583 7392 5595 7395
rect 9217 7395 9275 7401
rect 9217 7392 9229 7395
rect 5583 7364 9229 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 9217 7361 9229 7364
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 5810 7324 5816 7336
rect 4908 7296 5816 7324
rect 2685 7191 2743 7197
rect 2685 7157 2697 7191
rect 2731 7188 2743 7191
rect 4908 7188 4936 7296
rect 5810 7284 5816 7296
rect 5868 7324 5874 7336
rect 6546 7324 6552 7336
rect 5868 7296 6552 7324
rect 5868 7284 5874 7296
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 8352 7296 8585 7324
rect 8352 7284 8358 7296
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 8573 7287 8631 7293
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7324 8999 7327
rect 9306 7324 9312 7336
rect 8987 7296 9312 7324
rect 8987 7293 8999 7296
rect 8941 7287 8999 7293
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 5181 7259 5239 7265
rect 5181 7225 5193 7259
rect 5227 7256 5239 7259
rect 6822 7256 6828 7268
rect 5227 7228 6828 7256
rect 5227 7225 5239 7228
rect 5181 7219 5239 7225
rect 6822 7216 6828 7228
rect 6880 7216 6886 7268
rect 5902 7188 5908 7200
rect 2731 7160 4936 7188
rect 5863 7160 5908 7188
rect 2731 7157 2743 7160
rect 2685 7151 2743 7157
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 6512 7160 8033 7188
rect 6512 7148 6518 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 8570 7148 8576 7200
rect 8628 7188 8634 7200
rect 8846 7188 8852 7200
rect 8628 7160 8852 7188
rect 8628 7148 8634 7160
rect 8846 7148 8852 7160
rect 8904 7148 8910 7200
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 7566 7098
rect 7618 7046 7630 7098
rect 7682 7046 7694 7098
rect 7746 7046 7758 7098
rect 7810 7046 7822 7098
rect 7874 7046 9844 7098
rect 920 7024 9844 7046
rect 1752 6987 1810 6993
rect 1752 6953 1764 6987
rect 1798 6984 1810 6987
rect 3142 6984 3148 6996
rect 1798 6956 3148 6984
rect 1798 6953 1810 6956
rect 1752 6947 1810 6953
rect 3142 6944 3148 6956
rect 3200 6944 3206 6996
rect 4798 6944 4804 6996
rect 4856 6984 4862 6996
rect 4856 6956 6960 6984
rect 4856 6944 4862 6956
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 4157 6851 4215 6857
rect 4157 6848 4169 6851
rect 3283 6820 4169 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 4157 6817 4169 6820
rect 4203 6817 4215 6851
rect 6932 6848 6960 6956
rect 7466 6944 7472 6996
rect 7524 6993 7530 6996
rect 7524 6984 7535 6993
rect 7524 6956 7569 6984
rect 7524 6947 7535 6956
rect 7524 6944 7530 6947
rect 8846 6876 8852 6928
rect 8904 6876 8910 6928
rect 9493 6919 9551 6925
rect 9493 6885 9505 6919
rect 9539 6885 9551 6919
rect 9493 6879 9551 6885
rect 8864 6848 8892 6876
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 6932 6820 7880 6848
rect 8864 6820 8953 6848
rect 4157 6811 4215 6817
rect 1486 6780 1492 6792
rect 1447 6752 1492 6780
rect 1486 6740 1492 6752
rect 1544 6740 1550 6792
rect 3050 6740 3056 6792
rect 3108 6780 3114 6792
rect 3694 6780 3700 6792
rect 3108 6752 3700 6780
rect 3108 6740 3114 6752
rect 3694 6740 3700 6752
rect 3752 6780 3758 6792
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 3752 6752 4353 6780
rect 3752 6740 3758 6752
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 4522 6740 4528 6792
rect 4580 6780 4586 6792
rect 4801 6783 4859 6789
rect 4801 6780 4813 6783
rect 4580 6752 4813 6780
rect 4580 6740 4586 6752
rect 4801 6749 4813 6752
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6749 5135 6783
rect 5442 6780 5448 6792
rect 5403 6752 5448 6780
rect 5077 6743 5135 6749
rect 2406 6672 2412 6724
rect 2464 6672 2470 6724
rect 4246 6672 4252 6724
rect 4304 6712 4310 6724
rect 4617 6715 4675 6721
rect 4617 6712 4629 6715
rect 4304 6684 4629 6712
rect 4304 6672 4310 6684
rect 4617 6681 4629 6684
rect 4663 6681 4675 6715
rect 4617 6675 4675 6681
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 3605 6647 3663 6653
rect 3605 6644 3617 6647
rect 3200 6616 3617 6644
rect 3200 6604 3206 6616
rect 3605 6613 3617 6616
rect 3651 6613 3663 6647
rect 5092 6644 5120 6743
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6780 6975 6783
rect 7466 6780 7472 6792
rect 6963 6752 7472 6780
rect 6963 6749 6975 6752
rect 6917 6743 6975 6749
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7852 6789 7880 6820
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8570 6780 8576 6792
rect 8531 6752 8576 6780
rect 8113 6743 8171 6749
rect 5902 6672 5908 6724
rect 5960 6672 5966 6724
rect 7745 6715 7803 6721
rect 7745 6712 7757 6715
rect 6656 6684 7757 6712
rect 6656 6644 6684 6684
rect 7745 6681 7757 6684
rect 7791 6681 7803 6715
rect 7745 6675 7803 6681
rect 5092 6616 6684 6644
rect 3605 6607 3663 6613
rect 6822 6604 6828 6656
rect 6880 6644 6886 6656
rect 8128 6644 8156 6743
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 8956 6780 8984 6811
rect 9214 6780 9220 6792
rect 8956 6752 9220 6780
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9508 6780 9536 6879
rect 16574 6780 16580 6792
rect 9508 6752 16580 6780
rect 16574 6740 16580 6752
rect 16632 6740 16638 6792
rect 8297 6715 8355 6721
rect 8297 6681 8309 6715
rect 8343 6712 8355 6715
rect 8386 6712 8392 6724
rect 8343 6684 8392 6712
rect 8343 6681 8355 6684
rect 8297 6675 8355 6681
rect 8386 6672 8392 6684
rect 8444 6672 8450 6724
rect 9033 6715 9091 6721
rect 9033 6681 9045 6715
rect 9079 6712 9091 6715
rect 9306 6712 9312 6724
rect 9079 6684 9312 6712
rect 9079 6681 9091 6684
rect 9033 6675 9091 6681
rect 9306 6672 9312 6684
rect 9364 6672 9370 6724
rect 6880 6616 8156 6644
rect 9125 6647 9183 6653
rect 6880 6604 6886 6616
rect 9125 6613 9137 6647
rect 9171 6644 9183 6647
rect 9398 6644 9404 6656
rect 9171 6616 9404 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 920 6554 9844 6576
rect 920 6502 3816 6554
rect 3868 6502 3880 6554
rect 3932 6502 3944 6554
rect 3996 6502 4008 6554
rect 4060 6502 4072 6554
rect 4124 6502 8816 6554
rect 8868 6502 8880 6554
rect 8932 6502 8944 6554
rect 8996 6502 9008 6554
rect 9060 6502 9072 6554
rect 9124 6502 9844 6554
rect 920 6480 9844 6502
rect 13814 6468 13820 6520
rect 13872 6508 13878 6520
rect 16666 6508 16672 6520
rect 13872 6480 16672 6508
rect 13872 6468 13878 6480
rect 16666 6468 16672 6480
rect 16724 6468 16730 6520
rect 2225 6443 2283 6449
rect 2225 6409 2237 6443
rect 2271 6440 2283 6443
rect 3050 6440 3056 6452
rect 2271 6412 3056 6440
rect 2271 6409 2283 6412
rect 2225 6403 2283 6409
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 7524 6412 7788 6440
rect 7524 6400 7530 6412
rect 4252 6384 4304 6390
rect 2041 6375 2099 6381
rect 2041 6341 2053 6375
rect 2087 6372 2099 6375
rect 2406 6372 2412 6384
rect 2087 6344 2412 6372
rect 2087 6341 2099 6344
rect 2041 6335 2099 6341
rect 2406 6332 2412 6344
rect 2464 6332 2470 6384
rect 5353 6375 5411 6381
rect 5353 6341 5365 6375
rect 5399 6372 5411 6375
rect 5442 6372 5448 6384
rect 5399 6344 5448 6372
rect 5399 6341 5411 6344
rect 5353 6335 5411 6341
rect 5442 6332 5448 6344
rect 5500 6372 5506 6384
rect 6457 6375 6515 6381
rect 6457 6372 6469 6375
rect 5500 6344 6469 6372
rect 5500 6332 5506 6344
rect 6457 6341 6469 6344
rect 6503 6341 6515 6375
rect 7760 6372 7788 6412
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 7984 6412 8125 6440
rect 7984 6400 7990 6412
rect 8113 6409 8125 6412
rect 8159 6409 8171 6443
rect 8113 6403 8171 6409
rect 8662 6400 8668 6452
rect 8720 6400 8726 6452
rect 8846 6400 8852 6452
rect 8904 6440 8910 6452
rect 8941 6443 8999 6449
rect 8941 6440 8953 6443
rect 8904 6412 8953 6440
rect 8904 6400 8910 6412
rect 8941 6409 8953 6412
rect 8987 6409 8999 6443
rect 8941 6403 8999 6409
rect 9033 6443 9091 6449
rect 9033 6409 9045 6443
rect 9079 6409 9091 6443
rect 9033 6403 9091 6409
rect 8297 6375 8355 6381
rect 8297 6372 8309 6375
rect 7760 6344 8309 6372
rect 6457 6335 6515 6341
rect 8297 6341 8309 6344
rect 8343 6341 8355 6375
rect 8680 6372 8708 6400
rect 8757 6375 8815 6381
rect 8757 6372 8769 6375
rect 8680 6344 8769 6372
rect 8297 6335 8355 6341
rect 8757 6341 8769 6344
rect 8803 6341 8815 6375
rect 9048 6372 9076 6403
rect 8757 6335 8815 6341
rect 8956 6344 9076 6372
rect 9125 6375 9183 6381
rect 4252 6326 4304 6332
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 4614 6304 4620 6316
rect 2731 6276 2912 6304
rect 4575 6276 4620 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 2593 6239 2651 6245
rect 2593 6205 2605 6239
rect 2639 6236 2651 6239
rect 2777 6239 2835 6245
rect 2777 6236 2789 6239
rect 2639 6208 2789 6236
rect 2639 6205 2651 6208
rect 2593 6199 2651 6205
rect 2777 6205 2789 6208
rect 2823 6205 2835 6239
rect 2777 6199 2835 6205
rect 2884 6100 2912 6276
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 6181 6307 6239 6313
rect 6181 6304 6193 6307
rect 6052 6276 6193 6304
rect 6052 6264 6058 6276
rect 6181 6273 6193 6276
rect 6227 6273 6239 6307
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 7590 6276 8493 6304
rect 6181 6267 6239 6273
rect 8481 6273 8493 6276
rect 8527 6304 8539 6307
rect 8665 6307 8723 6313
rect 8527 6276 8616 6304
rect 8527 6273 8539 6276
rect 8481 6267 8539 6273
rect 8588 6248 8616 6276
rect 8665 6273 8677 6307
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 3142 6236 3148 6248
rect 3103 6208 3148 6236
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 5902 6236 5908 6248
rect 5863 6208 5908 6236
rect 5902 6196 5908 6208
rect 5960 6196 5966 6248
rect 6546 6196 6552 6248
rect 6604 6236 6610 6248
rect 7929 6239 7987 6245
rect 6604 6208 7880 6236
rect 6604 6196 6610 6208
rect 7852 6168 7880 6208
rect 7929 6205 7941 6239
rect 7975 6236 7987 6239
rect 8294 6236 8300 6248
rect 7975 6208 8300 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 8570 6196 8576 6248
rect 8628 6196 8634 6248
rect 8478 6168 8484 6180
rect 7852 6140 8484 6168
rect 8478 6128 8484 6140
rect 8536 6168 8542 6180
rect 8680 6168 8708 6267
rect 8536 6140 8708 6168
rect 8536 6128 8542 6140
rect 4982 6100 4988 6112
rect 2884 6072 4988 6100
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5181 6103 5239 6109
rect 5181 6069 5193 6103
rect 5227 6100 5239 6103
rect 5442 6100 5448 6112
rect 5227 6072 5448 6100
rect 5227 6069 5239 6072
rect 5181 6063 5239 6069
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 8956 6100 8984 6344
rect 9125 6341 9137 6375
rect 9171 6372 9183 6375
rect 9214 6372 9220 6384
rect 9171 6344 9220 6372
rect 9171 6341 9183 6344
rect 9125 6335 9183 6341
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 9309 6171 9367 6177
rect 9309 6137 9321 6171
rect 9355 6168 9367 6171
rect 19426 6168 19432 6180
rect 9355 6140 19432 6168
rect 9355 6137 9367 6140
rect 9309 6131 9367 6137
rect 19426 6128 19432 6140
rect 19484 6128 19490 6180
rect 8628 6072 8984 6100
rect 8628 6060 8634 6072
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9401 6103 9459 6109
rect 9401 6100 9413 6103
rect 9272 6072 9413 6100
rect 9272 6060 9278 6072
rect 9401 6069 9413 6072
rect 9447 6069 9459 6103
rect 9401 6063 9459 6069
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 7566 6010
rect 7618 5958 7630 6010
rect 7682 5958 7694 6010
rect 7746 5958 7758 6010
rect 7810 5958 7822 6010
rect 7874 5958 9844 6010
rect 920 5936 9844 5958
rect 1844 5899 1902 5905
rect 1844 5865 1856 5899
rect 1890 5896 1902 5899
rect 3142 5896 3148 5908
rect 1890 5868 3148 5896
rect 1890 5865 1902 5868
rect 1844 5859 1902 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3973 5899 4031 5905
rect 3973 5865 3985 5899
rect 4019 5896 4031 5899
rect 4614 5896 4620 5908
rect 4019 5868 4620 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5902 5896 5908 5908
rect 5863 5868 5908 5896
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 6880 5868 8432 5896
rect 6880 5856 6886 5868
rect 8404 5837 8432 5868
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 8536 5868 8581 5896
rect 8536 5856 8542 5868
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 9214 5896 9220 5908
rect 8720 5868 9220 5896
rect 8720 5856 8726 5868
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 8389 5831 8447 5837
rect 8389 5797 8401 5831
rect 8435 5828 8447 5831
rect 8435 5800 16574 5828
rect 8435 5797 8447 5800
rect 8389 5791 8447 5797
rect 1486 5720 1492 5772
rect 1544 5760 1550 5772
rect 1581 5763 1639 5769
rect 1581 5760 1593 5763
rect 1544 5732 1593 5760
rect 1544 5720 1550 5732
rect 1581 5729 1593 5732
rect 1627 5760 1639 5763
rect 4433 5763 4491 5769
rect 1627 5732 3372 5760
rect 1627 5729 1639 5732
rect 1581 5723 1639 5729
rect 3344 5704 3372 5732
rect 4433 5729 4445 5763
rect 4479 5760 4491 5763
rect 5718 5760 5724 5772
rect 4479 5732 5724 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 5994 5720 6000 5772
rect 6052 5760 6058 5772
rect 6181 5763 6239 5769
rect 6181 5760 6193 5763
rect 6052 5732 6193 5760
rect 6052 5720 6058 5732
rect 6181 5729 6193 5732
rect 6227 5729 6239 5763
rect 6454 5760 6460 5772
rect 6415 5732 6460 5760
rect 6181 5723 6239 5729
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 7929 5763 7987 5769
rect 7929 5729 7941 5763
rect 7975 5760 7987 5763
rect 8662 5760 8668 5772
rect 7975 5732 8668 5760
rect 7975 5729 7987 5732
rect 7929 5723 7987 5729
rect 8662 5720 8668 5732
rect 8720 5720 8726 5772
rect 8846 5760 8852 5772
rect 8807 5732 8852 5760
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 3326 5652 3332 5704
rect 3384 5692 3390 5704
rect 4157 5695 4215 5701
rect 4157 5692 4169 5695
rect 3384 5664 4169 5692
rect 3384 5652 3390 5664
rect 4157 5661 4169 5664
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 1489 5627 1547 5633
rect 1489 5593 1501 5627
rect 1535 5624 1547 5627
rect 2314 5624 2320 5636
rect 1535 5596 2320 5624
rect 1535 5593 1547 5596
rect 1489 5587 1547 5593
rect 2240 5556 2268 5596
rect 2314 5584 2320 5596
rect 2372 5584 2378 5636
rect 3697 5627 3755 5633
rect 3252 5596 3648 5624
rect 3252 5556 3280 5596
rect 2240 5528 3280 5556
rect 3329 5559 3387 5565
rect 3329 5525 3341 5559
rect 3375 5556 3387 5559
rect 3510 5556 3516 5568
rect 3375 5528 3516 5556
rect 3375 5525 3387 5528
rect 3329 5519 3387 5525
rect 3510 5516 3516 5528
rect 3568 5516 3574 5568
rect 3620 5556 3648 5596
rect 3697 5593 3709 5627
rect 3743 5624 3755 5627
rect 3786 5624 3792 5636
rect 3743 5596 3792 5624
rect 3743 5593 3755 5596
rect 3697 5587 3755 5593
rect 3786 5584 3792 5596
rect 3844 5584 3850 5636
rect 3881 5627 3939 5633
rect 3881 5593 3893 5627
rect 3927 5593 3939 5627
rect 3881 5587 3939 5593
rect 4540 5596 4922 5624
rect 7682 5596 8248 5624
rect 3896 5556 3924 5587
rect 4540 5568 4568 5596
rect 4154 5556 4160 5568
rect 3620 5528 4160 5556
rect 4154 5516 4160 5528
rect 4212 5556 4218 5568
rect 4522 5556 4528 5568
rect 4212 5528 4528 5556
rect 4212 5516 4218 5528
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 4816 5556 4844 5596
rect 7760 5556 7788 5596
rect 8220 5565 8248 5596
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 8941 5627 8999 5633
rect 8444 5596 8616 5624
rect 8444 5584 8450 5596
rect 4816 5528 7788 5556
rect 8205 5559 8263 5565
rect 8205 5525 8217 5559
rect 8251 5556 8263 5559
rect 8478 5556 8484 5568
rect 8251 5528 8484 5556
rect 8251 5525 8263 5528
rect 8205 5519 8263 5525
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 8588 5556 8616 5596
rect 8941 5593 8953 5627
rect 8987 5593 8999 5627
rect 9490 5624 9496 5636
rect 9451 5596 9496 5624
rect 8941 5587 8999 5593
rect 8956 5556 8984 5587
rect 9490 5584 9496 5596
rect 9548 5584 9554 5636
rect 8588 5528 8984 5556
rect 16546 5568 16574 5800
rect 16546 5528 16580 5568
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 920 5466 9844 5488
rect 920 5414 3816 5466
rect 3868 5414 3880 5466
rect 3932 5414 3944 5466
rect 3996 5414 4008 5466
rect 4060 5414 4072 5466
rect 4124 5414 8816 5466
rect 8868 5414 8880 5466
rect 8932 5414 8944 5466
rect 8996 5414 9008 5466
rect 9060 5414 9072 5466
rect 9124 5414 9844 5466
rect 920 5392 9844 5414
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 7064 5324 8309 5352
rect 7064 5312 7070 5324
rect 8297 5321 8309 5324
rect 8343 5321 8355 5355
rect 8297 5315 8355 5321
rect 4154 5244 4160 5296
rect 4212 5244 4218 5296
rect 8113 5287 8171 5293
rect 8113 5284 8125 5287
rect 7498 5256 8125 5284
rect 8113 5253 8125 5256
rect 8159 5284 8171 5287
rect 8478 5284 8484 5296
rect 8159 5256 8484 5284
rect 8159 5253 8171 5256
rect 8113 5247 8171 5253
rect 8478 5244 8484 5256
rect 8536 5284 8542 5296
rect 8536 5256 9260 5284
rect 8536 5244 8542 5256
rect 9232 5228 9260 5256
rect 5994 5216 6000 5228
rect 5955 5188 6000 5216
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 8352 5188 9045 5216
rect 8352 5176 8358 5188
rect 9033 5185 9045 5188
rect 9079 5185 9091 5219
rect 9214 5216 9220 5228
rect 9175 5188 9220 5216
rect 9033 5179 9091 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 3326 5148 3332 5160
rect 3287 5120 3332 5148
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 3602 5148 3608 5160
rect 3515 5120 3608 5148
rect 3602 5108 3608 5120
rect 3660 5148 3666 5160
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 3660 5120 5273 5148
rect 3660 5108 3666 5120
rect 5261 5117 5273 5120
rect 5307 5117 5319 5151
rect 5810 5148 5816 5160
rect 5771 5120 5816 5148
rect 5261 5111 5319 5117
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 6273 5151 6331 5157
rect 6273 5117 6285 5151
rect 6319 5148 6331 5151
rect 6914 5148 6920 5160
rect 6319 5120 6920 5148
rect 6319 5117 6331 5120
rect 6273 5111 6331 5117
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7745 5151 7803 5157
rect 7745 5117 7757 5151
rect 7791 5148 7803 5151
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 7791 5120 8861 5148
rect 7791 5117 7803 5120
rect 7745 5111 7803 5117
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5166 5012 5172 5024
rect 5123 4984 5172 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 8386 4972 8392 5024
rect 8444 5012 8450 5024
rect 9309 5015 9367 5021
rect 9309 5012 9321 5015
rect 8444 4984 9321 5012
rect 8444 4972 8450 4984
rect 9309 4981 9321 4984
rect 9355 4981 9367 5015
rect 9309 4975 9367 4981
rect 3036 4922 9844 4944
rect 3036 4870 7566 4922
rect 7618 4870 7630 4922
rect 7682 4870 7694 4922
rect 7746 4870 7758 4922
rect 7810 4870 7822 4922
rect 7874 4870 9844 4922
rect 3036 4848 9844 4870
rect 5077 4811 5135 4817
rect 5077 4777 5089 4811
rect 5123 4808 5135 4811
rect 5810 4808 5816 4820
rect 5123 4780 5816 4808
rect 5123 4777 5135 4780
rect 5077 4771 5135 4777
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9272 4780 9413 4808
rect 9272 4768 9278 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 5166 4700 5172 4752
rect 5224 4740 5230 4752
rect 5224 4712 6316 4740
rect 5224 4700 5230 4712
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 5353 4675 5411 4681
rect 5353 4672 5365 4675
rect 4212 4644 5365 4672
rect 4212 4632 4218 4644
rect 5353 4641 5365 4644
rect 5399 4641 5411 4675
rect 5718 4672 5724 4684
rect 5679 4644 5724 4672
rect 5353 4635 5411 4641
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 6288 4681 6316 4712
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4641 6331 4675
rect 6273 4635 6331 4641
rect 9582 4632 9588 4684
rect 9640 4632 9646 4684
rect 3326 4604 3332 4616
rect 3287 4576 3332 4604
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 4982 4564 4988 4616
rect 5040 4604 5046 4616
rect 5442 4604 5448 4616
rect 5040 4576 5448 4604
rect 5040 4564 5046 4576
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 6546 4604 6552 4616
rect 6507 4576 6552 4604
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 7006 4604 7012 4616
rect 6963 4576 7012 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 8386 4604 8392 4616
rect 8347 4576 8392 4604
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 9309 4607 9367 4613
rect 9309 4604 9321 4607
rect 8496 4576 9321 4604
rect 3605 4539 3663 4545
rect 3605 4505 3617 4539
rect 3651 4505 3663 4539
rect 3605 4499 3663 4505
rect 3620 4468 3648 4499
rect 4614 4496 4620 4548
rect 4672 4496 4678 4548
rect 7466 4496 7472 4548
rect 7524 4496 7530 4548
rect 8294 4496 8300 4548
rect 8352 4536 8358 4548
rect 8496 4536 8524 4576
rect 9309 4573 9321 4576
rect 9355 4604 9367 4607
rect 9600 4604 9628 4632
rect 9355 4576 9628 4604
rect 9355 4573 9367 4576
rect 9309 4567 9367 4573
rect 8352 4508 8524 4536
rect 8953 4539 9011 4545
rect 8352 4496 8358 4508
rect 8953 4505 8965 4539
rect 8999 4536 9011 4539
rect 9582 4536 9588 4548
rect 8999 4508 9588 4536
rect 8999 4505 9011 4508
rect 8953 4499 9011 4505
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 4246 4468 4252 4480
rect 3620 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 9214 4468 9220 4480
rect 9175 4440 9220 4468
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 3036 4378 9844 4400
rect 3036 4326 3816 4378
rect 3868 4326 3880 4378
rect 3932 4326 3944 4378
rect 3996 4326 4008 4378
rect 4060 4326 4072 4378
rect 4124 4326 8816 4378
rect 8868 4326 8880 4378
rect 8932 4326 8944 4378
rect 8996 4326 9008 4378
rect 9060 4326 9072 4378
rect 9124 4326 9844 4378
rect 3036 4304 9844 4326
rect 6365 4267 6423 4273
rect 6365 4233 6377 4267
rect 6411 4264 6423 4267
rect 6546 4264 6552 4276
rect 6411 4236 6552 4264
rect 6411 4233 6423 4236
rect 6365 4227 6423 4233
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 5810 4196 5816 4208
rect 5014 4168 5816 4196
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3292 4100 3341 4128
rect 3292 4088 3298 4100
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 5350 4128 5356 4140
rect 3559 4100 4016 4128
rect 5311 4100 5356 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 3602 4020 3608 4072
rect 3660 4060 3666 4072
rect 3881 4063 3939 4069
rect 3881 4060 3893 4063
rect 3660 4032 3893 4060
rect 3660 4020 3666 4032
rect 3881 4029 3893 4032
rect 3927 4029 3939 4063
rect 3988 4060 4016 4100
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 6273 4131 6331 4137
rect 6273 4128 6285 4131
rect 5500 4100 6285 4128
rect 5500 4088 5506 4100
rect 6273 4097 6285 4100
rect 6319 4097 6331 4131
rect 6273 4091 6331 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 9214 4128 9220 4140
rect 8159 4100 9220 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 9398 4128 9404 4140
rect 9359 4100 9404 4128
rect 9398 4088 9404 4100
rect 9456 4088 9462 4140
rect 4154 4060 4160 4072
rect 3988 4032 4160 4060
rect 3881 4023 3939 4029
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 6549 4063 6607 4069
rect 6549 4060 6561 4063
rect 5368 4032 6561 4060
rect 2682 3952 2688 4004
rect 2740 3992 2746 4004
rect 2740 3964 3648 3992
rect 2740 3952 2746 3964
rect 3620 3924 3648 3964
rect 5368 3924 5396 4032
rect 6549 4029 6561 4032
rect 6595 4029 6607 4063
rect 6549 4023 6607 4029
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 8297 4063 8355 4069
rect 8297 4060 8309 4063
rect 6972 4032 8309 4060
rect 6972 4020 6978 4032
rect 8297 4029 8309 4032
rect 8343 4029 8355 4063
rect 8297 4023 8355 4029
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 8720 4032 8861 4060
rect 8720 4020 8726 4032
rect 8849 4029 8861 4032
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 5442 3952 5448 4004
rect 5500 3992 5506 4004
rect 6089 3995 6147 4001
rect 6089 3992 6101 3995
rect 5500 3964 6101 3992
rect 5500 3952 5506 3964
rect 6089 3961 6101 3964
rect 6135 3961 6147 3995
rect 6089 3955 6147 3961
rect 8021 3995 8079 4001
rect 8021 3961 8033 3995
rect 8067 3992 8079 3995
rect 13814 3992 13820 4004
rect 8067 3964 13820 3992
rect 8067 3961 8079 3964
rect 8021 3955 8079 3961
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 5902 3924 5908 3936
rect 5960 3933 5966 3936
rect 3620 3896 5396 3924
rect 5871 3896 5908 3924
rect 5902 3884 5908 3896
rect 5960 3887 5971 3933
rect 5960 3884 5966 3887
rect 8386 3884 8392 3936
rect 8444 3924 8450 3936
rect 9125 3927 9183 3933
rect 9125 3924 9137 3927
rect 8444 3896 9137 3924
rect 8444 3884 8450 3896
rect 9125 3893 9137 3896
rect 9171 3924 9183 3927
rect 9217 3927 9275 3933
rect 9217 3924 9229 3927
rect 9171 3896 9229 3924
rect 9171 3893 9183 3896
rect 9125 3887 9183 3893
rect 9217 3893 9229 3896
rect 9263 3893 9275 3927
rect 9217 3887 9275 3893
rect 3036 3834 9844 3856
rect 3036 3782 7566 3834
rect 7618 3782 7630 3834
rect 7682 3782 7694 3834
rect 7746 3782 7758 3834
rect 7810 3782 7822 3834
rect 7874 3782 9844 3834
rect 3036 3760 9844 3782
rect 5350 3680 5356 3732
rect 5408 3720 5414 3732
rect 5445 3723 5503 3729
rect 5445 3720 5457 3723
rect 5408 3692 5457 3720
rect 5408 3680 5414 3692
rect 5445 3689 5457 3692
rect 5491 3689 5503 3723
rect 5810 3720 5816 3732
rect 5771 3692 5816 3720
rect 5445 3683 5503 3689
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 3421 3587 3479 3593
rect 3421 3584 3433 3587
rect 3384 3556 3433 3584
rect 3384 3544 3390 3556
rect 3421 3553 3433 3556
rect 3467 3553 3479 3587
rect 3421 3547 3479 3553
rect 5626 3544 5632 3596
rect 5684 3584 5690 3596
rect 6546 3584 6552 3596
rect 5684 3556 6552 3584
rect 5684 3544 5690 3556
rect 6546 3544 6552 3556
rect 6604 3584 6610 3596
rect 6604 3556 6776 3584
rect 6604 3544 6610 3556
rect 5074 3516 5080 3528
rect 5035 3488 5080 3516
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 6748 3525 6776 3556
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 7193 3587 7251 3593
rect 7193 3584 7205 3587
rect 6972 3556 7205 3584
rect 6972 3544 6978 3556
rect 7193 3553 7205 3556
rect 7239 3553 7251 3587
rect 7193 3547 7251 3553
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5184 3488 5733 3516
rect 5184 3460 5212 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3516 6239 3519
rect 6733 3519 6791 3525
rect 6227 3488 6592 3516
rect 6227 3485 6239 3488
rect 6181 3479 6239 3485
rect 4338 3408 4344 3460
rect 4396 3448 4402 3460
rect 5166 3448 5172 3460
rect 4396 3420 5172 3448
rect 4396 3408 4402 3420
rect 5166 3408 5172 3420
rect 5224 3408 5230 3460
rect 5353 3451 5411 3457
rect 5353 3417 5365 3451
rect 5399 3448 5411 3451
rect 5442 3448 5448 3460
rect 5399 3420 5448 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 4614 3340 4620 3392
rect 4672 3380 4678 3392
rect 5368 3380 5396 3411
rect 5442 3408 5448 3420
rect 5500 3448 5506 3460
rect 6196 3448 6224 3479
rect 5500 3420 6224 3448
rect 6365 3451 6423 3457
rect 5500 3408 5506 3420
rect 6365 3417 6377 3451
rect 6411 3448 6423 3451
rect 6454 3448 6460 3460
rect 6411 3420 6460 3448
rect 6411 3417 6423 3420
rect 6365 3411 6423 3417
rect 6454 3408 6460 3420
rect 6512 3408 6518 3460
rect 6564 3457 6592 3488
rect 6733 3485 6745 3519
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 7006 3516 7012 3528
rect 6871 3488 7012 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 7006 3476 7012 3488
rect 7064 3476 7070 3528
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8665 3519 8723 3525
rect 8665 3516 8677 3519
rect 8536 3488 8677 3516
rect 8536 3476 8542 3488
rect 8665 3485 8677 3488
rect 8711 3485 8723 3519
rect 8665 3479 8723 3485
rect 6549 3451 6607 3457
rect 6549 3417 6561 3451
rect 6595 3448 6607 3451
rect 6638 3448 6644 3460
rect 6595 3420 6644 3448
rect 6595 3417 6607 3420
rect 6549 3411 6607 3417
rect 6638 3408 6644 3420
rect 6696 3408 6702 3460
rect 7926 3408 7932 3460
rect 7984 3408 7990 3460
rect 8570 3408 8576 3460
rect 8628 3448 8634 3460
rect 9229 3451 9287 3457
rect 8628 3420 8984 3448
rect 8628 3408 8634 3420
rect 4672 3352 5396 3380
rect 4672 3340 4678 3352
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 8849 3383 8907 3389
rect 8849 3380 8861 3383
rect 8720 3352 8861 3380
rect 8720 3340 8726 3352
rect 8849 3349 8861 3352
rect 8895 3349 8907 3383
rect 8956 3380 8984 3420
rect 9229 3417 9241 3451
rect 9275 3448 9287 3451
rect 16574 3448 16580 3460
rect 9275 3420 16580 3448
rect 9275 3417 9287 3420
rect 9229 3411 9287 3417
rect 16574 3408 16580 3420
rect 16632 3408 16638 3460
rect 9398 3380 9404 3392
rect 8956 3352 9404 3380
rect 8849 3343 8907 3349
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 3036 3290 9844 3312
rect 3036 3238 3816 3290
rect 3868 3238 3880 3290
rect 3932 3238 3944 3290
rect 3996 3238 4008 3290
rect 4060 3238 4072 3290
rect 4124 3238 8816 3290
rect 8868 3238 8880 3290
rect 8932 3238 8944 3290
rect 8996 3238 9008 3290
rect 9060 3238 9072 3290
rect 9124 3238 9844 3290
rect 3036 3216 9844 3238
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 4246 3176 4252 3188
rect 4203 3148 4252 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 8386 3176 8392 3188
rect 8159 3148 8392 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 6092 3120 6144 3126
rect 3421 3111 3479 3117
rect 3421 3077 3433 3111
rect 3467 3108 3479 3111
rect 4338 3108 4344 3120
rect 3467 3080 4344 3108
rect 3467 3077 3479 3080
rect 3421 3071 3479 3077
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 7466 3108 7472 3120
rect 7427 3080 7472 3108
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 6092 3062 6144 3068
rect 3510 3040 3516 3052
rect 3471 3012 3516 3040
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 4890 3040 4896 3052
rect 4479 3012 4896 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 6454 3040 6460 3052
rect 6415 3012 6460 3040
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 6696 3012 7297 3040
rect 6696 3000 6702 3012
rect 7285 3009 7297 3012
rect 7331 3040 7343 3043
rect 8128 3040 8156 3139
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 8941 3179 8999 3185
rect 8941 3176 8953 3179
rect 8720 3148 8953 3176
rect 8720 3136 8726 3148
rect 8941 3145 8953 3148
rect 8987 3145 8999 3179
rect 8941 3139 8999 3145
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 9364 3148 9413 3176
rect 9364 3136 9370 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 8202 3068 8208 3120
rect 8260 3108 8266 3120
rect 8481 3111 8539 3117
rect 8481 3108 8493 3111
rect 8260 3080 8493 3108
rect 8260 3068 8266 3080
rect 8481 3077 8493 3080
rect 8527 3077 8539 3111
rect 8481 3071 8539 3077
rect 7331 3012 8156 3040
rect 7331 3009 7343 3012
rect 7285 3003 7343 3009
rect 4614 2972 4620 2984
rect 4575 2944 4620 2972
rect 4614 2932 4620 2944
rect 4672 2932 4678 2984
rect 4985 2975 5043 2981
rect 4985 2941 4997 2975
rect 5031 2972 5043 2975
rect 5626 2972 5632 2984
rect 5031 2944 5632 2972
rect 5031 2941 5043 2944
rect 4985 2935 5043 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 7021 2975 7079 2981
rect 7021 2941 7033 2975
rect 7067 2972 7079 2975
rect 7190 2972 7196 2984
rect 7067 2944 7196 2972
rect 7067 2941 7079 2944
rect 7021 2935 7079 2941
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 7607 2944 7941 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 7929 2941 7941 2944
rect 7975 2972 7987 2975
rect 8220 2972 8248 3068
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9306 3040 9312 3052
rect 9079 3012 9312 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 7975 2944 8248 2972
rect 8849 2975 8907 2981
rect 7975 2941 7987 2944
rect 7929 2935 7987 2941
rect 8849 2941 8861 2975
rect 8895 2972 8907 2975
rect 9214 2972 9220 2984
rect 8895 2944 9220 2972
rect 8895 2941 8907 2944
rect 8849 2935 8907 2941
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 4338 2836 4344 2848
rect 4299 2808 4344 2836
rect 4338 2796 4344 2808
rect 4396 2796 4402 2848
rect 3036 2746 9844 2768
rect 3036 2694 7566 2746
rect 7618 2694 7630 2746
rect 7682 2694 7694 2746
rect 7746 2694 7758 2746
rect 7810 2694 7822 2746
rect 7874 2694 9844 2746
rect 3036 2672 9844 2694
rect 4614 2592 4620 2644
rect 4672 2632 4678 2644
rect 4801 2635 4859 2641
rect 4801 2632 4813 2635
rect 4672 2604 4813 2632
rect 4672 2592 4678 2604
rect 4801 2601 4813 2604
rect 4847 2601 4859 2635
rect 5166 2632 5172 2644
rect 5127 2604 5172 2632
rect 4801 2595 4859 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 6086 2632 6092 2644
rect 6047 2604 6092 2632
rect 6086 2592 6092 2604
rect 6144 2592 6150 2644
rect 6546 2632 6552 2644
rect 6507 2604 6552 2632
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 7006 2632 7012 2644
rect 6967 2604 7012 2632
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2601 9091 2635
rect 9214 2632 9220 2644
rect 9175 2604 9220 2632
rect 9033 2595 9091 2601
rect 4522 2564 4528 2576
rect 3620 2536 4528 2564
rect 3620 2437 3648 2536
rect 3973 2499 4031 2505
rect 3973 2465 3985 2499
rect 4019 2496 4031 2499
rect 4154 2496 4160 2508
rect 4019 2468 4160 2496
rect 4019 2465 4031 2468
rect 3973 2459 4031 2465
rect 4154 2456 4160 2468
rect 4212 2456 4218 2508
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 3605 2431 3663 2437
rect 3605 2428 3617 2431
rect 3467 2400 3617 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 3605 2397 3617 2400
rect 3651 2397 3663 2431
rect 3605 2391 3663 2397
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2397 4123 2431
rect 4264 2428 4292 2536
rect 4522 2524 4528 2536
rect 4580 2564 4586 2576
rect 5258 2564 5264 2576
rect 4580 2536 5264 2564
rect 4580 2524 4586 2536
rect 5258 2524 5264 2536
rect 5316 2564 5322 2576
rect 5445 2567 5503 2573
rect 5445 2564 5457 2567
rect 5316 2536 5457 2564
rect 5316 2524 5322 2536
rect 5445 2533 5457 2536
rect 5491 2564 5503 2567
rect 6365 2567 6423 2573
rect 6365 2564 6377 2567
rect 5491 2536 6377 2564
rect 5491 2533 5503 2536
rect 5445 2527 5503 2533
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 4264 2400 4353 2428
rect 4065 2391 4123 2397
rect 4341 2397 4353 2400
rect 4387 2397 4399 2431
rect 4890 2428 4896 2440
rect 4851 2400 4896 2428
rect 4341 2391 4399 2397
rect 3234 2320 3240 2372
rect 3292 2360 3298 2372
rect 4080 2360 4108 2391
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 6196 2437 6224 2536
rect 6365 2533 6377 2536
rect 6411 2564 6423 2567
rect 6733 2567 6791 2573
rect 6733 2564 6745 2567
rect 6411 2536 6745 2564
rect 6411 2533 6423 2536
rect 6365 2527 6423 2533
rect 6733 2533 6745 2536
rect 6779 2564 6791 2567
rect 7193 2567 7251 2573
rect 7193 2564 7205 2567
rect 6779 2536 7205 2564
rect 6779 2533 6791 2536
rect 6733 2527 6791 2533
rect 7193 2533 7205 2536
rect 7239 2533 7251 2567
rect 8478 2564 8484 2576
rect 8439 2536 8484 2564
rect 7193 2527 7251 2533
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 7208 2428 7236 2527
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 9048 2564 9076 2595
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9582 2564 9588 2576
rect 9048 2536 9588 2564
rect 9582 2524 9588 2536
rect 9640 2524 9646 2576
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 9214 2496 9220 2508
rect 8352 2468 9220 2496
rect 8352 2456 8358 2468
rect 9214 2456 9220 2468
rect 9272 2496 9278 2508
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 9272 2468 9505 2496
rect 9272 2456 9278 2468
rect 9493 2465 9505 2468
rect 9539 2465 9551 2499
rect 9493 2459 9551 2465
rect 7561 2431 7619 2437
rect 7561 2428 7573 2431
rect 7208 2400 7573 2428
rect 6917 2391 6975 2397
rect 7561 2397 7573 2400
rect 7607 2397 7619 2431
rect 7834 2428 7840 2440
rect 7795 2400 7840 2428
rect 7561 2391 7619 2397
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 3292 2332 4169 2360
rect 3292 2320 3298 2332
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 4157 2323 4215 2329
rect 4525 2363 4583 2369
rect 4525 2329 4537 2363
rect 4571 2360 4583 2363
rect 5166 2360 5172 2372
rect 4571 2332 5172 2360
rect 4571 2329 4583 2332
rect 4525 2323 4583 2329
rect 4172 2292 4200 2323
rect 5166 2320 5172 2332
rect 5224 2320 5230 2372
rect 5920 2360 5948 2391
rect 5994 2360 6000 2372
rect 5907 2332 6000 2360
rect 5994 2320 6000 2332
rect 6052 2360 6058 2372
rect 6546 2360 6552 2372
rect 6052 2332 6552 2360
rect 6052 2320 6058 2332
rect 6546 2320 6552 2332
rect 6604 2320 6610 2372
rect 4430 2292 4436 2304
rect 4172 2264 4436 2292
rect 4430 2252 4436 2264
rect 4488 2252 4494 2304
rect 4890 2252 4896 2304
rect 4948 2292 4954 2304
rect 6932 2292 6960 2391
rect 7576 2360 7604 2391
rect 7834 2388 7840 2400
rect 7892 2428 7898 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7892 2400 8125 2428
rect 7892 2388 7898 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8662 2428 8668 2440
rect 8575 2400 8668 2428
rect 8113 2391 8171 2397
rect 8662 2388 8668 2400
rect 8720 2428 8726 2440
rect 8938 2428 8944 2440
rect 8720 2400 8944 2428
rect 8720 2388 8726 2400
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 9398 2388 9404 2440
rect 9456 2388 9462 2440
rect 8294 2360 8300 2372
rect 7576 2332 8300 2360
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 9079 2363 9137 2369
rect 9079 2329 9091 2363
rect 9125 2360 9137 2363
rect 9416 2360 9444 2388
rect 9125 2332 9444 2360
rect 9125 2329 9137 2332
rect 9079 2323 9137 2329
rect 4948 2264 6960 2292
rect 4948 2252 4954 2264
rect 3036 2202 9844 2224
rect 3036 2150 3816 2202
rect 3868 2150 3880 2202
rect 3932 2150 3944 2202
rect 3996 2150 4008 2202
rect 4060 2150 4072 2202
rect 4124 2150 8816 2202
rect 8868 2150 8880 2202
rect 8932 2150 8944 2202
rect 8996 2150 9008 2202
rect 9060 2150 9072 2202
rect 9124 2150 9844 2202
rect 3036 2128 9844 2150
rect 4338 2088 4344 2100
rect 3344 2060 4344 2088
rect 3344 1961 3372 2060
rect 4338 2048 4344 2060
rect 4396 2048 4402 2100
rect 5718 2088 5724 2100
rect 5776 2097 5782 2100
rect 5687 2060 5724 2088
rect 5718 2048 5724 2060
rect 5776 2051 5787 2097
rect 5994 2088 6000 2100
rect 5955 2060 6000 2088
rect 5776 2048 5782 2051
rect 5994 2048 6000 2060
rect 6052 2048 6058 2100
rect 8294 2088 8300 2100
rect 8255 2060 8300 2088
rect 8294 2048 8300 2060
rect 8352 2088 8358 2100
rect 8573 2091 8631 2097
rect 8573 2088 8585 2091
rect 8352 2060 8585 2088
rect 8352 2048 8358 2060
rect 8573 2057 8585 2060
rect 8619 2057 8631 2091
rect 8573 2051 8631 2057
rect 8662 2048 8668 2100
rect 8720 2088 8726 2100
rect 8757 2091 8815 2097
rect 8757 2088 8769 2091
rect 8720 2060 8769 2088
rect 8720 2048 8726 2060
rect 8757 2057 8769 2060
rect 8803 2057 8815 2091
rect 9306 2088 9312 2100
rect 9267 2060 9312 2088
rect 8757 2051 8815 2057
rect 9306 2048 9312 2060
rect 9364 2048 9370 2100
rect 4154 1980 4160 2032
rect 4212 1980 4218 2032
rect 5534 1980 5540 2032
rect 5592 2020 5598 2032
rect 7285 2023 7343 2029
rect 7285 2020 7297 2023
rect 5592 1992 7297 2020
rect 5592 1980 5598 1992
rect 7285 1989 7297 1992
rect 7331 2020 7343 2023
rect 7834 2020 7840 2032
rect 7331 1992 7840 2020
rect 7331 1989 7343 1992
rect 7285 1983 7343 1989
rect 7834 1980 7840 1992
rect 7892 2020 7898 2032
rect 7929 2023 7987 2029
rect 7929 2020 7941 2023
rect 7892 1992 7941 2020
rect 7892 1980 7898 1992
rect 7929 1989 7941 1992
rect 7975 1989 7987 2023
rect 7929 1983 7987 1989
rect 9214 1980 9220 2032
rect 9272 2020 9278 2032
rect 9401 2023 9459 2029
rect 9401 2020 9413 2023
rect 9272 1992 9413 2020
rect 9272 1980 9278 1992
rect 9401 1989 9413 1992
rect 9447 1989 9459 2023
rect 9401 1983 9459 1989
rect 3329 1955 3387 1961
rect 3329 1921 3341 1955
rect 3375 1921 3387 1955
rect 5166 1952 5172 1964
rect 5127 1924 5172 1952
rect 3329 1915 3387 1921
rect 5166 1912 5172 1924
rect 5224 1912 5230 1964
rect 3697 1887 3755 1893
rect 3697 1853 3709 1887
rect 3743 1884 3755 1887
rect 4246 1884 4252 1896
rect 3743 1856 4252 1884
rect 3743 1853 3755 1856
rect 3697 1847 3755 1853
rect 4246 1844 4252 1856
rect 4304 1844 4310 1896
rect 9122 1884 9128 1896
rect 9083 1856 9128 1884
rect 9122 1844 9128 1856
rect 9180 1844 9186 1896
rect 8941 1819 8999 1825
rect 8941 1785 8953 1819
rect 8987 1816 8999 1819
rect 9582 1816 9588 1828
rect 8987 1788 9588 1816
rect 8987 1785 8999 1788
rect 8941 1779 8999 1785
rect 9582 1776 9588 1788
rect 9640 1776 9646 1828
rect 3036 1658 9844 1680
rect 3036 1606 7566 1658
rect 7618 1606 7630 1658
rect 7682 1606 7694 1658
rect 7746 1606 7758 1658
rect 7810 1606 7822 1658
rect 7874 1606 9844 1658
rect 3036 1584 9844 1606
rect 4430 1504 4436 1556
rect 4488 1544 4494 1556
rect 5353 1547 5411 1553
rect 5353 1544 5365 1547
rect 4488 1516 5365 1544
rect 4488 1504 4494 1516
rect 5353 1513 5365 1516
rect 5399 1513 5411 1547
rect 9398 1544 9404 1556
rect 9359 1516 9404 1544
rect 5353 1507 5411 1513
rect 9398 1504 9404 1516
rect 9456 1504 9462 1556
rect 5258 1476 5264 1488
rect 5219 1448 5264 1476
rect 5258 1436 5264 1448
rect 5316 1436 5322 1488
rect 5077 1343 5135 1349
rect 5077 1309 5089 1343
rect 5123 1340 5135 1343
rect 6178 1340 6184 1352
rect 5123 1312 6184 1340
rect 5123 1309 5135 1312
rect 5077 1303 5135 1309
rect 6178 1300 6184 1312
rect 6236 1300 6242 1352
rect 3789 1207 3847 1213
rect 3789 1173 3801 1207
rect 3835 1204 3847 1207
rect 4890 1204 4896 1216
rect 3835 1176 4896 1204
rect 3835 1173 3847 1176
rect 3789 1167 3847 1173
rect 4890 1164 4896 1176
rect 4948 1164 4954 1216
rect 3036 1114 9844 1136
rect 3036 1062 3816 1114
rect 3868 1062 3880 1114
rect 3932 1062 3944 1114
rect 3996 1062 4008 1114
rect 4060 1062 4072 1114
rect 4124 1062 8816 1114
rect 8868 1062 8880 1114
rect 8932 1062 8944 1114
rect 8996 1062 9008 1114
rect 9060 1062 9072 1114
rect 9124 1062 9844 1114
rect 3036 1040 9844 1062
<< via1 >>
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 7566 11398 7618 11450
rect 7630 11398 7682 11450
rect 7694 11398 7746 11450
rect 7758 11398 7810 11450
rect 7822 11398 7874 11450
rect 1768 11296 1820 11348
rect 4344 11296 4396 11348
rect 6920 11296 6972 11348
rect 8116 11296 8168 11348
rect 4804 11160 4856 11212
rect 6368 11160 6420 11212
rect 8024 11160 8076 11212
rect 3148 11024 3200 11076
rect 4344 11135 4396 11144
rect 2964 10999 3016 11008
rect 2964 10965 2973 10999
rect 2973 10965 3007 10999
rect 3007 10965 3016 10999
rect 2964 10956 3016 10965
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 5356 11092 5408 11144
rect 4252 11067 4304 11076
rect 4252 11033 4261 11067
rect 4261 11033 4295 11067
rect 4295 11033 4304 11067
rect 4252 11024 4304 11033
rect 6092 11092 6144 11144
rect 6828 11092 6880 11144
rect 7012 11024 7064 11076
rect 4436 10956 4488 11008
rect 5540 10956 5592 11008
rect 6092 10956 6144 11008
rect 6368 10999 6420 11008
rect 6368 10965 6377 10999
rect 6377 10965 6411 10999
rect 6411 10965 6420 10999
rect 6368 10956 6420 10965
rect 7656 10956 7708 11008
rect 16580 11024 16632 11076
rect 3816 10854 3868 10906
rect 3880 10854 3932 10906
rect 3944 10854 3996 10906
rect 4008 10854 4060 10906
rect 4072 10854 4124 10906
rect 8816 10854 8868 10906
rect 8880 10854 8932 10906
rect 8944 10854 8996 10906
rect 9008 10854 9060 10906
rect 9072 10854 9124 10906
rect 4804 10752 4856 10804
rect 4712 10684 4764 10736
rect 5356 10727 5408 10736
rect 5356 10693 5365 10727
rect 5365 10693 5399 10727
rect 5399 10693 5408 10727
rect 5356 10684 5408 10693
rect 2964 10616 3016 10668
rect 4344 10616 4396 10668
rect 5264 10616 5316 10668
rect 7012 10752 7064 10804
rect 8024 10752 8076 10804
rect 1584 10548 1636 10600
rect 1768 10412 1820 10464
rect 6368 10616 6420 10668
rect 8208 10684 8260 10736
rect 5724 10523 5776 10532
rect 5724 10489 5733 10523
rect 5733 10489 5767 10523
rect 5767 10489 5776 10523
rect 5724 10480 5776 10489
rect 6092 10548 6144 10600
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 7472 10480 7524 10532
rect 5172 10455 5224 10464
rect 5172 10421 5189 10455
rect 5189 10421 5223 10455
rect 5223 10421 5224 10455
rect 5172 10412 5224 10421
rect 5908 10455 5960 10464
rect 5908 10421 5917 10455
rect 5917 10421 5951 10455
rect 5951 10421 5960 10455
rect 5908 10412 5960 10421
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 7104 10455 7156 10464
rect 7104 10421 7113 10455
rect 7113 10421 7147 10455
rect 7147 10421 7156 10455
rect 7104 10412 7156 10421
rect 7196 10412 7248 10464
rect 16580 10412 16632 10464
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 7566 10310 7618 10362
rect 7630 10310 7682 10362
rect 7694 10310 7746 10362
rect 7758 10310 7810 10362
rect 7822 10310 7874 10362
rect 4712 10251 4764 10260
rect 4712 10217 4721 10251
rect 4721 10217 4755 10251
rect 4755 10217 4764 10251
rect 4712 10208 4764 10217
rect 8116 10208 8168 10260
rect 3148 10140 3200 10192
rect 5264 10183 5316 10192
rect 1492 10004 1544 10056
rect 3148 10004 3200 10056
rect 4436 10072 4488 10124
rect 4712 10004 4764 10056
rect 5264 10149 5273 10183
rect 5273 10149 5307 10183
rect 5307 10149 5316 10183
rect 5264 10140 5316 10149
rect 5540 10072 5592 10124
rect 8024 10072 8076 10124
rect 5816 10047 5868 10056
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 5816 10004 5868 10013
rect 7104 10004 7156 10056
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 6368 9936 6420 9988
rect 8300 9979 8352 9988
rect 8300 9945 8309 9979
rect 8309 9945 8343 9979
rect 8343 9945 8352 9979
rect 8300 9936 8352 9945
rect 8668 9936 8720 9988
rect 3700 9868 3752 9920
rect 4160 9868 4212 9920
rect 8576 9868 8628 9920
rect 3816 9766 3868 9818
rect 3880 9766 3932 9818
rect 3944 9766 3996 9818
rect 4008 9766 4060 9818
rect 4072 9766 4124 9818
rect 8816 9766 8868 9818
rect 8880 9766 8932 9818
rect 8944 9766 8996 9818
rect 9008 9766 9060 9818
rect 9072 9766 9124 9818
rect 1492 9664 1544 9716
rect 2320 9596 2372 9648
rect 5264 9664 5316 9716
rect 7472 9664 7524 9716
rect 8116 9664 8168 9716
rect 4252 9596 4304 9648
rect 1584 9460 1636 9512
rect 3700 9503 3752 9512
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 3700 9460 3752 9469
rect 4160 9460 4212 9512
rect 5724 9460 5776 9512
rect 5816 9460 5868 9512
rect 6736 9503 6788 9512
rect 6736 9469 6745 9503
rect 6745 9469 6779 9503
rect 6779 9469 6788 9503
rect 6736 9460 6788 9469
rect 940 9324 992 9376
rect 6092 9392 6144 9444
rect 8300 9596 8352 9648
rect 7196 9528 7248 9580
rect 8668 9528 8720 9580
rect 8024 9460 8076 9512
rect 8484 9324 8536 9376
rect 9588 9324 9640 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 7566 9222 7618 9274
rect 7630 9222 7682 9274
rect 7694 9222 7746 9274
rect 7758 9222 7810 9274
rect 7822 9222 7874 9274
rect 1952 9120 2004 9172
rect 2412 9120 2464 9172
rect 2964 9120 3016 9172
rect 6736 9120 6788 9172
rect 8208 9163 8260 9172
rect 8208 9129 8217 9163
rect 8217 9129 8251 9163
rect 8251 9129 8260 9163
rect 8208 9120 8260 9129
rect 9496 9163 9548 9172
rect 9496 9129 9505 9163
rect 9505 9129 9539 9163
rect 9539 9129 9548 9163
rect 9496 9120 9548 9129
rect 4344 9052 4396 9104
rect 4436 8984 4488 9036
rect 6828 8984 6880 9036
rect 2964 8916 3016 8968
rect 3608 8916 3660 8968
rect 4344 8916 4396 8968
rect 4160 8891 4212 8900
rect 2320 8780 2372 8832
rect 2780 8780 2832 8832
rect 4160 8857 4169 8891
rect 4169 8857 4203 8891
rect 4203 8857 4212 8891
rect 4160 8848 4212 8857
rect 4988 8916 5040 8968
rect 7012 8848 7064 8900
rect 8116 8848 8168 8900
rect 8668 8848 8720 8900
rect 16764 8984 16816 9036
rect 9312 8823 9364 8832
rect 9312 8789 9321 8823
rect 9321 8789 9355 8823
rect 9355 8789 9364 8823
rect 9312 8780 9364 8789
rect 16580 8780 16632 8832
rect 3816 8678 3868 8730
rect 3880 8678 3932 8730
rect 3944 8678 3996 8730
rect 4008 8678 4060 8730
rect 4072 8678 4124 8730
rect 8816 8678 8868 8730
rect 8880 8678 8932 8730
rect 8944 8678 8996 8730
rect 9008 8678 9060 8730
rect 9072 8678 9124 8730
rect 4528 8576 4580 8628
rect 5632 8576 5684 8628
rect 6000 8576 6052 8628
rect 8024 8619 8076 8628
rect 1768 8551 1820 8560
rect 1768 8517 1777 8551
rect 1777 8517 1811 8551
rect 1811 8517 1820 8551
rect 1768 8508 1820 8517
rect 2780 8508 2832 8560
rect 4712 8508 4764 8560
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 8392 8508 8444 8560
rect 8668 8508 8720 8560
rect 4620 8440 4672 8492
rect 5816 8440 5868 8492
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 8208 8440 8260 8492
rect 1492 8415 1544 8424
rect 1492 8381 1501 8415
rect 1501 8381 1535 8415
rect 1535 8381 1544 8415
rect 1492 8372 1544 8381
rect 5080 8372 5132 8424
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 9312 8372 9364 8424
rect 4804 8304 4856 8356
rect 6092 8304 6144 8356
rect 6828 8304 6880 8356
rect 8300 8304 8352 8356
rect 16580 8304 16632 8356
rect 3148 8236 3200 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 7566 8134 7618 8186
rect 7630 8134 7682 8186
rect 7694 8134 7746 8186
rect 7758 8134 7810 8186
rect 7822 8134 7874 8186
rect 2964 8032 3016 8084
rect 3608 8032 3660 8084
rect 4712 8075 4764 8084
rect 4712 8041 4721 8075
rect 4721 8041 4755 8075
rect 4755 8041 4764 8075
rect 4712 8032 4764 8041
rect 5080 8032 5132 8084
rect 9312 8032 9364 8084
rect 3700 8007 3752 8016
rect 3700 7973 3709 8007
rect 3709 7973 3743 8007
rect 3743 7973 3752 8007
rect 3700 7964 3752 7973
rect 9496 7964 9548 8016
rect 4804 7896 4856 7948
rect 5908 7896 5960 7948
rect 8576 7896 8628 7948
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 4528 7828 4580 7880
rect 4988 7828 5040 7880
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 8300 7828 8352 7880
rect 2780 7692 2832 7744
rect 8116 7760 8168 7812
rect 8668 7692 8720 7744
rect 16672 7760 16724 7812
rect 16580 7692 16632 7744
rect 3816 7590 3868 7642
rect 3880 7590 3932 7642
rect 3944 7590 3996 7642
rect 4008 7590 4060 7642
rect 4072 7590 4124 7642
rect 8816 7590 8868 7642
rect 8880 7590 8932 7642
rect 8944 7590 8996 7642
rect 9008 7590 9060 7642
rect 9072 7590 9124 7642
rect 3056 7488 3108 7540
rect 9220 7488 9272 7540
rect 3700 7420 3752 7472
rect 6000 7420 6052 7472
rect 6184 7463 6236 7472
rect 6184 7429 6193 7463
rect 6193 7429 6227 7463
rect 6227 7429 6236 7463
rect 6184 7420 6236 7429
rect 7932 7463 7984 7472
rect 7932 7429 7941 7463
rect 7941 7429 7975 7463
rect 7975 7429 7984 7463
rect 7932 7420 7984 7429
rect 8116 7420 8168 7472
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 2780 7352 2832 7361
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 4160 7352 4212 7404
rect 4988 7352 5040 7404
rect 5816 7327 5868 7336
rect 5816 7293 5825 7327
rect 5825 7293 5859 7327
rect 5859 7293 5868 7327
rect 5816 7284 5868 7293
rect 6552 7284 6604 7336
rect 8300 7284 8352 7336
rect 9312 7284 9364 7336
rect 6828 7216 6880 7268
rect 5908 7191 5960 7200
rect 5908 7157 5917 7191
rect 5917 7157 5951 7191
rect 5951 7157 5960 7191
rect 5908 7148 5960 7157
rect 6460 7148 6512 7200
rect 8576 7148 8628 7200
rect 8852 7148 8904 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 7566 7046 7618 7098
rect 7630 7046 7682 7098
rect 7694 7046 7746 7098
rect 7758 7046 7810 7098
rect 7822 7046 7874 7098
rect 3148 6944 3200 6996
rect 4804 6944 4856 6996
rect 7472 6987 7524 6996
rect 7472 6953 7489 6987
rect 7489 6953 7523 6987
rect 7523 6953 7524 6987
rect 7472 6944 7524 6953
rect 8852 6876 8904 6928
rect 1492 6783 1544 6792
rect 1492 6749 1501 6783
rect 1501 6749 1535 6783
rect 1535 6749 1544 6783
rect 1492 6740 1544 6749
rect 3056 6740 3108 6792
rect 3700 6740 3752 6792
rect 4528 6740 4580 6792
rect 5448 6783 5500 6792
rect 2412 6672 2464 6724
rect 4252 6672 4304 6724
rect 3148 6604 3200 6656
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 7472 6740 7524 6792
rect 8576 6783 8628 6792
rect 5908 6672 5960 6724
rect 6828 6604 6880 6656
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 9220 6740 9272 6792
rect 16580 6740 16632 6792
rect 8392 6672 8444 6724
rect 9312 6672 9364 6724
rect 9404 6604 9456 6656
rect 3816 6502 3868 6554
rect 3880 6502 3932 6554
rect 3944 6502 3996 6554
rect 4008 6502 4060 6554
rect 4072 6502 4124 6554
rect 8816 6502 8868 6554
rect 8880 6502 8932 6554
rect 8944 6502 8996 6554
rect 9008 6502 9060 6554
rect 9072 6502 9124 6554
rect 13820 6468 13872 6520
rect 16672 6468 16724 6520
rect 3056 6400 3108 6452
rect 7472 6400 7524 6452
rect 2412 6375 2464 6384
rect 2412 6341 2421 6375
rect 2421 6341 2455 6375
rect 2455 6341 2464 6375
rect 2412 6332 2464 6341
rect 4252 6332 4304 6384
rect 5448 6332 5500 6384
rect 7932 6400 7984 6452
rect 8668 6400 8720 6452
rect 8852 6400 8904 6452
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 6000 6264 6052 6316
rect 3148 6239 3200 6248
rect 3148 6205 3157 6239
rect 3157 6205 3191 6239
rect 3191 6205 3200 6239
rect 3148 6196 3200 6205
rect 5908 6239 5960 6248
rect 5908 6205 5917 6239
rect 5917 6205 5951 6239
rect 5951 6205 5960 6239
rect 5908 6196 5960 6205
rect 6552 6196 6604 6248
rect 8300 6196 8352 6248
rect 8576 6196 8628 6248
rect 8484 6128 8536 6180
rect 4988 6060 5040 6112
rect 5448 6060 5500 6112
rect 8576 6060 8628 6112
rect 9220 6332 9272 6384
rect 19432 6128 19484 6180
rect 9220 6060 9272 6112
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 7566 5958 7618 6010
rect 7630 5958 7682 6010
rect 7694 5958 7746 6010
rect 7758 5958 7810 6010
rect 7822 5958 7874 6010
rect 3148 5856 3200 5908
rect 4620 5856 4672 5908
rect 5908 5899 5960 5908
rect 5908 5865 5917 5899
rect 5917 5865 5951 5899
rect 5951 5865 5960 5899
rect 5908 5856 5960 5865
rect 6828 5856 6880 5908
rect 8484 5899 8536 5908
rect 8484 5865 8493 5899
rect 8493 5865 8527 5899
rect 8527 5865 8536 5899
rect 8484 5856 8536 5865
rect 8668 5856 8720 5908
rect 9220 5856 9272 5908
rect 1492 5720 1544 5772
rect 5724 5720 5776 5772
rect 6000 5720 6052 5772
rect 6460 5763 6512 5772
rect 6460 5729 6469 5763
rect 6469 5729 6503 5763
rect 6503 5729 6512 5763
rect 6460 5720 6512 5729
rect 8668 5720 8720 5772
rect 8852 5763 8904 5772
rect 8852 5729 8861 5763
rect 8861 5729 8895 5763
rect 8895 5729 8904 5763
rect 8852 5720 8904 5729
rect 3332 5652 3384 5704
rect 2320 5584 2372 5636
rect 3516 5516 3568 5568
rect 3792 5584 3844 5636
rect 4160 5516 4212 5568
rect 4528 5516 4580 5568
rect 8392 5584 8444 5636
rect 8484 5516 8536 5568
rect 9496 5627 9548 5636
rect 9496 5593 9505 5627
rect 9505 5593 9539 5627
rect 9539 5593 9548 5627
rect 9496 5584 9548 5593
rect 16580 5516 16632 5568
rect 3816 5414 3868 5466
rect 3880 5414 3932 5466
rect 3944 5414 3996 5466
rect 4008 5414 4060 5466
rect 4072 5414 4124 5466
rect 8816 5414 8868 5466
rect 8880 5414 8932 5466
rect 8944 5414 8996 5466
rect 9008 5414 9060 5466
rect 9072 5414 9124 5466
rect 7012 5312 7064 5364
rect 4160 5244 4212 5296
rect 8484 5244 8536 5296
rect 6000 5219 6052 5228
rect 6000 5185 6009 5219
rect 6009 5185 6043 5219
rect 6043 5185 6052 5219
rect 6000 5176 6052 5185
rect 8300 5176 8352 5228
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 3332 5151 3384 5160
rect 3332 5117 3341 5151
rect 3341 5117 3375 5151
rect 3375 5117 3384 5151
rect 3332 5108 3384 5117
rect 3608 5151 3660 5160
rect 3608 5117 3617 5151
rect 3617 5117 3651 5151
rect 3651 5117 3660 5151
rect 3608 5108 3660 5117
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 6920 5108 6972 5160
rect 5172 4972 5224 5024
rect 8392 4972 8444 5024
rect 7566 4870 7618 4922
rect 7630 4870 7682 4922
rect 7694 4870 7746 4922
rect 7758 4870 7810 4922
rect 7822 4870 7874 4922
rect 5816 4768 5868 4820
rect 9220 4768 9272 4820
rect 5172 4700 5224 4752
rect 4160 4632 4212 4684
rect 5724 4675 5776 4684
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 9588 4632 9640 4684
rect 3332 4607 3384 4616
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 3332 4564 3384 4573
rect 4988 4564 5040 4616
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7012 4564 7064 4616
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 4620 4496 4672 4548
rect 7472 4496 7524 4548
rect 8300 4496 8352 4548
rect 9588 4496 9640 4548
rect 4252 4428 4304 4480
rect 9220 4471 9272 4480
rect 9220 4437 9229 4471
rect 9229 4437 9263 4471
rect 9263 4437 9272 4471
rect 9220 4428 9272 4437
rect 3816 4326 3868 4378
rect 3880 4326 3932 4378
rect 3944 4326 3996 4378
rect 4008 4326 4060 4378
rect 4072 4326 4124 4378
rect 8816 4326 8868 4378
rect 8880 4326 8932 4378
rect 8944 4326 8996 4378
rect 9008 4326 9060 4378
rect 9072 4326 9124 4378
rect 6552 4224 6604 4276
rect 5816 4156 5868 4208
rect 3240 4088 3292 4140
rect 5356 4131 5408 4140
rect 3608 4020 3660 4072
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 5448 4088 5500 4140
rect 9220 4088 9272 4140
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 4160 4020 4212 4072
rect 2688 3952 2740 4004
rect 6920 4020 6972 4072
rect 8668 4020 8720 4072
rect 5448 3952 5500 4004
rect 13820 3952 13872 4004
rect 5908 3927 5960 3936
rect 5908 3893 5925 3927
rect 5925 3893 5959 3927
rect 5959 3893 5960 3927
rect 5908 3884 5960 3893
rect 8392 3884 8444 3936
rect 7566 3782 7618 3834
rect 7630 3782 7682 3834
rect 7694 3782 7746 3834
rect 7758 3782 7810 3834
rect 7822 3782 7874 3834
rect 5356 3680 5408 3732
rect 5816 3723 5868 3732
rect 5816 3689 5825 3723
rect 5825 3689 5859 3723
rect 5859 3689 5868 3723
rect 5816 3680 5868 3689
rect 3332 3544 3384 3596
rect 5632 3544 5684 3596
rect 6552 3544 6604 3596
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 6920 3544 6972 3596
rect 4344 3408 4396 3460
rect 5172 3451 5224 3460
rect 5172 3417 5181 3451
rect 5181 3417 5215 3451
rect 5215 3417 5224 3451
rect 5172 3408 5224 3417
rect 4620 3340 4672 3392
rect 5448 3408 5500 3460
rect 6460 3408 6512 3460
rect 7012 3476 7064 3528
rect 8484 3476 8536 3528
rect 6644 3408 6696 3460
rect 7932 3408 7984 3460
rect 8576 3408 8628 3460
rect 8668 3340 8720 3392
rect 16580 3408 16632 3460
rect 9404 3383 9456 3392
rect 9404 3349 9413 3383
rect 9413 3349 9447 3383
rect 9447 3349 9456 3383
rect 9404 3340 9456 3349
rect 3816 3238 3868 3290
rect 3880 3238 3932 3290
rect 3944 3238 3996 3290
rect 4008 3238 4060 3290
rect 4072 3238 4124 3290
rect 8816 3238 8868 3290
rect 8880 3238 8932 3290
rect 8944 3238 8996 3290
rect 9008 3238 9060 3290
rect 9072 3238 9124 3290
rect 4252 3136 4304 3188
rect 8392 3179 8444 3188
rect 4344 3068 4396 3120
rect 6092 3068 6144 3120
rect 7472 3111 7524 3120
rect 7472 3077 7481 3111
rect 7481 3077 7515 3111
rect 7515 3077 7524 3111
rect 7472 3068 7524 3077
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 4896 3000 4948 3052
rect 6460 3043 6512 3052
rect 6460 3009 6469 3043
rect 6469 3009 6503 3043
rect 6503 3009 6512 3043
rect 6460 3000 6512 3009
rect 6644 3000 6696 3052
rect 8392 3145 8401 3179
rect 8401 3145 8435 3179
rect 8435 3145 8444 3179
rect 8392 3136 8444 3145
rect 8668 3136 8720 3188
rect 9312 3136 9364 3188
rect 8208 3068 8260 3120
rect 4620 2975 4672 2984
rect 4620 2941 4629 2975
rect 4629 2941 4663 2975
rect 4663 2941 4672 2975
rect 4620 2932 4672 2941
rect 5632 2932 5684 2984
rect 7196 2932 7248 2984
rect 9312 3000 9364 3052
rect 9220 2932 9272 2984
rect 4344 2839 4396 2848
rect 4344 2805 4353 2839
rect 4353 2805 4387 2839
rect 4387 2805 4396 2839
rect 4344 2796 4396 2805
rect 7566 2694 7618 2746
rect 7630 2694 7682 2746
rect 7694 2694 7746 2746
rect 7758 2694 7810 2746
rect 7822 2694 7874 2746
rect 4620 2592 4672 2644
rect 5172 2635 5224 2644
rect 5172 2601 5181 2635
rect 5181 2601 5215 2635
rect 5215 2601 5224 2635
rect 5172 2592 5224 2601
rect 6092 2635 6144 2644
rect 6092 2601 6101 2635
rect 6101 2601 6135 2635
rect 6135 2601 6144 2635
rect 6092 2592 6144 2601
rect 6552 2635 6604 2644
rect 6552 2601 6561 2635
rect 6561 2601 6595 2635
rect 6595 2601 6604 2635
rect 6552 2592 6604 2601
rect 7012 2635 7064 2644
rect 7012 2601 7021 2635
rect 7021 2601 7055 2635
rect 7055 2601 7064 2635
rect 7012 2592 7064 2601
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 9220 2635 9272 2644
rect 4160 2456 4212 2508
rect 4528 2524 4580 2576
rect 5264 2567 5316 2576
rect 5264 2533 5273 2567
rect 5273 2533 5307 2567
rect 5307 2533 5316 2567
rect 5264 2524 5316 2533
rect 4896 2431 4948 2440
rect 3240 2320 3292 2372
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 8484 2567 8536 2576
rect 8484 2533 8493 2567
rect 8493 2533 8527 2567
rect 8527 2533 8536 2567
rect 8484 2524 8536 2533
rect 9220 2601 9229 2635
rect 9229 2601 9263 2635
rect 9263 2601 9272 2635
rect 9220 2592 9272 2601
rect 9588 2524 9640 2576
rect 8300 2456 8352 2508
rect 9220 2456 9272 2508
rect 7840 2431 7892 2440
rect 5172 2320 5224 2372
rect 6000 2320 6052 2372
rect 6552 2320 6604 2372
rect 4436 2252 4488 2304
rect 4896 2252 4948 2304
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 8944 2388 8996 2440
rect 9404 2388 9456 2440
rect 8300 2363 8352 2372
rect 8300 2329 8309 2363
rect 8309 2329 8343 2363
rect 8343 2329 8352 2363
rect 8300 2320 8352 2329
rect 3816 2150 3868 2202
rect 3880 2150 3932 2202
rect 3944 2150 3996 2202
rect 4008 2150 4060 2202
rect 4072 2150 4124 2202
rect 8816 2150 8868 2202
rect 8880 2150 8932 2202
rect 8944 2150 8996 2202
rect 9008 2150 9060 2202
rect 9072 2150 9124 2202
rect 4344 2048 4396 2100
rect 5724 2091 5776 2100
rect 5724 2057 5741 2091
rect 5741 2057 5775 2091
rect 5775 2057 5776 2091
rect 5724 2048 5776 2057
rect 6000 2091 6052 2100
rect 6000 2057 6009 2091
rect 6009 2057 6043 2091
rect 6043 2057 6052 2091
rect 6000 2048 6052 2057
rect 8300 2091 8352 2100
rect 8300 2057 8309 2091
rect 8309 2057 8343 2091
rect 8343 2057 8352 2091
rect 8300 2048 8352 2057
rect 8668 2048 8720 2100
rect 9312 2091 9364 2100
rect 9312 2057 9321 2091
rect 9321 2057 9355 2091
rect 9355 2057 9364 2091
rect 9312 2048 9364 2057
rect 4160 1980 4212 2032
rect 5540 1980 5592 2032
rect 7840 1980 7892 2032
rect 9220 1980 9272 2032
rect 5172 1955 5224 1964
rect 5172 1921 5181 1955
rect 5181 1921 5215 1955
rect 5215 1921 5224 1955
rect 5172 1912 5224 1921
rect 4252 1844 4304 1896
rect 9128 1887 9180 1896
rect 9128 1853 9137 1887
rect 9137 1853 9171 1887
rect 9171 1853 9180 1887
rect 9128 1844 9180 1853
rect 9588 1776 9640 1828
rect 7566 1606 7618 1658
rect 7630 1606 7682 1658
rect 7694 1606 7746 1658
rect 7758 1606 7810 1658
rect 7822 1606 7874 1658
rect 4436 1504 4488 1556
rect 9404 1547 9456 1556
rect 9404 1513 9413 1547
rect 9413 1513 9447 1547
rect 9447 1513 9456 1547
rect 9404 1504 9456 1513
rect 5264 1479 5316 1488
rect 5264 1445 5273 1479
rect 5273 1445 5307 1479
rect 5307 1445 5316 1479
rect 5264 1436 5316 1445
rect 6184 1300 6236 1352
rect 4896 1164 4948 1216
rect 3816 1062 3868 1114
rect 3880 1062 3932 1114
rect 3944 1062 3996 1114
rect 4008 1062 4060 1114
rect 4072 1062 4124 1114
rect 8816 1062 8868 1114
rect 8880 1062 8932 1114
rect 8944 1062 8996 1114
rect 9008 1062 9060 1114
rect 9072 1062 9124 1114
<< obsm1 >>
rect 24000 0 34000 13000
<< metal2 >>
rect 938 12200 994 13000
rect 1398 12322 1454 13000
rect 1398 12294 1808 12322
rect 1398 12200 1454 12294
rect 952 9382 980 12200
rect 1780 11354 1808 12294
rect 1858 12200 1914 13000
rect 2318 12322 2374 13000
rect 2318 12294 2452 12322
rect 2318 12200 2374 12294
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1504 9722 1532 9998
rect 1492 9716 1544 9722
rect 1492 9658 1544 9664
rect 940 9376 992 9382
rect 940 9318 992 9324
rect 1504 8430 1532 9658
rect 1596 9518 1624 10542
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1780 8566 1808 10406
rect 1872 9738 1900 12200
rect 1872 9710 1992 9738
rect 1964 9178 1992 9710
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2332 8838 2360 9590
rect 2424 9178 2452 12294
rect 2778 12200 2834 13000
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12322 4214 13000
rect 4158 12294 4568 12322
rect 4158 12200 4214 12294
rect 2792 11642 2820 12200
rect 2792 11614 3096 11642
rect 2566 11452 2874 11461
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11387 2874 11396
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2976 10674 3004 10950
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2566 10364 2874 10373
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10299 2874 10308
rect 2566 9276 2874 9285
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9211 2874 9220
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2976 8974 3004 9114
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2792 8566 2820 8774
rect 1768 8560 1820 8566
rect 1768 8502 1820 8508
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 1504 6798 1532 8366
rect 2566 8188 2874 8197
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8123 2874 8132
rect 2976 8090 3004 8910
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2792 7410 2820 7686
rect 3068 7546 3096 11614
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 3160 10198 3188 11018
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3160 10062 3188 10134
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2566 7100 2874 7109
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7035 2874 7044
rect 3068 6798 3096 7482
rect 3160 7410 3188 8230
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3160 7002 3188 7346
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 1504 5778 1532 6734
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2424 6390 2452 6666
rect 3068 6458 3096 6734
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 2320 5636 2372 5642
rect 2424 5624 2452 6326
rect 3160 6254 3188 6598
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 2566 6012 2874 6021
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5947 2874 5956
rect 3160 5914 3188 6190
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 2372 5596 2452 5624
rect 2320 5578 2372 5584
rect 3252 4146 3280 12200
rect 3712 10010 3740 12200
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4356 11150 4384 11290
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 3816 10908 4124 10917
rect 3816 10906 3822 10908
rect 3878 10906 3902 10908
rect 3958 10906 3982 10908
rect 4038 10906 4062 10908
rect 4118 10906 4124 10908
rect 3878 10854 3880 10906
rect 4060 10854 4062 10906
rect 3816 10852 3822 10854
rect 3878 10852 3902 10854
rect 3958 10852 3982 10854
rect 4038 10852 4062 10854
rect 4118 10852 4124 10854
rect 3816 10843 4124 10852
rect 3620 9982 3740 10010
rect 3620 8974 3648 9982
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3712 9518 3740 9862
rect 3816 9820 4124 9829
rect 3816 9818 3822 9820
rect 3878 9818 3902 9820
rect 3958 9818 3982 9820
rect 4038 9818 4062 9820
rect 4118 9818 4124 9820
rect 3878 9766 3880 9818
rect 4060 9766 4062 9818
rect 3816 9764 3822 9766
rect 3878 9764 3902 9766
rect 3958 9764 3982 9766
rect 4038 9764 4062 9766
rect 4118 9764 4124 9766
rect 3816 9755 4124 9764
rect 4172 9518 4200 9862
rect 4264 9654 4292 11018
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4356 9110 4384 10610
rect 4448 10130 4476 10950
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4448 9042 4476 10066
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 3816 8732 4124 8741
rect 3816 8730 3822 8732
rect 3878 8730 3902 8732
rect 3958 8730 3982 8732
rect 4038 8730 4062 8732
rect 4118 8730 4124 8732
rect 3878 8678 3880 8730
rect 4060 8678 4062 8730
rect 3816 8676 3822 8678
rect 3878 8676 3902 8678
rect 3958 8676 3982 8678
rect 4038 8676 4062 8678
rect 4118 8676 4124 8678
rect 3816 8667 4124 8676
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3620 7886 3648 8026
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3712 7478 3740 7958
rect 3816 7644 4124 7653
rect 3816 7642 3822 7644
rect 3878 7642 3902 7644
rect 3958 7642 3982 7644
rect 4038 7642 4062 7644
rect 4118 7642 4124 7644
rect 3878 7590 3880 7642
rect 4060 7590 4062 7642
rect 3816 7588 3822 7590
rect 3878 7588 3902 7590
rect 3958 7588 3982 7590
rect 4038 7588 4062 7590
rect 4118 7588 4124 7590
rect 3816 7579 4124 7588
rect 3700 7472 3752 7478
rect 3700 7414 3752 7420
rect 4172 7410 4200 8842
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3344 5166 3372 5646
rect 3712 5624 3740 6734
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 3816 6556 4124 6565
rect 3816 6554 3822 6556
rect 3878 6554 3902 6556
rect 3958 6554 3982 6556
rect 4038 6554 4062 6556
rect 4118 6554 4124 6556
rect 3878 6502 3880 6554
rect 4060 6502 4062 6554
rect 3816 6500 3822 6502
rect 3878 6500 3902 6502
rect 3958 6500 3982 6502
rect 4038 6500 4062 6502
rect 4118 6500 4124 6502
rect 3816 6491 4124 6500
rect 4264 6390 4292 6666
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 3792 5636 3844 5642
rect 3712 5596 3792 5624
rect 3792 5578 3844 5584
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3344 4622 3372 5102
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2700 3437 2728 3946
rect 2686 3428 2742 3437
rect 2686 3363 2742 3372
rect 3252 2378 3280 4082
rect 3344 3602 3372 4558
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3528 3058 3556 5510
rect 3816 5468 4124 5477
rect 3816 5466 3822 5468
rect 3878 5466 3902 5468
rect 3958 5466 3982 5468
rect 4038 5466 4062 5468
rect 4118 5466 4124 5468
rect 3878 5414 3880 5466
rect 4060 5414 4062 5466
rect 3816 5412 3822 5414
rect 3878 5412 3902 5414
rect 3958 5412 3982 5414
rect 4038 5412 4062 5414
rect 4118 5412 4124 5414
rect 3816 5403 4124 5412
rect 4172 5302 4200 5510
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3620 4078 3648 5102
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 3816 4380 4124 4389
rect 3816 4378 3822 4380
rect 3878 4378 3902 4380
rect 3958 4378 3982 4380
rect 4038 4378 4062 4380
rect 4118 4378 4124 4380
rect 3878 4326 3880 4378
rect 4060 4326 4062 4378
rect 3816 4324 3822 4326
rect 3878 4324 3902 4326
rect 3958 4324 3982 4326
rect 4038 4324 4062 4326
rect 4118 4324 4124 4326
rect 3816 4315 4124 4324
rect 4172 4078 4200 4626
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 3816 3292 4124 3301
rect 3816 3290 3822 3292
rect 3878 3290 3902 3292
rect 3958 3290 3982 3292
rect 4038 3290 4062 3292
rect 4118 3290 4124 3292
rect 3878 3238 3880 3290
rect 4060 3238 4062 3290
rect 3816 3236 3822 3238
rect 3878 3236 3902 3238
rect 3958 3236 3982 3238
rect 4038 3236 4062 3238
rect 4118 3236 4124 3238
rect 3816 3227 4124 3236
rect 4264 3194 4292 4422
rect 4356 3466 4384 8910
rect 4540 8634 4568 12294
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6458 12200 6514 13000
rect 9402 12336 9458 12345
rect 6564 12294 6960 12322
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4632 8498 4660 12200
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4816 10810 4844 11154
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4724 10266 4752 10678
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4712 10056 4764 10062
rect 4816 10044 4844 10746
rect 4764 10016 4844 10044
rect 4712 9998 4764 10004
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4724 8090 4752 8502
rect 4816 8362 4844 10016
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4816 7954 4844 8298
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4540 6798 4568 7822
rect 4816 7002 4844 7890
rect 5000 7886 5028 8910
rect 5092 8430 5120 12200
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5552 11098 5580 12200
rect 5368 10742 5396 11086
rect 5552 11070 5672 11098
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5000 7410 5028 7822
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 5574 4568 6734
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4632 5914 4660 6258
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4540 4570 4568 5510
rect 5000 4622 5028 6054
rect 4988 4616 5040 4622
rect 4908 4576 4988 4604
rect 4540 4554 4660 4570
rect 4540 4548 4672 4554
rect 4540 4542 4620 4548
rect 4620 4490 4672 4496
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 3816 2204 4124 2213
rect 3816 2202 3822 2204
rect 3878 2202 3902 2204
rect 3958 2202 3982 2204
rect 4038 2202 4062 2204
rect 4118 2202 4124 2204
rect 3878 2150 3880 2202
rect 4060 2150 4062 2202
rect 3816 2148 3822 2150
rect 3878 2148 3902 2150
rect 3958 2148 3982 2150
rect 4038 2148 4062 2150
rect 4118 2148 4124 2150
rect 3816 2139 4124 2148
rect 4172 2038 4200 2450
rect 4160 2032 4212 2038
rect 4160 1974 4212 1980
rect 4264 1902 4292 3130
rect 4356 3126 4384 3402
rect 4632 3398 4660 4490
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4344 3120 4396 3126
rect 4632 3074 4660 3334
rect 4344 3062 4396 3068
rect 4540 3046 4660 3074
rect 4908 3058 4936 4576
rect 4988 4558 5040 4564
rect 5092 3534 5120 8026
rect 5184 6914 5212 10406
rect 5276 10198 5304 10610
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5276 9722 5304 10134
rect 5552 10130 5580 10950
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5644 8786 5672 11070
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5736 9518 5764 10474
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5828 9518 5856 9998
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5552 8758 5672 8786
rect 5184 6886 5304 6914
rect 5276 5137 5304 6886
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5460 6390 5488 6734
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5460 5273 5488 6054
rect 5446 5264 5502 5273
rect 5446 5199 5502 5208
rect 5262 5128 5318 5137
rect 5262 5063 5318 5072
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5184 4758 5212 4966
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5460 4146 5488 4558
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5368 3738 5396 4082
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5460 3466 5488 3946
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 4896 3052 4948 3058
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2106 4384 2790
rect 4540 2582 4568 3046
rect 4896 2994 4948 3000
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4632 2650 4660 2926
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 4908 2446 4936 2994
rect 5184 2650 5212 3402
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 4908 2310 4936 2382
rect 5172 2372 5224 2378
rect 5172 2314 5224 2320
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4344 2100 4396 2106
rect 4344 2042 4396 2048
rect 4252 1896 4304 1902
rect 4252 1838 4304 1844
rect 4448 1562 4476 2246
rect 4436 1556 4488 1562
rect 4436 1498 4488 1504
rect 4908 1222 4936 2246
rect 5184 1970 5212 2314
rect 5172 1964 5224 1970
rect 5172 1906 5224 1912
rect 5276 1494 5304 2518
rect 5552 2038 5580 8758
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5644 3602 5672 8570
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5828 7342 5856 8434
rect 5920 7954 5948 10406
rect 6012 8634 6040 12200
rect 6472 12050 6500 12200
rect 6564 12050 6592 12294
rect 6472 12022 6592 12050
rect 6932 11354 6960 12294
rect 9402 12271 9458 12280
rect 7566 11452 7874 11461
rect 7566 11450 7572 11452
rect 7628 11450 7652 11452
rect 7708 11450 7732 11452
rect 7788 11450 7812 11452
rect 7868 11450 7874 11452
rect 7628 11398 7630 11450
rect 7810 11398 7812 11450
rect 7566 11396 7572 11398
rect 7628 11396 7652 11398
rect 7708 11396 7732 11398
rect 7788 11396 7812 11398
rect 7868 11396 7874 11398
rect 7566 11387 7874 11396
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6104 11014 6132 11086
rect 6380 11014 6408 11154
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6104 10606 6132 10950
rect 6380 10674 6408 10950
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6104 9450 6132 10542
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 9994 6408 10406
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6092 9444 6144 9450
rect 6092 9386 6144 9392
rect 6748 9178 6776 9454
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6840 9042 6868 11086
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7024 10810 7052 11018
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7668 10674 7696 10950
rect 8036 10810 8064 11154
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 7930 10704 7986 10713
rect 7656 10668 7708 10674
rect 7930 10639 7986 10648
rect 7656 10610 7708 10616
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7116 10062 7144 10406
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7208 9586 7236 10406
rect 7484 9722 7512 10474
rect 7566 10364 7874 10373
rect 7566 10362 7572 10364
rect 7628 10362 7652 10364
rect 7708 10362 7732 10364
rect 7788 10362 7812 10364
rect 7868 10362 7874 10364
rect 7628 10310 7630 10362
rect 7810 10310 7812 10362
rect 7566 10308 7572 10310
rect 7628 10308 7652 10310
rect 7708 10308 7732 10310
rect 7788 10308 7812 10310
rect 7868 10308 7874 10310
rect 7566 10299 7874 10308
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7566 9276 7874 9285
rect 7566 9274 7572 9276
rect 7628 9274 7652 9276
rect 7708 9274 7732 9276
rect 7788 9274 7812 9276
rect 7868 9274 7874 9276
rect 7628 9222 7630 9274
rect 7810 9222 7812 9274
rect 7566 9220 7572 9222
rect 7628 9220 7652 9222
rect 7708 9220 7732 9222
rect 7788 9220 7812 9222
rect 7868 9220 7874 9222
rect 7566 9211 7874 9220
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 6012 7478 6040 8434
rect 6840 8362 6868 8978
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5920 6730 5948 7142
rect 6104 6914 6132 8298
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6012 6886 6132 6914
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 6012 6322 6040 6886
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5920 5914 5948 6190
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6012 5778 6040 6258
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5736 4690 5764 5714
rect 6012 5234 6040 5714
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5828 4826 5856 5102
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5736 3074 5764 4626
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5828 3738 5856 4150
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5920 3505 5948 3878
rect 5906 3496 5962 3505
rect 5906 3431 5962 3440
rect 5644 3046 5764 3074
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 5644 2990 5672 3046
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 6104 2650 6132 3062
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 5722 2544 5778 2553
rect 5722 2479 5778 2488
rect 5736 2106 5764 2479
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 6012 2106 6040 2314
rect 5724 2100 5776 2106
rect 5724 2042 5776 2048
rect 6000 2100 6052 2106
rect 6000 2042 6052 2048
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 5264 1488 5316 1494
rect 5264 1430 5316 1436
rect 6196 1358 6224 7414
rect 6472 7206 6500 7822
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 5778 6500 7142
rect 6564 6254 6592 7278
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 6840 6662 6868 7210
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6840 5914 6868 6598
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 7024 5370 7052 8842
rect 7566 8188 7874 8197
rect 7566 8186 7572 8188
rect 7628 8186 7652 8188
rect 7708 8186 7732 8188
rect 7788 8186 7812 8188
rect 7868 8186 7874 8188
rect 7628 8134 7630 8186
rect 7810 8134 7812 8186
rect 7566 8132 7572 8134
rect 7628 8132 7652 8134
rect 7708 8132 7732 8134
rect 7788 8132 7812 8134
rect 7868 8132 7874 8134
rect 7566 8123 7874 8132
rect 7944 7478 7972 10639
rect 8036 10130 8064 10746
rect 8128 10266 8156 11290
rect 8816 10908 9124 10917
rect 8816 10906 8822 10908
rect 8878 10906 8902 10908
rect 8958 10906 8982 10908
rect 9038 10906 9062 10908
rect 9118 10906 9124 10908
rect 8878 10854 8880 10906
rect 9060 10854 9062 10906
rect 8816 10852 8822 10854
rect 8878 10852 8902 10854
rect 8958 10852 8982 10854
rect 9038 10852 9062 10854
rect 9118 10852 9124 10854
rect 8816 10843 9124 10852
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8128 10062 8156 10202
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8036 8634 8064 9454
rect 8128 8906 8156 9658
rect 8220 9178 8248 10678
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8668 9988 8720 9994
rect 8668 9930 8720 9936
rect 8312 9654 8340 9930
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8220 8498 8248 9114
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8312 7886 8340 8298
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8128 7478 8156 7754
rect 7932 7472 7984 7478
rect 7470 7440 7526 7449
rect 7932 7414 7984 7420
rect 8116 7472 8168 7478
rect 8404 7426 8432 8502
rect 8116 7414 8168 7420
rect 7470 7375 7526 7384
rect 7484 7002 7512 7375
rect 7566 7100 7874 7109
rect 7566 7098 7572 7100
rect 7628 7098 7652 7100
rect 7708 7098 7732 7100
rect 7788 7098 7812 7100
rect 7868 7098 7874 7100
rect 7628 7046 7630 7098
rect 7810 7046 7812 7098
rect 7566 7044 7572 7046
rect 7628 7044 7652 7046
rect 7708 7044 7732 7046
rect 7788 7044 7812 7046
rect 7868 7044 7874 7046
rect 7566 7035 7874 7044
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7484 6458 7512 6734
rect 7944 6458 7972 7414
rect 8220 7398 8432 7426
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 8220 6066 8248 7398
rect 8300 7336 8352 7342
rect 8496 7324 8524 9318
rect 8588 7954 8616 9862
rect 8680 9586 8708 9930
rect 8816 9820 9124 9829
rect 8816 9818 8822 9820
rect 8878 9818 8902 9820
rect 8958 9818 8982 9820
rect 9038 9818 9062 9820
rect 9118 9818 9124 9820
rect 8878 9766 8880 9818
rect 9060 9766 9062 9818
rect 8816 9764 8822 9766
rect 8878 9764 8902 9766
rect 8958 9764 8982 9766
rect 9038 9764 9062 9766
rect 9118 9764 9124 9766
rect 8816 9755 9124 9764
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8680 8566 8708 8842
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 8816 8732 9124 8741
rect 8816 8730 8822 8732
rect 8878 8730 8902 8732
rect 8958 8730 8982 8732
rect 9038 8730 9062 8732
rect 9118 8730 9124 8732
rect 8878 8678 8880 8730
rect 9060 8678 9062 8730
rect 8816 8676 8822 8678
rect 8878 8676 8902 8678
rect 8958 8676 8982 8678
rect 9038 8676 9062 8678
rect 9118 8676 9124 8678
rect 8816 8667 9124 8676
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9232 8265 9260 8434
rect 9324 8430 9352 8774
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9218 8256 9274 8265
rect 9218 8191 9274 8200
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8300 7278 8352 7284
rect 8404 7296 8524 7324
rect 8312 6254 8340 7278
rect 8404 6914 8432 7296
rect 8588 7206 8616 7890
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8404 6886 8616 6914
rect 8588 6798 8616 6886
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8220 6038 8340 6066
rect 7566 6012 7874 6021
rect 7566 6010 7572 6012
rect 7628 6010 7652 6012
rect 7708 6010 7732 6012
rect 7788 6010 7812 6012
rect 7868 6010 7874 6012
rect 7628 5958 7630 6010
rect 7810 5958 7812 6010
rect 7566 5956 7572 5958
rect 7628 5956 7652 5958
rect 7708 5956 7732 5958
rect 7788 5956 7812 5958
rect 7868 5956 7874 5958
rect 7566 5947 7874 5956
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 4282 6592 4558
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6932 4078 6960 5102
rect 7024 4622 7052 5306
rect 8312 5234 8340 6038
rect 8404 5642 8432 6666
rect 8588 6338 8616 6734
rect 8680 6458 8708 7686
rect 8816 7644 9124 7653
rect 8816 7642 8822 7644
rect 8878 7642 8902 7644
rect 8958 7642 8982 7644
rect 9038 7642 9062 7644
rect 9118 7642 9124 7644
rect 8878 7590 8880 7642
rect 9060 7590 9062 7642
rect 8816 7588 8822 7590
rect 8878 7588 8902 7590
rect 8958 7588 8982 7590
rect 9038 7588 9062 7590
rect 9118 7588 9124 7590
rect 8816 7579 9124 7588
rect 9232 7546 9260 8191
rect 9324 8090 9352 8366
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9324 7342 9352 8026
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8864 6934 8892 7142
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 8816 6556 9124 6565
rect 8816 6554 8822 6556
rect 8878 6554 8902 6556
rect 8958 6554 8982 6556
rect 9038 6554 9062 6556
rect 9118 6554 9124 6556
rect 8878 6502 8880 6554
rect 9060 6502 9062 6554
rect 8816 6500 8822 6502
rect 8878 6500 8902 6502
rect 8958 6500 8982 6502
rect 9038 6500 9062 6502
rect 9118 6500 9124 6502
rect 8816 6491 9124 6500
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8864 6338 8892 6394
rect 9232 6390 9260 6734
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 8588 6310 8892 6338
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 8576 6248 8628 6254
rect 8628 6208 8708 6236
rect 8576 6190 8628 6196
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 8496 5914 8524 6122
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5302 8524 5510
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 7566 4924 7874 4933
rect 7566 4922 7572 4924
rect 7628 4922 7652 4924
rect 7708 4922 7732 4924
rect 7788 4922 7812 4924
rect 7868 4922 7874 4924
rect 7628 4870 7630 4922
rect 7810 4870 7812 4922
rect 7566 4868 7572 4870
rect 7628 4868 7652 4870
rect 7708 4868 7732 4870
rect 7788 4868 7812 4870
rect 7868 4868 7874 4870
rect 7566 4859 7874 4868
rect 8312 4706 8340 5170
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8220 4678 8340 4706
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6932 3602 6960 4014
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 3058 6500 3402
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6564 2650 6592 3538
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6656 3058 6684 3402
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 7024 2650 7052 3470
rect 7484 3126 7512 4490
rect 7566 3836 7874 3845
rect 7566 3834 7572 3836
rect 7628 3834 7652 3836
rect 7708 3834 7732 3836
rect 7788 3834 7812 3836
rect 7868 3834 7874 3836
rect 7628 3782 7630 3834
rect 7810 3782 7812 3834
rect 7566 3780 7572 3782
rect 7628 3780 7652 3782
rect 7708 3780 7732 3782
rect 7788 3780 7812 3782
rect 7868 3780 7874 3782
rect 7566 3771 7874 3780
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7196 2984 7248 2990
rect 7194 2952 7196 2961
rect 7248 2952 7250 2961
rect 7194 2887 7250 2896
rect 7566 2748 7874 2757
rect 7566 2746 7572 2748
rect 7628 2746 7652 2748
rect 7708 2746 7732 2748
rect 7788 2746 7812 2748
rect 7868 2746 7874 2748
rect 7628 2694 7630 2746
rect 7810 2694 7812 2746
rect 7566 2692 7572 2694
rect 7628 2692 7652 2694
rect 7708 2692 7732 2694
rect 7788 2692 7812 2694
rect 7868 2692 7874 2694
rect 7566 2683 7874 2692
rect 7944 2650 7972 3402
rect 8220 3126 8248 4678
rect 8404 4622 8432 4966
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 6564 2378 6592 2586
rect 8312 2514 8340 4490
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8404 3194 8432 3878
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8496 2582 8524 3470
rect 8588 3466 8616 6054
rect 8680 5914 8708 6208
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9232 5914 9260 6054
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 8850 5808 8906 5817
rect 8668 5772 8720 5778
rect 8850 5743 8852 5752
rect 8668 5714 8720 5720
rect 8904 5743 8906 5752
rect 8852 5714 8904 5720
rect 8680 4078 8708 5714
rect 8816 5468 9124 5477
rect 8816 5466 8822 5468
rect 8878 5466 8902 5468
rect 8958 5466 8982 5468
rect 9038 5466 9062 5468
rect 9118 5466 9124 5468
rect 8878 5414 8880 5466
rect 9060 5414 9062 5466
rect 8816 5412 8822 5414
rect 8878 5412 8902 5414
rect 8958 5412 8982 5414
rect 9038 5412 9062 5414
rect 9118 5412 9124 5414
rect 8816 5403 9124 5412
rect 9232 5234 9260 5850
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9232 4826 9260 5170
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 8816 4380 9124 4389
rect 8816 4378 8822 4380
rect 8878 4378 8902 4380
rect 8958 4378 8982 4380
rect 9038 4378 9062 4380
rect 9118 4378 9124 4380
rect 8878 4326 8880 4378
rect 9060 4326 9062 4378
rect 8816 4324 8822 4326
rect 8878 4324 8902 4326
rect 8958 4324 8982 4326
rect 9038 4324 9062 4326
rect 9118 4324 9124 4326
rect 8816 4315 9124 4324
rect 9126 4176 9182 4185
rect 9232 4146 9260 4422
rect 9126 4111 9182 4120
rect 9220 4140 9272 4146
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8576 3460 8628 3466
rect 9140 3448 9168 4111
rect 9220 4082 9272 4088
rect 9140 3420 9260 3448
rect 8576 3402 8628 3408
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8680 3194 8708 3334
rect 8816 3292 9124 3301
rect 8816 3290 8822 3292
rect 8878 3290 8902 3292
rect 8958 3290 8982 3292
rect 9038 3290 9062 3292
rect 9118 3290 9124 3292
rect 8878 3238 8880 3290
rect 9060 3238 9062 3290
rect 8816 3236 8822 3238
rect 8878 3236 8902 3238
rect 8958 3236 8982 3238
rect 9038 3236 9062 3238
rect 9118 3236 9124 3238
rect 8816 3227 9124 3236
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 9232 3074 9260 3420
rect 9324 3194 9352 6666
rect 9416 6662 9444 12271
rect 9494 11928 9550 11937
rect 9494 11863 9550 11872
rect 9508 9178 9536 11863
rect 16854 11520 16910 11529
rect 16854 11455 16910 11464
rect 16578 11112 16634 11121
rect 16578 11047 16580 11056
rect 16632 11047 16634 11056
rect 16580 11018 16632 11024
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16592 10305 16620 10406
rect 16578 10296 16634 10305
rect 16578 10231 16634 10240
rect 16762 9888 16818 9897
rect 16762 9823 16818 9832
rect 16578 9480 16634 9489
rect 16578 9415 16634 9424
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9508 8022 9536 9114
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9416 4146 9444 6598
rect 9600 5896 9628 9318
rect 16592 8838 16620 9415
rect 16670 9072 16726 9081
rect 16776 9042 16804 9823
rect 16670 9007 16726 9016
rect 16764 9036 16816 9042
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16578 8664 16634 8673
rect 16578 8599 16634 8608
rect 16592 8362 16620 8599
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16578 7848 16634 7857
rect 16684 7818 16712 9007
rect 16764 8978 16816 8984
rect 16578 7783 16634 7792
rect 16672 7812 16724 7818
rect 16592 7750 16620 7783
rect 16672 7754 16724 7760
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16868 6914 16896 11455
rect 19430 7032 19486 7041
rect 19430 6967 19486 6976
rect 16684 6886 16896 6914
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16592 6633 16620 6734
rect 16578 6624 16634 6633
rect 16578 6559 16634 6568
rect 16684 6526 16712 6886
rect 13820 6520 13872 6526
rect 13820 6462 13872 6468
rect 16672 6520 16724 6526
rect 16672 6462 16724 6468
rect 9600 5868 9720 5896
rect 9586 5808 9642 5817
rect 9586 5743 9642 5752
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 8956 3046 9260 3074
rect 9312 3052 9364 3058
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8956 2446 8984 3046
rect 9312 2994 9364 3000
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9232 2650 9260 2926
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 7852 2038 7880 2382
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8312 2106 8340 2314
rect 8680 2106 8708 2382
rect 8816 2204 9124 2213
rect 8816 2202 8822 2204
rect 8878 2202 8902 2204
rect 8958 2202 8982 2204
rect 9038 2202 9062 2204
rect 9118 2202 9124 2204
rect 8878 2150 8880 2202
rect 9060 2150 9062 2202
rect 8816 2148 8822 2150
rect 8878 2148 8902 2150
rect 8958 2148 8982 2150
rect 9038 2148 9062 2150
rect 9118 2148 9124 2150
rect 8816 2139 9124 2148
rect 8300 2100 8352 2106
rect 8300 2042 8352 2048
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 9232 2038 9260 2450
rect 9324 2145 9352 2994
rect 9416 2446 9444 3334
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9310 2136 9366 2145
rect 9310 2071 9312 2080
rect 9364 2071 9366 2080
rect 9312 2042 9364 2048
rect 7840 2032 7892 2038
rect 7840 1974 7892 1980
rect 9220 2032 9272 2038
rect 9324 2011 9352 2042
rect 9220 1974 9272 1980
rect 9128 1896 9180 1902
rect 9128 1838 9180 1844
rect 7566 1660 7874 1669
rect 7566 1658 7572 1660
rect 7628 1658 7652 1660
rect 7708 1658 7732 1660
rect 7788 1658 7812 1660
rect 7868 1658 7874 1660
rect 7628 1606 7630 1658
rect 7810 1606 7812 1658
rect 7566 1604 7572 1606
rect 7628 1604 7652 1606
rect 7708 1604 7732 1606
rect 7788 1604 7812 1606
rect 7868 1604 7874 1606
rect 7566 1595 7874 1604
rect 6184 1352 6236 1358
rect 9140 1329 9168 1838
rect 9416 1737 9444 2382
rect 9402 1728 9458 1737
rect 9402 1663 9458 1672
rect 9416 1562 9444 1663
rect 9404 1556 9456 1562
rect 9404 1498 9456 1504
rect 6184 1294 6236 1300
rect 9126 1320 9182 1329
rect 9126 1255 9182 1264
rect 4896 1216 4948 1222
rect 4896 1158 4948 1164
rect 3816 1116 4124 1125
rect 3816 1114 3822 1116
rect 3878 1114 3902 1116
rect 3958 1114 3982 1116
rect 4038 1114 4062 1116
rect 4118 1114 4124 1116
rect 3878 1062 3880 1114
rect 4060 1062 4062 1114
rect 3816 1060 3822 1062
rect 3878 1060 3902 1062
rect 3958 1060 3982 1062
rect 4038 1060 4062 1062
rect 4118 1060 4124 1062
rect 3816 1051 4124 1060
rect 8816 1116 9124 1125
rect 8816 1114 8822 1116
rect 8878 1114 8902 1116
rect 8958 1114 8982 1116
rect 9038 1114 9062 1116
rect 9118 1114 9124 1116
rect 8878 1062 8880 1114
rect 9060 1062 9062 1114
rect 8816 1060 8822 1062
rect 8878 1060 8902 1062
rect 8958 1060 8982 1062
rect 9038 1060 9062 1062
rect 9118 1060 9124 1062
rect 8816 1051 9124 1060
rect 9508 921 9536 5578
rect 9600 4690 9628 5743
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9692 4593 9720 5868
rect 9678 4584 9734 4593
rect 9588 4548 9640 4554
rect 9678 4519 9734 4528
rect 9588 4490 9640 4496
rect 9600 4185 9628 4490
rect 9586 4176 9642 4185
rect 9586 4111 9642 4120
rect 9600 2582 9628 4111
rect 13832 4010 13860 6462
rect 16578 6216 16634 6225
rect 19444 6186 19472 6967
rect 16578 6151 16634 6160
rect 19432 6180 19484 6186
rect 16592 5574 16620 6151
rect 19432 6122 19484 6128
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 16578 3768 16634 3777
rect 16578 3703 16634 3712
rect 16592 3466 16620 3703
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9588 1828 9640 1834
rect 9588 1770 9640 1776
rect 9494 912 9550 921
rect 9494 847 9550 856
rect 9600 513 9628 1770
rect 9586 504 9642 513
rect 9586 439 9642 448
<< via2 >>
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 3822 10906 3878 10908
rect 3902 10906 3958 10908
rect 3982 10906 4038 10908
rect 4062 10906 4118 10908
rect 3822 10854 3868 10906
rect 3868 10854 3878 10906
rect 3902 10854 3932 10906
rect 3932 10854 3944 10906
rect 3944 10854 3958 10906
rect 3982 10854 3996 10906
rect 3996 10854 4008 10906
rect 4008 10854 4038 10906
rect 4062 10854 4072 10906
rect 4072 10854 4118 10906
rect 3822 10852 3878 10854
rect 3902 10852 3958 10854
rect 3982 10852 4038 10854
rect 4062 10852 4118 10854
rect 3822 9818 3878 9820
rect 3902 9818 3958 9820
rect 3982 9818 4038 9820
rect 4062 9818 4118 9820
rect 3822 9766 3868 9818
rect 3868 9766 3878 9818
rect 3902 9766 3932 9818
rect 3932 9766 3944 9818
rect 3944 9766 3958 9818
rect 3982 9766 3996 9818
rect 3996 9766 4008 9818
rect 4008 9766 4038 9818
rect 4062 9766 4072 9818
rect 4072 9766 4118 9818
rect 3822 9764 3878 9766
rect 3902 9764 3958 9766
rect 3982 9764 4038 9766
rect 4062 9764 4118 9766
rect 3822 8730 3878 8732
rect 3902 8730 3958 8732
rect 3982 8730 4038 8732
rect 4062 8730 4118 8732
rect 3822 8678 3868 8730
rect 3868 8678 3878 8730
rect 3902 8678 3932 8730
rect 3932 8678 3944 8730
rect 3944 8678 3958 8730
rect 3982 8678 3996 8730
rect 3996 8678 4008 8730
rect 4008 8678 4038 8730
rect 4062 8678 4072 8730
rect 4072 8678 4118 8730
rect 3822 8676 3878 8678
rect 3902 8676 3958 8678
rect 3982 8676 4038 8678
rect 4062 8676 4118 8678
rect 3822 7642 3878 7644
rect 3902 7642 3958 7644
rect 3982 7642 4038 7644
rect 4062 7642 4118 7644
rect 3822 7590 3868 7642
rect 3868 7590 3878 7642
rect 3902 7590 3932 7642
rect 3932 7590 3944 7642
rect 3944 7590 3958 7642
rect 3982 7590 3996 7642
rect 3996 7590 4008 7642
rect 4008 7590 4038 7642
rect 4062 7590 4072 7642
rect 4072 7590 4118 7642
rect 3822 7588 3878 7590
rect 3902 7588 3958 7590
rect 3982 7588 4038 7590
rect 4062 7588 4118 7590
rect 3822 6554 3878 6556
rect 3902 6554 3958 6556
rect 3982 6554 4038 6556
rect 4062 6554 4118 6556
rect 3822 6502 3868 6554
rect 3868 6502 3878 6554
rect 3902 6502 3932 6554
rect 3932 6502 3944 6554
rect 3944 6502 3958 6554
rect 3982 6502 3996 6554
rect 3996 6502 4008 6554
rect 4008 6502 4038 6554
rect 4062 6502 4072 6554
rect 4072 6502 4118 6554
rect 3822 6500 3878 6502
rect 3902 6500 3958 6502
rect 3982 6500 4038 6502
rect 4062 6500 4118 6502
rect 2686 3372 2742 3428
rect 3822 5466 3878 5468
rect 3902 5466 3958 5468
rect 3982 5466 4038 5468
rect 4062 5466 4118 5468
rect 3822 5414 3868 5466
rect 3868 5414 3878 5466
rect 3902 5414 3932 5466
rect 3932 5414 3944 5466
rect 3944 5414 3958 5466
rect 3982 5414 3996 5466
rect 3996 5414 4008 5466
rect 4008 5414 4038 5466
rect 4062 5414 4072 5466
rect 4072 5414 4118 5466
rect 3822 5412 3878 5414
rect 3902 5412 3958 5414
rect 3982 5412 4038 5414
rect 4062 5412 4118 5414
rect 3822 4378 3878 4380
rect 3902 4378 3958 4380
rect 3982 4378 4038 4380
rect 4062 4378 4118 4380
rect 3822 4326 3868 4378
rect 3868 4326 3878 4378
rect 3902 4326 3932 4378
rect 3932 4326 3944 4378
rect 3944 4326 3958 4378
rect 3982 4326 3996 4378
rect 3996 4326 4008 4378
rect 4008 4326 4038 4378
rect 4062 4326 4072 4378
rect 4072 4326 4118 4378
rect 3822 4324 3878 4326
rect 3902 4324 3958 4326
rect 3982 4324 4038 4326
rect 4062 4324 4118 4326
rect 3822 3290 3878 3292
rect 3902 3290 3958 3292
rect 3982 3290 4038 3292
rect 4062 3290 4118 3292
rect 3822 3238 3868 3290
rect 3868 3238 3878 3290
rect 3902 3238 3932 3290
rect 3932 3238 3944 3290
rect 3944 3238 3958 3290
rect 3982 3238 3996 3290
rect 3996 3238 4008 3290
rect 4008 3238 4038 3290
rect 4062 3238 4072 3290
rect 4072 3238 4118 3290
rect 3822 3236 3878 3238
rect 3902 3236 3958 3238
rect 3982 3236 4038 3238
rect 4062 3236 4118 3238
rect 3822 2202 3878 2204
rect 3902 2202 3958 2204
rect 3982 2202 4038 2204
rect 4062 2202 4118 2204
rect 3822 2150 3868 2202
rect 3868 2150 3878 2202
rect 3902 2150 3932 2202
rect 3932 2150 3944 2202
rect 3944 2150 3958 2202
rect 3982 2150 3996 2202
rect 3996 2150 4008 2202
rect 4008 2150 4038 2202
rect 4062 2150 4072 2202
rect 4072 2150 4118 2202
rect 3822 2148 3878 2150
rect 3902 2148 3958 2150
rect 3982 2148 4038 2150
rect 4062 2148 4118 2150
rect 5446 5208 5502 5264
rect 5262 5072 5318 5128
rect 9402 12280 9458 12336
rect 7572 11450 7628 11452
rect 7652 11450 7708 11452
rect 7732 11450 7788 11452
rect 7812 11450 7868 11452
rect 7572 11398 7618 11450
rect 7618 11398 7628 11450
rect 7652 11398 7682 11450
rect 7682 11398 7694 11450
rect 7694 11398 7708 11450
rect 7732 11398 7746 11450
rect 7746 11398 7758 11450
rect 7758 11398 7788 11450
rect 7812 11398 7822 11450
rect 7822 11398 7868 11450
rect 7572 11396 7628 11398
rect 7652 11396 7708 11398
rect 7732 11396 7788 11398
rect 7812 11396 7868 11398
rect 7930 10648 7986 10704
rect 7572 10362 7628 10364
rect 7652 10362 7708 10364
rect 7732 10362 7788 10364
rect 7812 10362 7868 10364
rect 7572 10310 7618 10362
rect 7618 10310 7628 10362
rect 7652 10310 7682 10362
rect 7682 10310 7694 10362
rect 7694 10310 7708 10362
rect 7732 10310 7746 10362
rect 7746 10310 7758 10362
rect 7758 10310 7788 10362
rect 7812 10310 7822 10362
rect 7822 10310 7868 10362
rect 7572 10308 7628 10310
rect 7652 10308 7708 10310
rect 7732 10308 7788 10310
rect 7812 10308 7868 10310
rect 7572 9274 7628 9276
rect 7652 9274 7708 9276
rect 7732 9274 7788 9276
rect 7812 9274 7868 9276
rect 7572 9222 7618 9274
rect 7618 9222 7628 9274
rect 7652 9222 7682 9274
rect 7682 9222 7694 9274
rect 7694 9222 7708 9274
rect 7732 9222 7746 9274
rect 7746 9222 7758 9274
rect 7758 9222 7788 9274
rect 7812 9222 7822 9274
rect 7822 9222 7868 9274
rect 7572 9220 7628 9222
rect 7652 9220 7708 9222
rect 7732 9220 7788 9222
rect 7812 9220 7868 9222
rect 5906 3440 5962 3496
rect 5722 2488 5778 2544
rect 7572 8186 7628 8188
rect 7652 8186 7708 8188
rect 7732 8186 7788 8188
rect 7812 8186 7868 8188
rect 7572 8134 7618 8186
rect 7618 8134 7628 8186
rect 7652 8134 7682 8186
rect 7682 8134 7694 8186
rect 7694 8134 7708 8186
rect 7732 8134 7746 8186
rect 7746 8134 7758 8186
rect 7758 8134 7788 8186
rect 7812 8134 7822 8186
rect 7822 8134 7868 8186
rect 7572 8132 7628 8134
rect 7652 8132 7708 8134
rect 7732 8132 7788 8134
rect 7812 8132 7868 8134
rect 8822 10906 8878 10908
rect 8902 10906 8958 10908
rect 8982 10906 9038 10908
rect 9062 10906 9118 10908
rect 8822 10854 8868 10906
rect 8868 10854 8878 10906
rect 8902 10854 8932 10906
rect 8932 10854 8944 10906
rect 8944 10854 8958 10906
rect 8982 10854 8996 10906
rect 8996 10854 9008 10906
rect 9008 10854 9038 10906
rect 9062 10854 9072 10906
rect 9072 10854 9118 10906
rect 8822 10852 8878 10854
rect 8902 10852 8958 10854
rect 8982 10852 9038 10854
rect 9062 10852 9118 10854
rect 7470 7384 7526 7440
rect 7572 7098 7628 7100
rect 7652 7098 7708 7100
rect 7732 7098 7788 7100
rect 7812 7098 7868 7100
rect 7572 7046 7618 7098
rect 7618 7046 7628 7098
rect 7652 7046 7682 7098
rect 7682 7046 7694 7098
rect 7694 7046 7708 7098
rect 7732 7046 7746 7098
rect 7746 7046 7758 7098
rect 7758 7046 7788 7098
rect 7812 7046 7822 7098
rect 7822 7046 7868 7098
rect 7572 7044 7628 7046
rect 7652 7044 7708 7046
rect 7732 7044 7788 7046
rect 7812 7044 7868 7046
rect 8822 9818 8878 9820
rect 8902 9818 8958 9820
rect 8982 9818 9038 9820
rect 9062 9818 9118 9820
rect 8822 9766 8868 9818
rect 8868 9766 8878 9818
rect 8902 9766 8932 9818
rect 8932 9766 8944 9818
rect 8944 9766 8958 9818
rect 8982 9766 8996 9818
rect 8996 9766 9008 9818
rect 9008 9766 9038 9818
rect 9062 9766 9072 9818
rect 9072 9766 9118 9818
rect 8822 9764 8878 9766
rect 8902 9764 8958 9766
rect 8982 9764 9038 9766
rect 9062 9764 9118 9766
rect 8822 8730 8878 8732
rect 8902 8730 8958 8732
rect 8982 8730 9038 8732
rect 9062 8730 9118 8732
rect 8822 8678 8868 8730
rect 8868 8678 8878 8730
rect 8902 8678 8932 8730
rect 8932 8678 8944 8730
rect 8944 8678 8958 8730
rect 8982 8678 8996 8730
rect 8996 8678 9008 8730
rect 9008 8678 9038 8730
rect 9062 8678 9072 8730
rect 9072 8678 9118 8730
rect 8822 8676 8878 8678
rect 8902 8676 8958 8678
rect 8982 8676 9038 8678
rect 9062 8676 9118 8678
rect 9218 8200 9274 8256
rect 7572 6010 7628 6012
rect 7652 6010 7708 6012
rect 7732 6010 7788 6012
rect 7812 6010 7868 6012
rect 7572 5958 7618 6010
rect 7618 5958 7628 6010
rect 7652 5958 7682 6010
rect 7682 5958 7694 6010
rect 7694 5958 7708 6010
rect 7732 5958 7746 6010
rect 7746 5958 7758 6010
rect 7758 5958 7788 6010
rect 7812 5958 7822 6010
rect 7822 5958 7868 6010
rect 7572 5956 7628 5958
rect 7652 5956 7708 5958
rect 7732 5956 7788 5958
rect 7812 5956 7868 5958
rect 8822 7642 8878 7644
rect 8902 7642 8958 7644
rect 8982 7642 9038 7644
rect 9062 7642 9118 7644
rect 8822 7590 8868 7642
rect 8868 7590 8878 7642
rect 8902 7590 8932 7642
rect 8932 7590 8944 7642
rect 8944 7590 8958 7642
rect 8982 7590 8996 7642
rect 8996 7590 9008 7642
rect 9008 7590 9038 7642
rect 9062 7590 9072 7642
rect 9072 7590 9118 7642
rect 8822 7588 8878 7590
rect 8902 7588 8958 7590
rect 8982 7588 9038 7590
rect 9062 7588 9118 7590
rect 8822 6554 8878 6556
rect 8902 6554 8958 6556
rect 8982 6554 9038 6556
rect 9062 6554 9118 6556
rect 8822 6502 8868 6554
rect 8868 6502 8878 6554
rect 8902 6502 8932 6554
rect 8932 6502 8944 6554
rect 8944 6502 8958 6554
rect 8982 6502 8996 6554
rect 8996 6502 9008 6554
rect 9008 6502 9038 6554
rect 9062 6502 9072 6554
rect 9072 6502 9118 6554
rect 8822 6500 8878 6502
rect 8902 6500 8958 6502
rect 8982 6500 9038 6502
rect 9062 6500 9118 6502
rect 7572 4922 7628 4924
rect 7652 4922 7708 4924
rect 7732 4922 7788 4924
rect 7812 4922 7868 4924
rect 7572 4870 7618 4922
rect 7618 4870 7628 4922
rect 7652 4870 7682 4922
rect 7682 4870 7694 4922
rect 7694 4870 7708 4922
rect 7732 4870 7746 4922
rect 7746 4870 7758 4922
rect 7758 4870 7788 4922
rect 7812 4870 7822 4922
rect 7822 4870 7868 4922
rect 7572 4868 7628 4870
rect 7652 4868 7708 4870
rect 7732 4868 7788 4870
rect 7812 4868 7868 4870
rect 7572 3834 7628 3836
rect 7652 3834 7708 3836
rect 7732 3834 7788 3836
rect 7812 3834 7868 3836
rect 7572 3782 7618 3834
rect 7618 3782 7628 3834
rect 7652 3782 7682 3834
rect 7682 3782 7694 3834
rect 7694 3782 7708 3834
rect 7732 3782 7746 3834
rect 7746 3782 7758 3834
rect 7758 3782 7788 3834
rect 7812 3782 7822 3834
rect 7822 3782 7868 3834
rect 7572 3780 7628 3782
rect 7652 3780 7708 3782
rect 7732 3780 7788 3782
rect 7812 3780 7868 3782
rect 7194 2932 7196 2952
rect 7196 2932 7248 2952
rect 7248 2932 7250 2952
rect 7194 2896 7250 2932
rect 7572 2746 7628 2748
rect 7652 2746 7708 2748
rect 7732 2746 7788 2748
rect 7812 2746 7868 2748
rect 7572 2694 7618 2746
rect 7618 2694 7628 2746
rect 7652 2694 7682 2746
rect 7682 2694 7694 2746
rect 7694 2694 7708 2746
rect 7732 2694 7746 2746
rect 7746 2694 7758 2746
rect 7758 2694 7788 2746
rect 7812 2694 7822 2746
rect 7822 2694 7868 2746
rect 7572 2692 7628 2694
rect 7652 2692 7708 2694
rect 7732 2692 7788 2694
rect 7812 2692 7868 2694
rect 8850 5772 8906 5808
rect 8850 5752 8852 5772
rect 8852 5752 8904 5772
rect 8904 5752 8906 5772
rect 8822 5466 8878 5468
rect 8902 5466 8958 5468
rect 8982 5466 9038 5468
rect 9062 5466 9118 5468
rect 8822 5414 8868 5466
rect 8868 5414 8878 5466
rect 8902 5414 8932 5466
rect 8932 5414 8944 5466
rect 8944 5414 8958 5466
rect 8982 5414 8996 5466
rect 8996 5414 9008 5466
rect 9008 5414 9038 5466
rect 9062 5414 9072 5466
rect 9072 5414 9118 5466
rect 8822 5412 8878 5414
rect 8902 5412 8958 5414
rect 8982 5412 9038 5414
rect 9062 5412 9118 5414
rect 8822 4378 8878 4380
rect 8902 4378 8958 4380
rect 8982 4378 9038 4380
rect 9062 4378 9118 4380
rect 8822 4326 8868 4378
rect 8868 4326 8878 4378
rect 8902 4326 8932 4378
rect 8932 4326 8944 4378
rect 8944 4326 8958 4378
rect 8982 4326 8996 4378
rect 8996 4326 9008 4378
rect 9008 4326 9038 4378
rect 9062 4326 9072 4378
rect 9072 4326 9118 4378
rect 8822 4324 8878 4326
rect 8902 4324 8958 4326
rect 8982 4324 9038 4326
rect 9062 4324 9118 4326
rect 9126 4120 9182 4176
rect 8822 3290 8878 3292
rect 8902 3290 8958 3292
rect 8982 3290 9038 3292
rect 9062 3290 9118 3292
rect 8822 3238 8868 3290
rect 8868 3238 8878 3290
rect 8902 3238 8932 3290
rect 8932 3238 8944 3290
rect 8944 3238 8958 3290
rect 8982 3238 8996 3290
rect 8996 3238 9008 3290
rect 9008 3238 9038 3290
rect 9062 3238 9072 3290
rect 9072 3238 9118 3290
rect 8822 3236 8878 3238
rect 8902 3236 8958 3238
rect 8982 3236 9038 3238
rect 9062 3236 9118 3238
rect 9494 11872 9550 11928
rect 16854 11464 16910 11520
rect 16578 11076 16634 11112
rect 16578 11056 16580 11076
rect 16580 11056 16632 11076
rect 16632 11056 16634 11076
rect 16578 10240 16634 10296
rect 16762 9832 16818 9888
rect 16578 9424 16634 9480
rect 16670 9016 16726 9072
rect 16578 8608 16634 8664
rect 16578 7792 16634 7848
rect 19430 6976 19486 7032
rect 16578 6568 16634 6624
rect 9586 5752 9642 5808
rect 8822 2202 8878 2204
rect 8902 2202 8958 2204
rect 8982 2202 9038 2204
rect 9062 2202 9118 2204
rect 8822 2150 8868 2202
rect 8868 2150 8878 2202
rect 8902 2150 8932 2202
rect 8932 2150 8944 2202
rect 8944 2150 8958 2202
rect 8982 2150 8996 2202
rect 8996 2150 9008 2202
rect 9008 2150 9038 2202
rect 9062 2150 9072 2202
rect 9072 2150 9118 2202
rect 8822 2148 8878 2150
rect 8902 2148 8958 2150
rect 8982 2148 9038 2150
rect 9062 2148 9118 2150
rect 9310 2100 9366 2136
rect 9310 2080 9312 2100
rect 9312 2080 9364 2100
rect 9364 2080 9366 2100
rect 7572 1658 7628 1660
rect 7652 1658 7708 1660
rect 7732 1658 7788 1660
rect 7812 1658 7868 1660
rect 7572 1606 7618 1658
rect 7618 1606 7628 1658
rect 7652 1606 7682 1658
rect 7682 1606 7694 1658
rect 7694 1606 7708 1658
rect 7732 1606 7746 1658
rect 7746 1606 7758 1658
rect 7758 1606 7788 1658
rect 7812 1606 7822 1658
rect 7822 1606 7868 1658
rect 7572 1604 7628 1606
rect 7652 1604 7708 1606
rect 7732 1604 7788 1606
rect 7812 1604 7868 1606
rect 9402 1672 9458 1728
rect 9126 1264 9182 1320
rect 3822 1114 3878 1116
rect 3902 1114 3958 1116
rect 3982 1114 4038 1116
rect 4062 1114 4118 1116
rect 3822 1062 3868 1114
rect 3868 1062 3878 1114
rect 3902 1062 3932 1114
rect 3932 1062 3944 1114
rect 3944 1062 3958 1114
rect 3982 1062 3996 1114
rect 3996 1062 4008 1114
rect 4008 1062 4038 1114
rect 4062 1062 4072 1114
rect 4072 1062 4118 1114
rect 3822 1060 3878 1062
rect 3902 1060 3958 1062
rect 3982 1060 4038 1062
rect 4062 1060 4118 1062
rect 8822 1114 8878 1116
rect 8902 1114 8958 1116
rect 8982 1114 9038 1116
rect 9062 1114 9118 1116
rect 8822 1062 8868 1114
rect 8868 1062 8878 1114
rect 8902 1062 8932 1114
rect 8932 1062 8944 1114
rect 8944 1062 8958 1114
rect 8982 1062 8996 1114
rect 8996 1062 9008 1114
rect 9008 1062 9038 1114
rect 9062 1062 9072 1114
rect 9072 1062 9118 1114
rect 8822 1060 8878 1062
rect 8902 1060 8958 1062
rect 8982 1060 9038 1062
rect 9062 1060 9118 1062
rect 9678 4528 9734 4584
rect 9586 4120 9642 4176
rect 16578 6160 16634 6216
rect 16578 3712 16634 3768
rect 9494 856 9550 912
rect 9586 448 9642 504
<< obsm2 >>
rect 24000 0 34000 13000
<< metal3 >>
rect 9397 12338 9463 12341
rect 14000 12338 34000 12368
rect 9397 12336 34000 12338
rect 9397 12280 9402 12336
rect 9458 12280 34000 12336
rect 9397 12278 34000 12280
rect 9397 12275 9463 12278
rect 14000 12248 34000 12278
rect 9489 11930 9555 11933
rect 14000 11930 34000 11960
rect 9489 11928 34000 11930
rect 9489 11872 9494 11928
rect 9550 11872 34000 11928
rect 9489 11870 34000 11872
rect 9489 11867 9555 11870
rect 14000 11840 34000 11870
rect 14000 11520 34000 11552
rect 14000 11464 16854 11520
rect 16910 11464 34000 11520
rect 2562 11456 2878 11457
rect 2562 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2878 11456
rect 2562 11391 2878 11392
rect 7562 11456 7878 11457
rect 7562 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7878 11456
rect 14000 11432 34000 11464
rect 7562 11391 7878 11392
rect 14000 11112 34000 11144
rect 14000 11056 16578 11112
rect 16634 11056 34000 11112
rect 14000 11024 34000 11056
rect 3812 10912 4128 10913
rect 3812 10848 3818 10912
rect 3882 10848 3898 10912
rect 3962 10848 3978 10912
rect 4042 10848 4058 10912
rect 4122 10848 4128 10912
rect 3812 10847 4128 10848
rect 8812 10912 9128 10913
rect 8812 10848 8818 10912
rect 8882 10848 8898 10912
rect 8962 10848 8978 10912
rect 9042 10848 9058 10912
rect 9122 10848 9128 10912
rect 8812 10847 9128 10848
rect 7925 10706 7991 10709
rect 14000 10706 34000 10736
rect 7925 10704 34000 10706
rect 7925 10648 7930 10704
rect 7986 10648 34000 10704
rect 7925 10646 34000 10648
rect 7925 10643 7991 10646
rect 14000 10616 34000 10646
rect 2562 10368 2878 10369
rect 2562 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2878 10368
rect 2562 10303 2878 10304
rect 7562 10368 7878 10369
rect 7562 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7878 10368
rect 7562 10303 7878 10304
rect 14000 10296 34000 10328
rect 14000 10240 16578 10296
rect 16634 10240 34000 10296
rect 14000 10208 34000 10240
rect 14000 9888 34000 9920
rect 14000 9832 16762 9888
rect 16818 9832 34000 9888
rect 3812 9824 4128 9825
rect 3812 9760 3818 9824
rect 3882 9760 3898 9824
rect 3962 9760 3978 9824
rect 4042 9760 4058 9824
rect 4122 9760 4128 9824
rect 3812 9759 4128 9760
rect 8812 9824 9128 9825
rect 8812 9760 8818 9824
rect 8882 9760 8898 9824
rect 8962 9760 8978 9824
rect 9042 9760 9058 9824
rect 9122 9760 9128 9824
rect 14000 9800 34000 9832
rect 8812 9759 9128 9760
rect 14000 9480 34000 9512
rect 14000 9424 16578 9480
rect 16634 9424 34000 9480
rect 14000 9392 34000 9424
rect 2562 9280 2878 9281
rect 2562 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2878 9280
rect 2562 9215 2878 9216
rect 7562 9280 7878 9281
rect 7562 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7878 9280
rect 7562 9215 7878 9216
rect 14000 9072 34000 9104
rect 14000 9016 16670 9072
rect 16726 9016 34000 9072
rect 14000 8984 34000 9016
rect 3812 8736 4128 8737
rect 3812 8672 3818 8736
rect 3882 8672 3898 8736
rect 3962 8672 3978 8736
rect 4042 8672 4058 8736
rect 4122 8672 4128 8736
rect 3812 8671 4128 8672
rect 8812 8736 9128 8737
rect 8812 8672 8818 8736
rect 8882 8672 8898 8736
rect 8962 8672 8978 8736
rect 9042 8672 9058 8736
rect 9122 8672 9128 8736
rect 8812 8671 9128 8672
rect 14000 8664 34000 8696
rect 14000 8608 16578 8664
rect 16634 8608 34000 8664
rect 14000 8576 34000 8608
rect 9213 8258 9279 8261
rect 14000 8258 34000 8288
rect 9213 8256 34000 8258
rect 9213 8200 9218 8256
rect 9274 8200 34000 8256
rect 9213 8198 34000 8200
rect 9213 8195 9279 8198
rect 2562 8192 2878 8193
rect 2562 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2878 8192
rect 2562 8127 2878 8128
rect 7562 8192 7878 8193
rect 7562 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7878 8192
rect 14000 8168 34000 8198
rect 7562 8127 7878 8128
rect 14000 7848 34000 7880
rect 14000 7792 16578 7848
rect 16634 7792 34000 7848
rect 14000 7760 34000 7792
rect 3812 7648 4128 7649
rect 3812 7584 3818 7648
rect 3882 7584 3898 7648
rect 3962 7584 3978 7648
rect 4042 7584 4058 7648
rect 4122 7584 4128 7648
rect 3812 7583 4128 7584
rect 8812 7648 9128 7649
rect 8812 7584 8818 7648
rect 8882 7584 8898 7648
rect 8962 7584 8978 7648
rect 9042 7584 9058 7648
rect 9122 7584 9128 7648
rect 8812 7583 9128 7584
rect 7465 7442 7531 7445
rect 14000 7442 34000 7472
rect 7465 7440 34000 7442
rect 7465 7384 7470 7440
rect 7526 7384 34000 7440
rect 7465 7382 34000 7384
rect 7465 7379 7531 7382
rect 14000 7352 34000 7382
rect 2562 7104 2878 7105
rect 2562 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2878 7104
rect 2562 7039 2878 7040
rect 7562 7104 7878 7105
rect 7562 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7878 7104
rect 7562 7039 7878 7040
rect 14000 7032 34000 7064
rect 14000 6976 19430 7032
rect 19486 6976 34000 7032
rect 14000 6944 34000 6976
rect 14000 6624 34000 6656
rect 14000 6568 16578 6624
rect 16634 6568 34000 6624
rect 3812 6560 4128 6561
rect 3812 6496 3818 6560
rect 3882 6496 3898 6560
rect 3962 6496 3978 6560
rect 4042 6496 4058 6560
rect 4122 6496 4128 6560
rect 3812 6495 4128 6496
rect 8812 6560 9128 6561
rect 8812 6496 8818 6560
rect 8882 6496 8898 6560
rect 8962 6496 8978 6560
rect 9042 6496 9058 6560
rect 9122 6496 9128 6560
rect 14000 6536 34000 6568
rect 8812 6495 9128 6496
rect 14000 6216 34000 6248
rect 14000 6160 16578 6216
rect 16634 6160 34000 6216
rect 14000 6128 34000 6160
rect 2562 6016 2878 6017
rect 2562 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2878 6016
rect 2562 5951 2878 5952
rect 7562 6016 7878 6017
rect 7562 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7878 6016
rect 7562 5951 7878 5952
rect 8845 5810 8911 5813
rect 9581 5810 9647 5813
rect 14000 5810 34000 5840
rect 8845 5808 34000 5810
rect 8845 5752 8850 5808
rect 8906 5752 9586 5808
rect 9642 5752 34000 5808
rect 8845 5750 34000 5752
rect 8845 5747 8911 5750
rect 9581 5747 9647 5750
rect 14000 5720 34000 5750
rect 3812 5472 4128 5473
rect 3812 5408 3818 5472
rect 3882 5408 3898 5472
rect 3962 5408 3978 5472
rect 4042 5408 4058 5472
rect 4122 5408 4128 5472
rect 3812 5407 4128 5408
rect 8812 5472 9128 5473
rect 8812 5408 8818 5472
rect 8882 5408 8898 5472
rect 8962 5408 8978 5472
rect 9042 5408 9058 5472
rect 9122 5408 9128 5472
rect 8812 5407 9128 5408
rect 14000 5402 34000 5432
rect 10366 5342 34000 5402
rect 5441 5266 5507 5269
rect 10366 5266 10426 5342
rect 14000 5312 34000 5342
rect 5441 5264 10426 5266
rect 5441 5208 5446 5264
rect 5502 5208 10426 5264
rect 5441 5206 10426 5208
rect 5441 5203 5507 5206
rect 5257 5130 5323 5133
rect 5257 5128 9322 5130
rect 5257 5072 5262 5128
rect 5318 5072 9322 5128
rect 5257 5070 9322 5072
rect 5257 5067 5323 5070
rect 9262 4994 9322 5070
rect 14000 4994 34000 5024
rect 9262 4934 34000 4994
rect 7562 4928 7878 4929
rect 7562 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7878 4928
rect 14000 4904 34000 4934
rect 7562 4863 7878 4864
rect 9673 4586 9739 4589
rect 14000 4586 34000 4616
rect 9262 4584 34000 4586
rect 9262 4528 9678 4584
rect 9734 4528 34000 4584
rect 9262 4526 34000 4528
rect 3812 4384 4128 4385
rect 3812 4320 3818 4384
rect 3882 4320 3898 4384
rect 3962 4320 3978 4384
rect 4042 4320 4058 4384
rect 4122 4320 4128 4384
rect 3812 4319 4128 4320
rect 8812 4384 9128 4385
rect 8812 4320 8818 4384
rect 8882 4320 8898 4384
rect 8962 4320 8978 4384
rect 9042 4320 9058 4384
rect 9122 4320 9128 4384
rect 8812 4319 9128 4320
rect 9121 4178 9187 4181
rect 9262 4178 9322 4526
rect 9673 4523 9739 4526
rect 14000 4496 34000 4526
rect 9121 4176 9322 4178
rect 9121 4120 9126 4176
rect 9182 4120 9322 4176
rect 9121 4118 9322 4120
rect 9581 4178 9647 4181
rect 14000 4178 34000 4208
rect 9581 4176 34000 4178
rect 9581 4120 9586 4176
rect 9642 4120 34000 4176
rect 9581 4118 34000 4120
rect 9121 4115 9187 4118
rect 9581 4115 9647 4118
rect 14000 4088 34000 4118
rect 7562 3840 7878 3841
rect 7562 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7878 3840
rect 7562 3775 7878 3776
rect 14000 3768 34000 3800
rect 14000 3712 16578 3768
rect 16634 3712 34000 3768
rect 14000 3680 34000 3712
rect 5901 3498 5967 3501
rect 5901 3496 10426 3498
rect 5901 3440 5906 3496
rect 5962 3440 10426 3496
rect 5901 3438 10426 3440
rect 5901 3435 5967 3438
rect 2681 3430 2747 3433
rect 2484 3428 2747 3430
rect 2484 3372 2686 3428
rect 2742 3372 2747 3428
rect 2484 3370 2747 3372
rect 2681 3367 2747 3370
rect 10366 3362 10426 3438
rect 14000 3362 34000 3392
rect 10366 3302 34000 3362
rect 3812 3296 4128 3297
rect 3812 3232 3818 3296
rect 3882 3232 3898 3296
rect 3962 3232 3978 3296
rect 4042 3232 4058 3296
rect 4122 3232 4128 3296
rect 3812 3231 4128 3232
rect 8812 3296 9128 3297
rect 8812 3232 8818 3296
rect 8882 3232 8898 3296
rect 8962 3232 8978 3296
rect 9042 3232 9058 3296
rect 9122 3232 9128 3296
rect 14000 3272 34000 3302
rect 8812 3231 9128 3232
rect 7189 2954 7255 2957
rect 14000 2954 34000 2984
rect 7189 2952 34000 2954
rect 7189 2896 7194 2952
rect 7250 2896 34000 2952
rect 7189 2894 34000 2896
rect 7189 2891 7255 2894
rect 14000 2864 34000 2894
rect 7562 2752 7878 2753
rect 7562 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7878 2752
rect 7562 2687 7878 2688
rect 5717 2546 5783 2549
rect 14000 2546 34000 2576
rect 5717 2544 34000 2546
rect 5717 2488 5722 2544
rect 5778 2488 34000 2544
rect 5717 2486 34000 2488
rect 5717 2483 5783 2486
rect 14000 2456 34000 2486
rect 3812 2208 4128 2209
rect 3812 2144 3818 2208
rect 3882 2144 3898 2208
rect 3962 2144 3978 2208
rect 4042 2144 4058 2208
rect 4122 2144 4128 2208
rect 3812 2143 4128 2144
rect 8812 2208 9128 2209
rect 8812 2144 8818 2208
rect 8882 2144 8898 2208
rect 8962 2144 8978 2208
rect 9042 2144 9058 2208
rect 9122 2144 9128 2208
rect 8812 2143 9128 2144
rect 9305 2138 9371 2141
rect 14000 2138 34000 2168
rect 9305 2136 34000 2138
rect 9305 2080 9310 2136
rect 9366 2080 34000 2136
rect 9305 2078 34000 2080
rect 9305 2075 9371 2078
rect 14000 2048 34000 2078
rect 9397 1730 9463 1733
rect 14000 1730 34000 1760
rect 9397 1728 34000 1730
rect 9397 1672 9402 1728
rect 9458 1672 34000 1728
rect 9397 1670 34000 1672
rect 9397 1667 9463 1670
rect 7562 1664 7878 1665
rect 7562 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7878 1664
rect 14000 1640 34000 1670
rect 7562 1599 7878 1600
rect 9121 1322 9187 1325
rect 14000 1322 34000 1352
rect 9121 1320 34000 1322
rect 9121 1264 9126 1320
rect 9182 1264 34000 1320
rect 9121 1262 34000 1264
rect 9121 1259 9187 1262
rect 14000 1232 34000 1262
rect 3812 1120 4128 1121
rect 3812 1056 3818 1120
rect 3882 1056 3898 1120
rect 3962 1056 3978 1120
rect 4042 1056 4058 1120
rect 4122 1056 4128 1120
rect 3812 1055 4128 1056
rect 8812 1120 9128 1121
rect 8812 1056 8818 1120
rect 8882 1056 8898 1120
rect 8962 1056 8978 1120
rect 9042 1056 9058 1120
rect 9122 1056 9128 1120
rect 8812 1055 9128 1056
rect 9489 914 9555 917
rect 14000 914 34000 944
rect 9489 912 34000 914
rect 9489 856 9494 912
rect 9550 856 34000 912
rect 9489 854 34000 856
rect 9489 851 9555 854
rect 14000 824 34000 854
rect 9581 506 9647 509
rect 14000 506 34000 536
rect 9581 504 34000 506
rect 9581 448 9586 504
rect 9642 448 34000 504
rect 9581 446 34000 448
rect 9581 443 9647 446
rect 14000 416 34000 446
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 7568 11452 7632 11456
rect 7568 11396 7572 11452
rect 7572 11396 7628 11452
rect 7628 11396 7632 11452
rect 7568 11392 7632 11396
rect 7648 11452 7712 11456
rect 7648 11396 7652 11452
rect 7652 11396 7708 11452
rect 7708 11396 7712 11452
rect 7648 11392 7712 11396
rect 7728 11452 7792 11456
rect 7728 11396 7732 11452
rect 7732 11396 7788 11452
rect 7788 11396 7792 11452
rect 7728 11392 7792 11396
rect 7808 11452 7872 11456
rect 7808 11396 7812 11452
rect 7812 11396 7868 11452
rect 7868 11396 7872 11452
rect 7808 11392 7872 11396
rect 3818 10908 3882 10912
rect 3818 10852 3822 10908
rect 3822 10852 3878 10908
rect 3878 10852 3882 10908
rect 3818 10848 3882 10852
rect 3898 10908 3962 10912
rect 3898 10852 3902 10908
rect 3902 10852 3958 10908
rect 3958 10852 3962 10908
rect 3898 10848 3962 10852
rect 3978 10908 4042 10912
rect 3978 10852 3982 10908
rect 3982 10852 4038 10908
rect 4038 10852 4042 10908
rect 3978 10848 4042 10852
rect 4058 10908 4122 10912
rect 4058 10852 4062 10908
rect 4062 10852 4118 10908
rect 4118 10852 4122 10908
rect 4058 10848 4122 10852
rect 8818 10908 8882 10912
rect 8818 10852 8822 10908
rect 8822 10852 8878 10908
rect 8878 10852 8882 10908
rect 8818 10848 8882 10852
rect 8898 10908 8962 10912
rect 8898 10852 8902 10908
rect 8902 10852 8958 10908
rect 8958 10852 8962 10908
rect 8898 10848 8962 10852
rect 8978 10908 9042 10912
rect 8978 10852 8982 10908
rect 8982 10852 9038 10908
rect 9038 10852 9042 10908
rect 8978 10848 9042 10852
rect 9058 10908 9122 10912
rect 9058 10852 9062 10908
rect 9062 10852 9118 10908
rect 9118 10852 9122 10908
rect 9058 10848 9122 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 7568 10364 7632 10368
rect 7568 10308 7572 10364
rect 7572 10308 7628 10364
rect 7628 10308 7632 10364
rect 7568 10304 7632 10308
rect 7648 10364 7712 10368
rect 7648 10308 7652 10364
rect 7652 10308 7708 10364
rect 7708 10308 7712 10364
rect 7648 10304 7712 10308
rect 7728 10364 7792 10368
rect 7728 10308 7732 10364
rect 7732 10308 7788 10364
rect 7788 10308 7792 10364
rect 7728 10304 7792 10308
rect 7808 10364 7872 10368
rect 7808 10308 7812 10364
rect 7812 10308 7868 10364
rect 7868 10308 7872 10364
rect 7808 10304 7872 10308
rect 3818 9820 3882 9824
rect 3818 9764 3822 9820
rect 3822 9764 3878 9820
rect 3878 9764 3882 9820
rect 3818 9760 3882 9764
rect 3898 9820 3962 9824
rect 3898 9764 3902 9820
rect 3902 9764 3958 9820
rect 3958 9764 3962 9820
rect 3898 9760 3962 9764
rect 3978 9820 4042 9824
rect 3978 9764 3982 9820
rect 3982 9764 4038 9820
rect 4038 9764 4042 9820
rect 3978 9760 4042 9764
rect 4058 9820 4122 9824
rect 4058 9764 4062 9820
rect 4062 9764 4118 9820
rect 4118 9764 4122 9820
rect 4058 9760 4122 9764
rect 8818 9820 8882 9824
rect 8818 9764 8822 9820
rect 8822 9764 8878 9820
rect 8878 9764 8882 9820
rect 8818 9760 8882 9764
rect 8898 9820 8962 9824
rect 8898 9764 8902 9820
rect 8902 9764 8958 9820
rect 8958 9764 8962 9820
rect 8898 9760 8962 9764
rect 8978 9820 9042 9824
rect 8978 9764 8982 9820
rect 8982 9764 9038 9820
rect 9038 9764 9042 9820
rect 8978 9760 9042 9764
rect 9058 9820 9122 9824
rect 9058 9764 9062 9820
rect 9062 9764 9118 9820
rect 9118 9764 9122 9820
rect 9058 9760 9122 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 7568 9276 7632 9280
rect 7568 9220 7572 9276
rect 7572 9220 7628 9276
rect 7628 9220 7632 9276
rect 7568 9216 7632 9220
rect 7648 9276 7712 9280
rect 7648 9220 7652 9276
rect 7652 9220 7708 9276
rect 7708 9220 7712 9276
rect 7648 9216 7712 9220
rect 7728 9276 7792 9280
rect 7728 9220 7732 9276
rect 7732 9220 7788 9276
rect 7788 9220 7792 9276
rect 7728 9216 7792 9220
rect 7808 9276 7872 9280
rect 7808 9220 7812 9276
rect 7812 9220 7868 9276
rect 7868 9220 7872 9276
rect 7808 9216 7872 9220
rect 3818 8732 3882 8736
rect 3818 8676 3822 8732
rect 3822 8676 3878 8732
rect 3878 8676 3882 8732
rect 3818 8672 3882 8676
rect 3898 8732 3962 8736
rect 3898 8676 3902 8732
rect 3902 8676 3958 8732
rect 3958 8676 3962 8732
rect 3898 8672 3962 8676
rect 3978 8732 4042 8736
rect 3978 8676 3982 8732
rect 3982 8676 4038 8732
rect 4038 8676 4042 8732
rect 3978 8672 4042 8676
rect 4058 8732 4122 8736
rect 4058 8676 4062 8732
rect 4062 8676 4118 8732
rect 4118 8676 4122 8732
rect 4058 8672 4122 8676
rect 8818 8732 8882 8736
rect 8818 8676 8822 8732
rect 8822 8676 8878 8732
rect 8878 8676 8882 8732
rect 8818 8672 8882 8676
rect 8898 8732 8962 8736
rect 8898 8676 8902 8732
rect 8902 8676 8958 8732
rect 8958 8676 8962 8732
rect 8898 8672 8962 8676
rect 8978 8732 9042 8736
rect 8978 8676 8982 8732
rect 8982 8676 9038 8732
rect 9038 8676 9042 8732
rect 8978 8672 9042 8676
rect 9058 8732 9122 8736
rect 9058 8676 9062 8732
rect 9062 8676 9118 8732
rect 9118 8676 9122 8732
rect 9058 8672 9122 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 7568 8188 7632 8192
rect 7568 8132 7572 8188
rect 7572 8132 7628 8188
rect 7628 8132 7632 8188
rect 7568 8128 7632 8132
rect 7648 8188 7712 8192
rect 7648 8132 7652 8188
rect 7652 8132 7708 8188
rect 7708 8132 7712 8188
rect 7648 8128 7712 8132
rect 7728 8188 7792 8192
rect 7728 8132 7732 8188
rect 7732 8132 7788 8188
rect 7788 8132 7792 8188
rect 7728 8128 7792 8132
rect 7808 8188 7872 8192
rect 7808 8132 7812 8188
rect 7812 8132 7868 8188
rect 7868 8132 7872 8188
rect 7808 8128 7872 8132
rect 3818 7644 3882 7648
rect 3818 7588 3822 7644
rect 3822 7588 3878 7644
rect 3878 7588 3882 7644
rect 3818 7584 3882 7588
rect 3898 7644 3962 7648
rect 3898 7588 3902 7644
rect 3902 7588 3958 7644
rect 3958 7588 3962 7644
rect 3898 7584 3962 7588
rect 3978 7644 4042 7648
rect 3978 7588 3982 7644
rect 3982 7588 4038 7644
rect 4038 7588 4042 7644
rect 3978 7584 4042 7588
rect 4058 7644 4122 7648
rect 4058 7588 4062 7644
rect 4062 7588 4118 7644
rect 4118 7588 4122 7644
rect 4058 7584 4122 7588
rect 8818 7644 8882 7648
rect 8818 7588 8822 7644
rect 8822 7588 8878 7644
rect 8878 7588 8882 7644
rect 8818 7584 8882 7588
rect 8898 7644 8962 7648
rect 8898 7588 8902 7644
rect 8902 7588 8958 7644
rect 8958 7588 8962 7644
rect 8898 7584 8962 7588
rect 8978 7644 9042 7648
rect 8978 7588 8982 7644
rect 8982 7588 9038 7644
rect 9038 7588 9042 7644
rect 8978 7584 9042 7588
rect 9058 7644 9122 7648
rect 9058 7588 9062 7644
rect 9062 7588 9118 7644
rect 9118 7588 9122 7644
rect 9058 7584 9122 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 7568 7100 7632 7104
rect 7568 7044 7572 7100
rect 7572 7044 7628 7100
rect 7628 7044 7632 7100
rect 7568 7040 7632 7044
rect 7648 7100 7712 7104
rect 7648 7044 7652 7100
rect 7652 7044 7708 7100
rect 7708 7044 7712 7100
rect 7648 7040 7712 7044
rect 7728 7100 7792 7104
rect 7728 7044 7732 7100
rect 7732 7044 7788 7100
rect 7788 7044 7792 7100
rect 7728 7040 7792 7044
rect 7808 7100 7872 7104
rect 7808 7044 7812 7100
rect 7812 7044 7868 7100
rect 7868 7044 7872 7100
rect 7808 7040 7872 7044
rect 3818 6556 3882 6560
rect 3818 6500 3822 6556
rect 3822 6500 3878 6556
rect 3878 6500 3882 6556
rect 3818 6496 3882 6500
rect 3898 6556 3962 6560
rect 3898 6500 3902 6556
rect 3902 6500 3958 6556
rect 3958 6500 3962 6556
rect 3898 6496 3962 6500
rect 3978 6556 4042 6560
rect 3978 6500 3982 6556
rect 3982 6500 4038 6556
rect 4038 6500 4042 6556
rect 3978 6496 4042 6500
rect 4058 6556 4122 6560
rect 4058 6500 4062 6556
rect 4062 6500 4118 6556
rect 4118 6500 4122 6556
rect 4058 6496 4122 6500
rect 8818 6556 8882 6560
rect 8818 6500 8822 6556
rect 8822 6500 8878 6556
rect 8878 6500 8882 6556
rect 8818 6496 8882 6500
rect 8898 6556 8962 6560
rect 8898 6500 8902 6556
rect 8902 6500 8958 6556
rect 8958 6500 8962 6556
rect 8898 6496 8962 6500
rect 8978 6556 9042 6560
rect 8978 6500 8982 6556
rect 8982 6500 9038 6556
rect 9038 6500 9042 6556
rect 8978 6496 9042 6500
rect 9058 6556 9122 6560
rect 9058 6500 9062 6556
rect 9062 6500 9118 6556
rect 9118 6500 9122 6556
rect 9058 6496 9122 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 7568 6012 7632 6016
rect 7568 5956 7572 6012
rect 7572 5956 7628 6012
rect 7628 5956 7632 6012
rect 7568 5952 7632 5956
rect 7648 6012 7712 6016
rect 7648 5956 7652 6012
rect 7652 5956 7708 6012
rect 7708 5956 7712 6012
rect 7648 5952 7712 5956
rect 7728 6012 7792 6016
rect 7728 5956 7732 6012
rect 7732 5956 7788 6012
rect 7788 5956 7792 6012
rect 7728 5952 7792 5956
rect 7808 6012 7872 6016
rect 7808 5956 7812 6012
rect 7812 5956 7868 6012
rect 7868 5956 7872 6012
rect 7808 5952 7872 5956
rect 3818 5468 3882 5472
rect 3818 5412 3822 5468
rect 3822 5412 3878 5468
rect 3878 5412 3882 5468
rect 3818 5408 3882 5412
rect 3898 5468 3962 5472
rect 3898 5412 3902 5468
rect 3902 5412 3958 5468
rect 3958 5412 3962 5468
rect 3898 5408 3962 5412
rect 3978 5468 4042 5472
rect 3978 5412 3982 5468
rect 3982 5412 4038 5468
rect 4038 5412 4042 5468
rect 3978 5408 4042 5412
rect 4058 5468 4122 5472
rect 4058 5412 4062 5468
rect 4062 5412 4118 5468
rect 4118 5412 4122 5468
rect 4058 5408 4122 5412
rect 8818 5468 8882 5472
rect 8818 5412 8822 5468
rect 8822 5412 8878 5468
rect 8878 5412 8882 5468
rect 8818 5408 8882 5412
rect 8898 5468 8962 5472
rect 8898 5412 8902 5468
rect 8902 5412 8958 5468
rect 8958 5412 8962 5468
rect 8898 5408 8962 5412
rect 8978 5468 9042 5472
rect 8978 5412 8982 5468
rect 8982 5412 9038 5468
rect 9038 5412 9042 5468
rect 8978 5408 9042 5412
rect 9058 5468 9122 5472
rect 9058 5412 9062 5468
rect 9062 5412 9118 5468
rect 9118 5412 9122 5468
rect 9058 5408 9122 5412
rect 7568 4924 7632 4928
rect 7568 4868 7572 4924
rect 7572 4868 7628 4924
rect 7628 4868 7632 4924
rect 7568 4864 7632 4868
rect 7648 4924 7712 4928
rect 7648 4868 7652 4924
rect 7652 4868 7708 4924
rect 7708 4868 7712 4924
rect 7648 4864 7712 4868
rect 7728 4924 7792 4928
rect 7728 4868 7732 4924
rect 7732 4868 7788 4924
rect 7788 4868 7792 4924
rect 7728 4864 7792 4868
rect 7808 4924 7872 4928
rect 7808 4868 7812 4924
rect 7812 4868 7868 4924
rect 7868 4868 7872 4924
rect 7808 4864 7872 4868
rect 3818 4380 3882 4384
rect 3818 4324 3822 4380
rect 3822 4324 3878 4380
rect 3878 4324 3882 4380
rect 3818 4320 3882 4324
rect 3898 4380 3962 4384
rect 3898 4324 3902 4380
rect 3902 4324 3958 4380
rect 3958 4324 3962 4380
rect 3898 4320 3962 4324
rect 3978 4380 4042 4384
rect 3978 4324 3982 4380
rect 3982 4324 4038 4380
rect 4038 4324 4042 4380
rect 3978 4320 4042 4324
rect 4058 4380 4122 4384
rect 4058 4324 4062 4380
rect 4062 4324 4118 4380
rect 4118 4324 4122 4380
rect 4058 4320 4122 4324
rect 8818 4380 8882 4384
rect 8818 4324 8822 4380
rect 8822 4324 8878 4380
rect 8878 4324 8882 4380
rect 8818 4320 8882 4324
rect 8898 4380 8962 4384
rect 8898 4324 8902 4380
rect 8902 4324 8958 4380
rect 8958 4324 8962 4380
rect 8898 4320 8962 4324
rect 8978 4380 9042 4384
rect 8978 4324 8982 4380
rect 8982 4324 9038 4380
rect 9038 4324 9042 4380
rect 8978 4320 9042 4324
rect 9058 4380 9122 4384
rect 9058 4324 9062 4380
rect 9062 4324 9118 4380
rect 9118 4324 9122 4380
rect 9058 4320 9122 4324
rect 7568 3836 7632 3840
rect 7568 3780 7572 3836
rect 7572 3780 7628 3836
rect 7628 3780 7632 3836
rect 7568 3776 7632 3780
rect 7648 3836 7712 3840
rect 7648 3780 7652 3836
rect 7652 3780 7708 3836
rect 7708 3780 7712 3836
rect 7648 3776 7712 3780
rect 7728 3836 7792 3840
rect 7728 3780 7732 3836
rect 7732 3780 7788 3836
rect 7788 3780 7792 3836
rect 7728 3776 7792 3780
rect 7808 3836 7872 3840
rect 7808 3780 7812 3836
rect 7812 3780 7868 3836
rect 7868 3780 7872 3836
rect 7808 3776 7872 3780
rect 3818 3292 3882 3296
rect 3818 3236 3822 3292
rect 3822 3236 3878 3292
rect 3878 3236 3882 3292
rect 3818 3232 3882 3236
rect 3898 3292 3962 3296
rect 3898 3236 3902 3292
rect 3902 3236 3958 3292
rect 3958 3236 3962 3292
rect 3898 3232 3962 3236
rect 3978 3292 4042 3296
rect 3978 3236 3982 3292
rect 3982 3236 4038 3292
rect 4038 3236 4042 3292
rect 3978 3232 4042 3236
rect 4058 3292 4122 3296
rect 4058 3236 4062 3292
rect 4062 3236 4118 3292
rect 4118 3236 4122 3292
rect 4058 3232 4122 3236
rect 8818 3292 8882 3296
rect 8818 3236 8822 3292
rect 8822 3236 8878 3292
rect 8878 3236 8882 3292
rect 8818 3232 8882 3236
rect 8898 3292 8962 3296
rect 8898 3236 8902 3292
rect 8902 3236 8958 3292
rect 8958 3236 8962 3292
rect 8898 3232 8962 3236
rect 8978 3292 9042 3296
rect 8978 3236 8982 3292
rect 8982 3236 9038 3292
rect 9038 3236 9042 3292
rect 8978 3232 9042 3236
rect 9058 3292 9122 3296
rect 9058 3236 9062 3292
rect 9062 3236 9118 3292
rect 9118 3236 9122 3292
rect 9058 3232 9122 3236
rect 7568 2748 7632 2752
rect 7568 2692 7572 2748
rect 7572 2692 7628 2748
rect 7628 2692 7632 2748
rect 7568 2688 7632 2692
rect 7648 2748 7712 2752
rect 7648 2692 7652 2748
rect 7652 2692 7708 2748
rect 7708 2692 7712 2748
rect 7648 2688 7712 2692
rect 7728 2748 7792 2752
rect 7728 2692 7732 2748
rect 7732 2692 7788 2748
rect 7788 2692 7792 2748
rect 7728 2688 7792 2692
rect 7808 2748 7872 2752
rect 7808 2692 7812 2748
rect 7812 2692 7868 2748
rect 7868 2692 7872 2748
rect 7808 2688 7872 2692
rect 3818 2204 3882 2208
rect 3818 2148 3822 2204
rect 3822 2148 3878 2204
rect 3878 2148 3882 2204
rect 3818 2144 3882 2148
rect 3898 2204 3962 2208
rect 3898 2148 3902 2204
rect 3902 2148 3958 2204
rect 3958 2148 3962 2204
rect 3898 2144 3962 2148
rect 3978 2204 4042 2208
rect 3978 2148 3982 2204
rect 3982 2148 4038 2204
rect 4038 2148 4042 2204
rect 3978 2144 4042 2148
rect 4058 2204 4122 2208
rect 4058 2148 4062 2204
rect 4062 2148 4118 2204
rect 4118 2148 4122 2204
rect 4058 2144 4122 2148
rect 8818 2204 8882 2208
rect 8818 2148 8822 2204
rect 8822 2148 8878 2204
rect 8878 2148 8882 2204
rect 8818 2144 8882 2148
rect 8898 2204 8962 2208
rect 8898 2148 8902 2204
rect 8902 2148 8958 2204
rect 8958 2148 8962 2204
rect 8898 2144 8962 2148
rect 8978 2204 9042 2208
rect 8978 2148 8982 2204
rect 8982 2148 9038 2204
rect 9038 2148 9042 2204
rect 8978 2144 9042 2148
rect 9058 2204 9122 2208
rect 9058 2148 9062 2204
rect 9062 2148 9118 2204
rect 9118 2148 9122 2204
rect 9058 2144 9122 2148
rect 7568 1660 7632 1664
rect 7568 1604 7572 1660
rect 7572 1604 7628 1660
rect 7628 1604 7632 1660
rect 7568 1600 7632 1604
rect 7648 1660 7712 1664
rect 7648 1604 7652 1660
rect 7652 1604 7708 1660
rect 7708 1604 7712 1660
rect 7648 1600 7712 1604
rect 7728 1660 7792 1664
rect 7728 1604 7732 1660
rect 7732 1604 7788 1660
rect 7788 1604 7792 1660
rect 7728 1600 7792 1604
rect 7808 1660 7872 1664
rect 7808 1604 7812 1660
rect 7812 1604 7868 1660
rect 7868 1604 7872 1660
rect 7808 1600 7872 1604
rect 3818 1116 3882 1120
rect 3818 1060 3822 1116
rect 3822 1060 3878 1116
rect 3878 1060 3882 1116
rect 3818 1056 3882 1060
rect 3898 1116 3962 1120
rect 3898 1060 3902 1116
rect 3902 1060 3958 1116
rect 3958 1060 3962 1116
rect 3898 1056 3962 1060
rect 3978 1116 4042 1120
rect 3978 1060 3982 1116
rect 3982 1060 4038 1116
rect 4038 1060 4042 1116
rect 3978 1056 4042 1060
rect 4058 1116 4122 1120
rect 4058 1060 4062 1116
rect 4062 1060 4118 1116
rect 4118 1060 4122 1116
rect 4058 1056 4122 1060
rect 8818 1116 8882 1120
rect 8818 1060 8822 1116
rect 8822 1060 8878 1116
rect 8878 1060 8882 1116
rect 8818 1056 8882 1060
rect 8898 1116 8962 1120
rect 8898 1060 8902 1116
rect 8902 1060 8958 1116
rect 8958 1060 8962 1116
rect 8898 1056 8962 1060
rect 8978 1116 9042 1120
rect 8978 1060 8982 1116
rect 8982 1060 9038 1116
rect 9038 1060 9042 1116
rect 8978 1056 9042 1060
rect 9058 1116 9122 1120
rect 9058 1060 9062 1116
rect 9062 1060 9118 1116
rect 9118 1060 9122 1116
rect 9058 1056 9122 1060
<< metal4 >>
rect 2560 11456 2880 11472
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8266 2880 9216
rect 2560 8192 2602 8266
rect 2838 8192 2880 8266
rect 2560 8128 2568 8192
rect 2872 8128 2880 8192
rect 2560 8030 2602 8128
rect 2838 8030 2880 8128
rect 2560 7104 2880 8030
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5280 2880 5952
rect 3810 10912 4130 11472
rect 3810 10848 3818 10912
rect 3882 10848 3898 10912
rect 3962 10848 3978 10912
rect 4042 10848 4058 10912
rect 4122 10848 4130 10912
rect 3810 9824 4130 10848
rect 3810 9760 3818 9824
rect 3882 9760 3898 9824
rect 3962 9760 3978 9824
rect 4042 9760 4058 9824
rect 4122 9760 4130 9824
rect 3810 9111 4130 9760
rect 3810 8875 3852 9111
rect 4088 8875 4130 9111
rect 3810 8736 4130 8875
rect 3810 8672 3818 8736
rect 3882 8672 3898 8736
rect 3962 8672 3978 8736
rect 4042 8672 4058 8736
rect 4122 8672 4130 8736
rect 3810 7648 4130 8672
rect 3810 7584 3818 7648
rect 3882 7584 3898 7648
rect 3962 7584 3978 7648
rect 4042 7584 4058 7648
rect 4122 7584 4130 7648
rect 3810 6560 4130 7584
rect 3810 6496 3818 6560
rect 3882 6496 3898 6560
rect 3962 6496 3978 6560
rect 4042 6496 4058 6560
rect 4122 6496 4130 6560
rect 3810 5731 4130 6496
rect 3810 5495 3852 5731
rect 4088 5495 4130 5731
rect 3810 5472 4130 5495
rect 3810 5408 3818 5472
rect 3882 5408 3898 5472
rect 3962 5408 3978 5472
rect 4042 5408 4058 5472
rect 4122 5408 4130 5472
rect 3810 4384 4130 5408
rect 3810 4320 3818 4384
rect 3882 4320 3898 4384
rect 3962 4320 3978 4384
rect 4042 4320 4058 4384
rect 4122 4320 4130 4384
rect 1996 4041 2276 4083
rect 1996 3805 2018 4041
rect 2254 3805 2276 4041
rect 1996 3763 2276 3805
rect 3810 3296 4130 4320
rect 1256 3196 1536 3238
rect 1256 2960 1278 3196
rect 1514 2960 1536 3196
rect 1256 2918 1536 2960
rect 3810 3232 3818 3296
rect 3882 3232 3898 3296
rect 3962 3232 3978 3296
rect 4042 3232 4058 3296
rect 4122 3232 4130 3296
rect 3810 2351 4130 3232
rect 3810 2208 3852 2351
rect 4088 2208 4130 2351
rect 3810 2144 3818 2208
rect 4122 2144 4130 2208
rect 3810 2115 3852 2144
rect 4088 2115 4130 2144
rect 3810 1120 4130 2115
rect 3810 1056 3818 1120
rect 3882 1056 3898 1120
rect 3962 1056 3978 1120
rect 4042 1056 4058 1120
rect 4122 1056 4130 1120
rect 3810 1040 4130 1056
rect 5060 3196 5380 11472
rect 5060 2960 5102 3196
rect 5338 2960 5380 3196
rect 5060 1040 5380 2960
rect 6310 4041 6630 11472
rect 6310 3805 6352 4041
rect 6588 3805 6630 4041
rect 6310 1040 6630 3805
rect 7560 11456 7880 11472
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 7560 10368 7880 11392
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 9280 7880 10304
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 8266 7880 9216
rect 7560 8192 7602 8266
rect 7838 8192 7880 8266
rect 7560 8128 7568 8192
rect 7872 8128 7880 8192
rect 7560 8030 7602 8128
rect 7838 8030 7880 8128
rect 7560 7104 7880 8030
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 6016 7880 7040
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 4928 7880 5952
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 7560 3840 7880 4864
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 2752 7880 3776
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 1664 7880 2688
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 7560 1506 7880 1600
rect 7560 1270 7602 1506
rect 7838 1270 7880 1506
rect 7560 1040 7880 1270
rect 8810 10912 9130 11472
rect 8810 10848 8818 10912
rect 8882 10848 8898 10912
rect 8962 10848 8978 10912
rect 9042 10848 9058 10912
rect 9122 10848 9130 10912
rect 8810 9824 9130 10848
rect 8810 9760 8818 9824
rect 8882 9760 8898 9824
rect 8962 9760 8978 9824
rect 9042 9760 9058 9824
rect 9122 9760 9130 9824
rect 8810 9111 9130 9760
rect 8810 8875 8852 9111
rect 9088 8875 9130 9111
rect 8810 8736 9130 8875
rect 8810 8672 8818 8736
rect 8882 8672 8898 8736
rect 8962 8672 8978 8736
rect 9042 8672 9058 8736
rect 9122 8672 9130 8736
rect 8810 7648 9130 8672
rect 8810 7584 8818 7648
rect 8882 7584 8898 7648
rect 8962 7584 8978 7648
rect 9042 7584 9058 7648
rect 9122 7584 9130 7648
rect 8810 6560 9130 7584
rect 8810 6496 8818 6560
rect 8882 6496 8898 6560
rect 8962 6496 8978 6560
rect 9042 6496 9058 6560
rect 9122 6496 9130 6560
rect 8810 5731 9130 6496
rect 8810 5495 8852 5731
rect 9088 5495 9130 5731
rect 8810 5472 9130 5495
rect 8810 5408 8818 5472
rect 8882 5408 8898 5472
rect 8962 5408 8978 5472
rect 9042 5408 9058 5472
rect 9122 5408 9130 5472
rect 8810 4384 9130 5408
rect 8810 4320 8818 4384
rect 8882 4320 8898 4384
rect 8962 4320 8978 4384
rect 9042 4320 9058 4384
rect 9122 4320 9130 4384
rect 8810 3296 9130 4320
rect 8810 3232 8818 3296
rect 8882 3232 8898 3296
rect 8962 3232 8978 3296
rect 9042 3232 9058 3296
rect 9122 3232 9130 3296
rect 8810 2351 9130 3232
rect 8810 2208 8852 2351
rect 9088 2208 9130 2351
rect 8810 2144 8818 2208
rect 9122 2144 9130 2208
rect 8810 2115 8852 2144
rect 9088 2115 9130 2144
rect 8810 1120 9130 2115
rect 8810 1056 8818 1120
rect 8882 1056 8898 1120
rect 8962 1056 8978 1120
rect 9042 1056 9058 1120
rect 9122 1056 9130 1120
rect 8810 1040 9130 1056
<< obsm4 >>
rect 13400 0 34000 13000
<< via4 >>
rect 2602 8192 2838 8266
rect 2602 8128 2632 8192
rect 2632 8128 2648 8192
rect 2648 8128 2712 8192
rect 2712 8128 2728 8192
rect 2728 8128 2792 8192
rect 2792 8128 2808 8192
rect 2808 8128 2838 8192
rect 2602 8030 2838 8128
rect 3852 8875 4088 9111
rect 3852 5495 4088 5731
rect 2018 3805 2254 4041
rect 1278 2960 1514 3196
rect 3852 2208 4088 2351
rect 3852 2144 3882 2208
rect 3882 2144 3898 2208
rect 3898 2144 3962 2208
rect 3962 2144 3978 2208
rect 3978 2144 4042 2208
rect 4042 2144 4058 2208
rect 4058 2144 4088 2208
rect 3852 2115 4088 2144
rect 5102 2960 5338 3196
rect 6352 3805 6588 4041
rect 7602 8192 7838 8266
rect 7602 8128 7632 8192
rect 7632 8128 7648 8192
rect 7648 8128 7712 8192
rect 7712 8128 7728 8192
rect 7728 8128 7792 8192
rect 7792 8128 7808 8192
rect 7808 8128 7838 8192
rect 7602 8030 7838 8128
rect 7602 1270 7838 1506
rect 8852 8875 9088 9111
rect 8852 5495 9088 5731
rect 8852 2208 9088 2351
rect 8852 2144 8882 2208
rect 8882 2144 8898 2208
rect 8898 2144 8962 2208
rect 8962 2144 8978 2208
rect 8978 2144 9042 2208
rect 9042 2144 9058 2208
rect 9058 2144 9088 2208
rect 8852 2115 9088 2144
<< metal5 >>
rect 872 9111 9892 9153
rect 872 8875 3852 9111
rect 4088 8875 8852 9111
rect 9088 8875 9892 9111
rect 872 8833 9892 8875
rect 872 8266 9892 8308
rect 872 8030 2602 8266
rect 2838 8030 7602 8266
rect 7838 8030 9892 8266
rect 872 7988 9892 8030
rect 872 5731 9892 5773
rect 872 5495 3852 5731
rect 4088 5495 8852 5731
rect 9088 5495 9892 5731
rect 872 5453 9892 5495
rect 872 4041 9892 4083
rect 872 3805 2018 4041
rect 2254 3805 6352 4041
rect 6588 3805 9892 4041
rect 872 3763 9892 3805
rect 872 3196 9892 3238
rect 872 2960 1278 3196
rect 1514 2960 5102 3196
rect 5338 2960 9892 3196
rect 872 2918 9892 2960
rect 872 2351 9892 2393
rect 872 2115 3852 2351
rect 4088 2115 8852 2351
rect 9088 2115 9892 2351
rect 872 2073 9892 2115
rect 872 1506 9892 1548
rect 872 1270 7602 1506
rect 7838 1270 9892 1506
rect 872 1228 9892 1270
<< obsm5 >>
rect 13400 0 34000 13000
use sky130_fd_sc_hd__diode_2  ANTENNA__058__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 9568 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A_N
timestamp 1659098407
transform -1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__B
timestamp 1659098407
transform 1 0 9384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A2
timestamp 1659098407
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A_N
timestamp 1659098407
transform -1 0 8924 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__C
timestamp 1659098407
transform -1 0 9568 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A0
timestamp 1659098407
transform -1 0 9384 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A0
timestamp 1659098407
transform -1 0 9568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1659098407
transform -1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__B
timestamp 1659098407
transform 1 0 6624 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A_N
timestamp 1659098407
transform -1 0 6992 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__B
timestamp 1659098407
transform 1 0 6164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1659098407
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__B
timestamp 1659098407
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A_N
timestamp 1659098407
transform 1 0 5244 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__B
timestamp 1659098407
transform 1 0 4600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1659098407
transform 1 0 9016 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__B
timestamp 1659098407
transform -1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A_N
timestamp 1659098407
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__B
timestamp 1659098407
transform -1 0 2760 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1659098407
transform 1 0 9384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__B
timestamp 1659098407
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A_N
timestamp 1659098407
transform 1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__B
timestamp 1659098407
transform -1 0 9568 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1659098407
transform 1 0 3588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__B
timestamp 1659098407
transform 1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A_N
timestamp 1659098407
transform 1 0 4232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__B
timestamp 1659098407
transform 1 0 2668 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1659098407
transform -1 0 1564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__B
timestamp 1659098407
transform -1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A_N
timestamp 1659098407
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__B
timestamp 1659098407
transform 1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1659098407
transform -1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__B
timestamp 1659098407
transform 1 0 5152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A_N
timestamp 1659098407
transform -1 0 4968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__B
timestamp 1659098407
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1659098407
transform 1 0 8556 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__B
timestamp 1659098407
transform -1 0 8096 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A_N
timestamp 1659098407
transform 1 0 8280 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__B
timestamp 1659098407
transform -1 0 7452 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1659098407
transform 1 0 8280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__B
timestamp 1659098407
transform -1 0 8648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A_N
timestamp 1659098407
transform 1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__B
timestamp 1659098407
transform -1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1659098407
transform -1 0 8464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__B
timestamp 1659098407
transform -1 0 9384 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A_N
timestamp 1659098407
transform -1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B
timestamp 1659098407
transform 1 0 8004 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1659098407
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__B
timestamp 1659098407
transform -1 0 5520 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A_N
timestamp 1659098407
transform -1 0 5336 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__B
timestamp 1659098407
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1659098407
transform 1 0 5428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__B
timestamp 1659098407
transform -1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A_N
timestamp 1659098407
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__B
timestamp 1659098407
transform -1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1659098407
transform 1 0 7176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__B
timestamp 1659098407
transform -1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A_N
timestamp 1659098407
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__B
timestamp 1659098407
transform -1 0 6072 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__D
timestamp 1659098407
transform -1 0 8556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__RESET_B
timestamp 1659098407
transform 1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__RESET_B
timestamp 1659098407
transform -1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__RESET_B
timestamp 1659098407
transform -1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__RESET_B
timestamp 1659098407
transform 1 0 2852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__RESET_B
timestamp 1659098407
transform 1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__RESET_B
timestamp 1659098407
transform 1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__RESET_B
timestamp 1659098407
transform 1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__RESET_B
timestamp 1659098407
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__RESET_B
timestamp 1659098407
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__RESET_B
timestamp 1659098407
transform 1 0 9384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__RESET_B
timestamp 1659098407
transform 1 0 8004 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__RESET_B
timestamp 1659098407
transform 1 0 9200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__RESET_B
timestamp 1659098407
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__RESET_B
timestamp 1659098407
transform -1 0 7728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1659098407
transform -1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1659098407
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1659098407
transform -1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_load_A
timestamp 1659098407
transform -1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 5520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_52 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 5704 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_64
timestamp 1659098407
transform 1 0 6808 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 7912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_80
timestamp 1659098407
transform 1 0 8280 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1659098407
transform 1 0 6072 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_68
timestamp 1659098407
transform 1 0 7176 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 7452 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 1659098407
transform 1 0 7820 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1659098407
transform 1 0 8096 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_82
timestamp 1659098407
transform 1 0 8464 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_40
timestamp 1659098407
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 1659098407
transform 1 0 4968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_70
timestamp 1659098407
transform 1 0 7360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1659098407
transform 1 0 8556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_39
timestamp 1659098407
transform 1 0 4508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_93
timestamp 1659098407
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_50
timestamp 1659098407
transform 1 0 5520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_60
timestamp 1659098407
transform 1 0 6440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_76
timestamp 1659098407
transform 1 0 7912 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_93
timestamp 1659098407
transform 1 0 9476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 1196 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1659098407
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 1196 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1659098407
transform 1 0 1196 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1659098407
transform 1 0 3404 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_44
timestamp 1659098407
transform 1 0 4968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_76
timestamp 1659098407
transform 1 0 7912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1659098407
transform 1 0 1196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1659098407
transform 1 0 2300 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_48
timestamp 1659098407
transform 1 0 5336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1659098407
transform 1 0 1196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1659098407
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1659098407
transform 1 0 1196 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_35
timestamp 1659098407
transform 1 0 4140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1659098407
transform 1 0 1196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_38
timestamp 1659098407
transform 1 0 4416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1659098407
transform 1 0 8556 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1659098407
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1659098407
transform 1 0 1196 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_65
timestamp 1659098407
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1659098407
transform 1 0 1196 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1659098407
transform 1 0 1196 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1659098407
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_72
timestamp 1659098407
transform 1 0 7544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1659098407
transform 1 0 1196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 2300 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_24
timestamp 1659098407
transform 1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1659098407
transform 1 0 4968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_48
timestamp 1659098407
transform 1 0 5336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_52
timestamp 1659098407
transform 1 0 5704 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_61
timestamp 1659098407
transform 1 0 6532 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_66
timestamp 1659098407
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_71
timestamp 1659098407
transform 1 0 7452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_79
timestamp 1659098407
transform 1 0 8188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1659098407
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1659098407
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1659098407
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1659098407
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1659098407
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1659098407
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1659098407
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1659098407
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1659098407
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1659098407
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1659098407
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1659098407
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1659098407
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1659098407
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1659098407
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1659098407
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1659098407
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1659098407
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1659098407
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1659098407
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1659098407
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1659098407
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1659098407
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1659098407
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1659098407
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1659098407
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1659098407
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1659098407
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1659098407
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1659098407
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1659098407
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1659098407
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1659098407
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1659098407
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1659098407
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1659098407
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1659098407
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1659098407
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1659098407
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1659098407
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1659098407
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1659098407
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1659098407
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1659098407
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1659098407
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1659098407
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1659098407
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1659098407
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1659098407
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1659098407
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1659098407
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1659098407
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1659098407
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1659098407
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1659098407
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1659098407
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1659098407
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1659098407
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1659098407
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1659098407
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1659098407
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1659098407
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1659098407
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1659098407
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1659098407
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1659098407
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _058_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059__1
timestamp 1659098407
transform -1 0 6072 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _060__14
timestamp 1659098407
transform -1 0 8004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 8004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 9384 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 9384 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 8648 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 9476 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _066_
timestamp 1659098407
transform -1 0 9568 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 6808 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _068_
timestamp 1659098407
transform 1 0 6164 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _069_
timestamp 1659098407
transform 1 0 3036 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _070_
timestamp 1659098407
transform -1 0 5244 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _071_
timestamp 1659098407
transform -1 0 8740 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _072_
timestamp 1659098407
transform 1 0 5428 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _073_
timestamp 1659098407
transform -1 0 9200 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _074_
timestamp 1659098407
transform -1 0 9384 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _075_
timestamp 1659098407
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _076_
timestamp 1659098407
transform -1 0 4232 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _077_
timestamp 1659098407
transform 1 0 3680 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _078_
timestamp 1659098407
transform -1 0 4968 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _079_
timestamp 1659098407
transform 1 0 5336 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _080_
timestamp 1659098407
transform 1 0 3956 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _081_
timestamp 1659098407
transform 1 0 8096 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _082_
timestamp 1659098407
transform 1 0 7452 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _083_
timestamp 1659098407
transform 1 0 9016 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _084_
timestamp 1659098407
transform 1 0 7176 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _085_
timestamp 1659098407
transform -1 0 9200 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _086_
timestamp 1659098407
transform -1 0 8648 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _087_
timestamp 1659098407
transform 1 0 4140 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _088_
timestamp 1659098407
transform 1 0 3496 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _089_
timestamp 1659098407
transform 1 0 5152 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _090_
timestamp 1659098407
transform -1 0 6348 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _091_
timestamp 1659098407
transform -1 0 6808 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _092_
timestamp 1659098407
transform -1 0 6348 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _093__2
timestamp 1659098407
transform -1 0 3128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _094__3
timestamp 1659098407
transform -1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095__4
timestamp 1659098407
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096__5
timestamp 1659098407
transform -1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097__6
timestamp 1659098407
transform -1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098__7
timestamp 1659098407
transform -1 0 4600 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099__8
timestamp 1659098407
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100__9
timestamp 1659098407
transform 1 0 6256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101__10
timestamp 1659098407
transform -1 0 7544 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102__11
timestamp 1659098407
transform -1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103__12
timestamp 1659098407
transform -1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104__13
timestamp 1659098407
transform -1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_2  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 5428 0 1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _106_
timestamp 1659098407
transform 1 0 2760 0 -1 10880
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _107_
timestamp 1659098407
transform 1 0 5060 0 1 6528
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _108_
timestamp 1659098407
transform 1 0 6072 0 1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _109_
timestamp 1659098407
transform 1 0 2760 0 -1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _110_
timestamp 1659098407
transform 1 0 2760 0 -1 6528
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _111_
timestamp 1659098407
transform 1 0 3312 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _112_
timestamp 1659098407
transform 1 0 6808 0 1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _113_
timestamp 1659098407
transform 1 0 6532 0 1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _114_
timestamp 1659098407
transform 1 0 6992 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _115_
timestamp 1659098407
transform 1 0 3312 0 -1 2176
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _116_
timestamp 1659098407
transform 1 0 3496 0 -1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _117_
timestamp 1659098407
transform 1 0 4600 0 -1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_2  _118_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 6440 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _119_
timestamp 1659098407
transform 1 0 1564 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _120_
timestamp 1659098407
transform -1 0 3312 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _121_
timestamp 1659098407
transform 1 0 1472 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _122_
timestamp 1659098407
transform 1 0 1472 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _123_
timestamp 1659098407
transform 1 0 1564 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _124_
timestamp 1659098407
transform 1 0 3312 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _125_
timestamp 1659098407
transform 1 0 3312 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _126_
timestamp 1659098407
transform 1 0 4140 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _127_
timestamp 1659098407
transform 1 0 6164 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _128_
timestamp 1659098407
transform 1 0 6164 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _129_
timestamp 1659098407
transform 1 0 5980 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _130_
timestamp 1659098407
transform 1 0 6440 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _131_
timestamp 1659098407
transform 1 0 7636 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 9200 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1659098407
transform 1 0 8832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1659098407
transform 1 0 8832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _135_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 8740 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 6072 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 1659098407
transform -1 0 8004 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_clock
timestamp 1659098407
transform -1 0 5152 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_load
timestamp 1659098407
transform -1 0 5152 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_clock
timestamp 1659098407
transform 1 0 6164 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_load
timestamp 1659098407
transform -1 0 6072 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 9200 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform 1 0 6532 0 -1 4352
box -38 -48 1694 592
use gpio_logic_high  gpio_logic_high
timestamp 0
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659098407
transform -1 0 8740 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1659098407
transform -1 0 8740 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1659098407
transform 1 0 2024 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1659098407
transform -1 0 4140 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1659098407
transform -1 0 4324 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1659098407
transform -1 0 6900 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1659098407
transform -1 0 6072 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1659098407
transform -1 0 9016 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1659098407
transform -1 0 4324 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1659098407
transform -1 0 5980 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1659098407
transform -1 0 6440 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1659098407
transform 1 0 3496 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1659098407
transform -1 0 9016 0 -1 5440
box -38 -48 774 592
<< labels >>
flabel metal2 s 938 12200 994 13000 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 0 nsew signal input
flabel metal2 s 5538 12200 5594 13000 0 FreeSans 224 90 0 0 gpio_defaults[10]
port 1 nsew signal input
flabel metal2 s 5998 12200 6054 13000 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 2 nsew signal input
flabel metal2 s 6458 12200 6514 13000 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 3 nsew signal input
flabel metal2 s 1398 12200 1454 13000 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 4 nsew signal input
flabel metal2 s 1858 12200 1914 13000 0 FreeSans 224 90 0 0 gpio_defaults[2]
port 5 nsew signal input
flabel metal2 s 2318 12200 2374 13000 0 FreeSans 224 90 0 0 gpio_defaults[3]
port 6 nsew signal input
flabel metal2 s 2778 12200 2834 13000 0 FreeSans 224 90 0 0 gpio_defaults[4]
port 7 nsew signal input
flabel metal2 s 3238 12200 3294 13000 0 FreeSans 224 90 0 0 gpio_defaults[5]
port 8 nsew signal input
flabel metal2 s 3698 12200 3754 13000 0 FreeSans 224 90 0 0 gpio_defaults[6]
port 9 nsew signal input
flabel metal2 s 4158 12200 4214 13000 0 FreeSans 224 90 0 0 gpio_defaults[7]
port 10 nsew signal input
flabel metal2 s 4618 12200 4674 13000 0 FreeSans 224 90 0 0 gpio_defaults[8]
port 11 nsew signal input
flabel metal2 s 5078 12200 5134 13000 0 FreeSans 224 90 0 0 gpio_defaults[9]
port 12 nsew signal input
flabel metal3 s 14000 824 34000 944 0 FreeSans 480 0 0 0 mgmt_gpio_in
port 13 nsew signal tristate
flabel metal3 s 14000 1640 34000 1760 0 FreeSans 480 0 0 0 mgmt_gpio_oeb
port 14 nsew signal input
flabel metal3 s 14000 2048 34000 2168 0 FreeSans 480 0 0 0 mgmt_gpio_out
port 15 nsew signal input
flabel metal3 s 14000 1232 34000 1352 0 FreeSans 480 0 0 0 one
port 16 nsew signal tristate
flabel metal3 s 14000 2456 34000 2576 0 FreeSans 480 0 0 0 pad_gpio_ana_en
port 17 nsew signal tristate
flabel metal3 s 14000 2864 34000 2984 0 FreeSans 480 0 0 0 pad_gpio_ana_pol
port 18 nsew signal tristate
flabel metal3 s 14000 3272 34000 3392 0 FreeSans 480 0 0 0 pad_gpio_ana_sel
port 19 nsew signal tristate
flabel metal3 s 14000 3680 34000 3800 0 FreeSans 480 0 0 0 pad_gpio_dm[0]
port 20 nsew signal tristate
flabel metal3 s 14000 4088 34000 4208 0 FreeSans 480 0 0 0 pad_gpio_dm[1]
port 21 nsew signal tristate
flabel metal3 s 14000 4496 34000 4616 0 FreeSans 480 0 0 0 pad_gpio_dm[2]
port 22 nsew signal tristate
flabel metal3 s 14000 4904 34000 5024 0 FreeSans 480 0 0 0 pad_gpio_holdover
port 23 nsew signal tristate
flabel metal3 s 14000 5312 34000 5432 0 FreeSans 480 0 0 0 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
flabel metal3 s 14000 5720 34000 5840 0 FreeSans 480 0 0 0 pad_gpio_in
port 25 nsew signal input
flabel metal3 s 14000 6128 34000 6248 0 FreeSans 480 0 0 0 pad_gpio_inenb
port 26 nsew signal tristate
flabel metal3 s 14000 6536 34000 6656 0 FreeSans 480 0 0 0 pad_gpio_out
port 27 nsew signal tristate
flabel metal3 s 14000 6944 34000 7064 0 FreeSans 480 0 0 0 pad_gpio_outenb
port 28 nsew signal tristate
flabel metal3 s 14000 7352 34000 7472 0 FreeSans 480 0 0 0 pad_gpio_slow_sel
port 29 nsew signal tristate
flabel metal3 s 14000 7760 34000 7880 0 FreeSans 480 0 0 0 pad_gpio_vtrip_sel
port 30 nsew signal tristate
flabel metal3 s 14000 8168 34000 8288 0 FreeSans 480 0 0 0 resetn
port 31 nsew signal input
flabel metal3 s 14000 8576 34000 8696 0 FreeSans 480 0 0 0 resetn_out
port 32 nsew signal tristate
flabel metal3 s 14000 8984 34000 9104 0 FreeSans 480 0 0 0 serial_clock
port 33 nsew signal input
flabel metal3 s 14000 9392 34000 9512 0 FreeSans 480 0 0 0 serial_clock_out
port 34 nsew signal tristate
flabel metal3 s 14000 9800 34000 9920 0 FreeSans 480 0 0 0 serial_data_in
port 35 nsew signal input
flabel metal3 s 14000 10208 34000 10328 0 FreeSans 480 0 0 0 serial_data_out
port 36 nsew signal tristate
flabel metal3 s 14000 10616 34000 10736 0 FreeSans 480 0 0 0 serial_load
port 37 nsew signal input
flabel metal3 s 14000 11024 34000 11144 0 FreeSans 480 0 0 0 serial_load_out
port 38 nsew signal tristate
flabel metal3 s 14000 11432 34000 11552 0 FreeSans 480 0 0 0 user_gpio_in
port 39 nsew signal tristate
flabel metal3 s 14000 11840 34000 11960 0 FreeSans 480 0 0 0 user_gpio_oeb
port 40 nsew signal input
flabel metal3 s 14000 12248 34000 12368 0 FreeSans 480 0 0 0 user_gpio_out
port 41 nsew signal input
flabel metal4 s 2560 5280 2880 11472 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 7560 1040 7880 11472 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 1228 9892 1548 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 7988 9892 8308 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 5060 1040 5380 11472 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 2918 9892 3238 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 3810 1040 4130 11472 0 FreeSans 1920 90 0 0 vssd
port 44 nsew ground bidirectional
flabel metal4 s 8810 1040 9130 11472 0 FreeSans 1920 90 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 2073 9892 2393 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 5453 9892 5773 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 8833 9892 9153 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal4 s 6310 1040 6630 11472 0 FreeSans 1920 90 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 3763 9892 4083 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal3 s 14000 416 34000 536 0 FreeSans 480 0 0 0 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
