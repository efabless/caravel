module caravan_power_routing ();
endmodule
