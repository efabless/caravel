* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_1 abstract view
.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb sram_ro_addr[0] sram_ro_addr[1] sram_ro_addr[2]
+ sram_ro_addr[3] sram_ro_addr[4] sram_ro_addr[5] sram_ro_addr[6] sram_ro_addr[7]
+ sram_ro_clk sram_ro_csb sram_ro_data[0] sram_ro_data[10] sram_ro_data[11] sram_ro_data[12]
+ sram_ro_data[13] sram_ro_data[14] sram_ro_data[15] sram_ro_data[16] sram_ro_data[17]
+ sram_ro_data[18] sram_ro_data[19] sram_ro_data[1] sram_ro_data[20] sram_ro_data[21]
+ sram_ro_data[22] sram_ro_data[23] sram_ro_data[24] sram_ro_data[25] sram_ro_data[26]
+ sram_ro_data[27] sram_ro_data[28] sram_ro_data[29] sram_ro_data[2] sram_ro_data[30]
+ sram_ro_data[31] sram_ro_data[3] sram_ro_data[4] sram_ro_data[5] sram_ro_data[6]
+ sram_ro_data[7] sram_ro_data[8] sram_ro_data[9] trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_100_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7963_ _8505_/A _7963_/B VGND VGND VPWR VPWR _7964_/B sky130_fd_sc_hd__or2_1
X_9702_ _9705_/CLK _9702_/D _6177_/A VGND VGND VPWR VPWR _9702_/Q sky130_fd_sc_hd__dfrtp_1
X_6914_ _9228_/Q VGND VGND VPWR VPWR _6914_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7894_ _8118_/A _8312_/B VGND VGND VPWR VPWR _8641_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9633_ _9651_/CLK _9633_/D _9563_/SET_B VGND VGND VPWR VPWR _9633_/Q sky130_fd_sc_hd__dfrtp_1
X_6845_ _9762_/Q VGND VGND VPWR VPWR _6845_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9564_ _9569_/CLK _9564_/D _9563_/SET_B VGND VGND VPWR VPWR _9564_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6776_ _9685_/Q VGND VGND VPWR VPWR _6776_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9495_ _9569_/CLK hold45/X _9563_/SET_B VGND VGND VPWR VPWR _9495_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8515_ _8513_/Y _8514_/Y _8102_/A _8750_/C VGND VGND VPWR VPWR _8516_/B sky130_fd_sc_hd__a31o_1
X_5727_ _5727_/A VGND VGND VPWR VPWR _5727_/X sky130_fd_sc_hd__buf_4
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8446_ _8707_/B _8613_/A VGND VGND VPWR VPWR _8447_/A sky130_fd_sc_hd__or2_1
XFILLER_190_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5658_ _5698_/A _5658_/B VGND VGND VPWR VPWR _5658_/X sky130_fd_sc_hd__or2_1
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8377_ _8377_/A _8376_/X VGND VGND VPWR VPWR _8378_/B sky130_fd_sc_hd__or2b_1
X_4609_ _4689_/A _4750_/D _4689_/C _4750_/B VGND VGND VPWR VPWR _4818_/B sky130_fd_sc_hd__or4_4
X_5589_ _5698_/A _5589_/B VGND VGND VPWR VPWR _5590_/A sky130_fd_sc_hd__or2_1
Xhold340 hold340/A VGND VGND VPWR VPWR hold341/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold351 _4536_/X VGND VGND VPWR VPWR _4537_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold362 hold362/A VGND VGND VPWR VPWR _4643_/A sky130_fd_sc_hd__clkbuf_2
X_7328_ _4770_/Y _7155_/X _4912_/Y _7156_/X _7327_/X VGND VGND VPWR VPWR _7331_/C
+ sky130_fd_sc_hd__o221a_1
Xhold373 hold373/A VGND VGND VPWR VPWR _9641_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7259_ _6271_/Y _7151_/X _6302_/Y _7152_/X VGND VGND VPWR VPWR _7259_/X sky130_fd_sc_hd__o22a_1
XFILLER_131_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold384 hold384/A VGND VGND VPWR VPWR hold385/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 hold395/A VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_89_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4960_ _4969_/A VGND VGND VPWR VPWR _4961_/A sky130_fd_sc_hd__clkbuf_1
X_4891_ input4/X VGND VGND VPWR VPWR _4891_/Y sky130_fd_sc_hd__inv_2
X_6630_ _9771_/Q VGND VGND VPWR VPWR _6630_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6561_ _6559_/Y _5927_/B _6560_/Y _5047_/B VGND VGND VPWR VPWR _6561_/X sky130_fd_sc_hd__o22a_1
XFILLER_118_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8300_ _8552_/A _8304_/B VGND VGND VPWR VPWR _8409_/B sky130_fd_sc_hd__nor2_1
X_5512_ _9427_/Q _5507_/A _6008_/B1 _5507_/Y VGND VGND VPWR VPWR _9427_/D sky130_fd_sc_hd__a22o_1
X_6492_ _9384_/Q VGND VGND VPWR VPWR _6492_/Y sky130_fd_sc_hd__inv_2
X_9280_ _9420_/CLK _9280_/D _9537_/SET_B VGND VGND VPWR VPWR _9280_/Q sky130_fd_sc_hd__dfrtp_1
X_8231_ _8230_/A _8255_/A _8230_/Y VGND VGND VPWR VPWR _8387_/A sky130_fd_sc_hd__a21oi_1
XFILLER_145_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5443_ _9474_/Q _5437_/X _6008_/B1 _5438_/Y VGND VGND VPWR VPWR _5443_/X sky130_fd_sc_hd__a22o_1
X_5374_ _9521_/Q _5369_/A hold42/X _5369_/Y VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__a22o_1
X_8162_ _8439_/A _8439_/B _8139_/A VGND VGND VPWR VPWR _8162_/Y sky130_fd_sc_hd__o21ai_2
X_7113_ _7113_/A _7129_/B _7129_/C VGND VGND VPWR VPWR _7162_/A sky130_fd_sc_hd__or3_4
X_8093_ _8563_/A _8209_/A VGND VGND VPWR VPWR _8434_/A sky130_fd_sc_hd__or2_1
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7044_ _7044_/A VGND VGND VPWR VPWR _7045_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_101_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8995_ _9755_/Q _6660_/Y _8999_/S VGND VGND VPWR VPWR _8995_/X sky130_fd_sc_hd__mux2_1
X_7946_ _7903_/X _8272_/A _7926_/Y _7932_/X _7945_/X VGND VGND VPWR VPWR _7946_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7877_ _8140_/A VGND VGND VPWR VPWR _8236_/A sky130_fd_sc_hd__buf_4
X_9616_ _9731_/CLK _9616_/D _9731_/SET_B VGND VGND VPWR VPWR _9616_/Q sky130_fd_sc_hd__dfrtp_1
X_6828_ _6826_/Y _4558_/B _6827_/Y _4585_/B VGND VGND VPWR VPWR _6828_/X sky130_fd_sc_hd__o22a_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9547_ _9550_/CLK _9547_/D _9563_/SET_B VGND VGND VPWR VPWR _9547_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6759_ _6754_/Y _5428_/B _6755_/Y _5521_/B _6758_/X VGND VGND VPWR VPWR _6772_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9478_ _9483_/CLK _9478_/D _9727_/SET_B VGND VGND VPWR VPWR _9478_/Q sky130_fd_sc_hd__dfrtp_1
X_8429_ _8429_/A _8674_/B VGND VGND VPWR VPWR _8729_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold170 _5120_/X VGND VGND VPWR VPWR hold171/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 hold512/X VGND VGND VPWR VPWR hold511/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold181 hold181/A VGND VGND VPWR VPWR _9112_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5090_ _5090_/A VGND VGND VPWR VPWR _9707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7800_ _8230_/A VGND VGND VPWR VPWR _7904_/D sky130_fd_sc_hd__clkbuf_4
X_8780_ _8780_/A VGND VGND VPWR VPWR _8780_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5992_ _5992_/A VGND VGND VPWR VPWR _5992_/Y sky130_fd_sc_hd__inv_2
X_7731_ _7731_/A VGND VGND VPWR VPWR _7732_/A sky130_fd_sc_hd__clkbuf_1
X_4943_ _4943_/A _4953_/B VGND VGND VPWR VPWR _5543_/B sky130_fd_sc_hd__or2_4
XFILLER_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7662_ _6963_/Y _7491_/X _6831_/Y _7492_/X _7661_/X VGND VGND VPWR VPWR _7676_/B
+ sky130_fd_sc_hd__o221a_1
X_6613_ _9331_/Q VGND VGND VPWR VPWR _6613_/Y sky130_fd_sc_hd__clkinv_4
X_4874_ _9804_/Q VGND VGND VPWR VPWR _4874_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9401_ _9729_/CLK _9401_/D _9727_/SET_B VGND VGND VPWR VPWR _9401_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7593_ _6335_/Y _7500_/X _6294_/Y _7501_/X _7592_/X VGND VGND VPWR VPWR _7593_/X
+ sky130_fd_sc_hd__o221a_1
X_9332_ _9569_/CLK hold68/X _9563_/SET_B VGND VGND VPWR VPWR _9332_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6544_ _6539_/Y _5581_/B _8805_/A _5598_/B _6543_/X VGND VGND VPWR VPWR _6557_/B
+ sky130_fd_sc_hd__o221a_1
X_9263_ _9731_/CLK _9263_/D _9731_/SET_B VGND VGND VPWR VPWR _9263_/Q sky130_fd_sc_hd__dfrtp_1
X_6475_ _6475_/A VGND VGND VPWR VPWR _6475_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_173_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8214_ _8730_/A _8214_/B VGND VGND VPWR VPWR _8215_/B sky130_fd_sc_hd__or2_1
X_5426_ _9485_/Q _5419_/A _8969_/A1 _5419_/Y VGND VGND VPWR VPWR _9485_/D sky130_fd_sc_hd__a22o_1
Xoutput231 _8836_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_2
Xoutput220 _8816_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput253 _9036_/Z VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_2
X_9194_ _9416_/CLK _9194_/D _9731_/SET_B VGND VGND VPWR VPWR _9194_/Q sky130_fd_sc_hd__dfstp_1
Xoutput242 _7732_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_2
Xoutput264 _9046_/Z VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_2
Xoutput275 _8872_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_2
X_8145_ _8145_/A VGND VGND VPWR VPWR _8145_/Y sky130_fd_sc_hd__inv_2
Xoutput286 _7041_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_2
X_5357_ _9532_/Q _5353_/A _6067_/B1 _5353_/Y VGND VGND VPWR VPWR _9532_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8076_ _8076_/A _8502_/A VGND VGND VPWR VPWR _8076_/X sky130_fd_sc_hd__and2_1
Xoutput297 _9762_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_2
X_5288_ _9579_/Q _5284_/A _6067_/B1 _5284_/Y VGND VGND VPWR VPWR _9579_/D sky130_fd_sc_hd__a22o_1
X_7027_ _7092_/A _7106_/B VGND VGND VPWR VPWR _7027_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8978_ hold403/X hold405/X _9093_/Q VGND VGND VPWR VPWR _8978_/X sky130_fd_sc_hd__mux2_2
X_7929_ _7929_/A VGND VGND VPWR VPWR _8347_/B sky130_fd_sc_hd__buf_4
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4590_ _9795_/Q _4587_/A hold696/A _4587_/Y VGND VGND VPWR VPWR _9795_/D sky130_fd_sc_hd__a22o_1
XFILLER_155_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6260_ _6255_/Y _5935_/B _6256_/Y _4937_/X _6259_/X VGND VGND VPWR VPWR _6267_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5211_ _9629_/Q _5969_/A _5131_/X _4572_/X VGND VGND VPWR VPWR _9629_/D sky130_fd_sc_hd__a211o_1
XFILLER_142_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6191_ _9542_/Q VGND VGND VPWR VPWR _6191_/Y sky130_fd_sc_hd__inv_2
X_5142_ _9675_/Q _5135_/A _8969_/A1 _5135_/Y VGND VGND VPWR VPWR _9675_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5073_ _9714_/Q _5070_/A hold696/X _5070_/Y VGND VGND VPWR VPWR _9714_/D sky130_fd_sc_hd__a22o_1
XFILLER_111_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8901_ _7622_/Y _9680_/Q _9020_/S VGND VGND VPWR VPWR _8901_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8832_ _8832_/A VGND VGND VPWR VPWR _8832_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8763_ _8763_/A _8763_/B _8763_/C _8763_/D VGND VGND VPWR VPWR _8764_/C sky130_fd_sc_hd__or4_1
X_5975_ _9159_/Q _5973_/A _8964_/A1 _5973_/Y VGND VGND VPWR VPWR _9159_/D sky130_fd_sc_hd__a22o_1
X_8694_ _8723_/A _8764_/B _8723_/C VGND VGND VPWR VPWR _8694_/X sky130_fd_sc_hd__or3_1
X_4926_ _6189_/A _4848_/B _4923_/Y _4924_/Y _5436_/B VGND VGND VPWR VPWR _4926_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_40_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7714_ _6455_/Y _7485_/A _6393_/Y _7486_/A _7713_/X VGND VGND VPWR VPWR _7730_/A
+ sky130_fd_sc_hd__o221a_1
X_4857_ _9123_/Q VGND VGND VPWR VPWR _4857_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7645_ _4880_/Y _7498_/X _4739_/Y _5727_/X VGND VGND VPWR VPWR _7645_/X sky130_fd_sc_hd__o22a_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7576_ _6487_/Y _7497_/X _7573_/X _7575_/X VGND VGND VPWR VPWR _7586_/C sky130_fd_sc_hd__o211a_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9315_ _9574_/CLK _9315_/D _9571_/SET_B VGND VGND VPWR VPWR _9315_/Q sky130_fd_sc_hd__dfrtp_1
X_6527_ _9170_/Q VGND VGND VPWR VPWR _7733_/A sky130_fd_sc_hd__clkinv_4
X_4788_ _4784_/Y _5589_/B _4786_/Y _5990_/B VGND VGND VPWR VPWR _4788_/X sky130_fd_sc_hd__o22a_1
XFILLER_134_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9246_ _9695_/CLK _9246_/D _9537_/SET_B VGND VGND VPWR VPWR _9246_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_161_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6458_ _9540_/Q VGND VGND VPWR VPWR _6458_/Y sky130_fd_sc_hd__inv_2
X_5409_ _9499_/Q _5408_/A hold516/X _5408_/Y VGND VGND VPWR VPWR _5409_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6389_ _9814_/Q _6282_/Y _6388_/Y _4937_/X VGND VGND VPWR VPWR _6389_/X sky130_fd_sc_hd__o2bb2a_1
X_9177_ _9679_/CLK _9177_/D _9730_/SET_B VGND VGND VPWR VPWR _9177_/Q sky130_fd_sc_hd__dfstp_1
X_8128_ _8556_/B _8127_/Y VGND VGND VPWR VPWR _8338_/A sky130_fd_sc_hd__or2b_1
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8059_ _8654_/A _8056_/X _8059_/C _8483_/B VGND VGND VPWR VPWR _8059_/X sky130_fd_sc_hd__and4bb_1
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5760_ _9291_/Q _5759_/Y _5752_/Y VGND VGND VPWR VPWR _9291_/D sky130_fd_sc_hd__o21ba_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5691_ _9317_/Q _5689_/A hold510/X _5689_/Y VGND VGND VPWR VPWR _5691_/X sky130_fd_sc_hd__a22o_1
X_4711_ _4941_/A _4806_/B VGND VGND VPWR VPWR _5047_/B sky130_fd_sc_hd__or2_4
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4642_ _4689_/A _4642_/B _4689_/C _4708_/B VGND VGND VPWR VPWR _4915_/B sky130_fd_sc_hd__or4_4
X_7430_ _7467_/A _7471_/A _9297_/Q VGND VGND VPWR VPWR _9020_/S sky130_fd_sc_hd__nor3_4
XFILLER_175_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4573_ _7763_/A _5085_/D _9801_/Q _9002_/X _4572_/X VGND VGND VPWR VPWR _9801_/D
+ sky130_fd_sc_hd__a32o_1
Xhold703 _9319_/Q VGND VGND VPWR VPWR hold703/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_7361_ _6903_/Y _7180_/X _6916_/Y _7181_/X _7360_/X VGND VGND VPWR VPWR _7362_/D
+ sky130_fd_sc_hd__o221a_2
X_6312_ _8843_/A VGND VGND VPWR VPWR _6312_/Y sky130_fd_sc_hd__inv_2
X_7292_ _7292_/A _7380_/B VGND VGND VPWR VPWR _7292_/X sky130_fd_sc_hd__or2_1
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9100_ _9100_/CLK _9100_/D _6072_/X VGND VGND VPWR VPWR _9100_/Q sky130_fd_sc_hd__dfstp_2
X_9031_ _9616_/Q _8797_/A VGND VGND VPWR VPWR _9031_/Z sky130_fd_sc_hd__ebufn_1
X_6243_ _9199_/Q VGND VGND VPWR VPWR _6243_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6174_ _7314_/A _5636_/B _6170_/Y _5706_/B _6173_/X VGND VGND VPWR VPWR _6175_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5125_ _5125_/A VGND VGND VPWR VPWR _5125_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5056_ _5056_/A VGND VGND VPWR VPWR _5056_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8815_ _8815_/A VGND VGND VPWR VPWR _8816_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_111_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_9795_ _9798_/CLK _9795_/D _9797_/SET_B VGND VGND VPWR VPWR _9795_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5958_ _7809_/C _7809_/D _5958_/C VGND VGND VPWR VPWR _5966_/C sky130_fd_sc_hd__or3_1
X_8746_ _8746_/A _8746_/B VGND VGND VPWR VPWR _8747_/C sky130_fd_sc_hd__or2_1
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4909_ _9774_/Q VGND VGND VPWR VPWR _4909_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8677_ _8755_/B _8756_/A VGND VGND VPWR VPWR _8677_/Y sky130_fd_sc_hd__nor2_1
X_5889_ _5889_/A VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7628_ _6140_/Y _7502_/X _6141_/Y _7503_/X VGND VGND VPWR VPWR _7628_/X sky130_fd_sc_hd__o22a_1
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7559_ _8813_/A _7509_/X _8811_/A _7510_/X VGND VGND VPWR VPWR _7559_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_2_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9229_ _9418_/CLK _9229_/D _9730_/SET_B VGND VGND VPWR VPWR _9229_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_136_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold41 hold41/A VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold30 hold30/A VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold52 hold52/A VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold85 hold85/A VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_188_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_5 _5250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6930_ _6928_/Y _5839_/B _6929_/Y _5581_/B VGND VGND VPWR VPWR _6930_/X sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_6_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9574_/CLK sky130_fd_sc_hd__clkbuf_16
X_6861_ _6861_/A _6861_/B _6861_/C _6861_/D VGND VGND VPWR VPWR _6977_/A sky130_fd_sc_hd__and4_1
XFILLER_62_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8600_ _8600_/A VGND VGND VPWR VPWR _8730_/B sky130_fd_sc_hd__inv_2
X_5812_ _9263_/Q _5807_/A _8964_/A1 _5807_/Y VGND VGND VPWR VPWR _9263_/D sky130_fd_sc_hd__a22o_1
X_6792_ _9590_/Q VGND VGND VPWR VPWR _6792_/Y sky130_fd_sc_hd__inv_4
X_9580_ _9819_/CLK _9580_/D _7042_/B VGND VGND VPWR VPWR _9580_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8531_ _8762_/A _8755_/A _8745_/A VGND VGND VPWR VPWR _8645_/A sky130_fd_sc_hd__or3_1
Xclkbuf_1_0_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_1_0_1_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_62_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5743_ _9292_/Q VGND VGND VPWR VPWR _7025_/A sky130_fd_sc_hd__inv_2
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8462_ _8657_/B _8620_/A VGND VGND VPWR VPWR _8672_/C sky130_fd_sc_hd__or2_1
X_5674_ _9322_/Q VGND VGND VPWR VPWR _5675_/A sky130_fd_sc_hd__inv_2
X_8393_ _8682_/A _8420_/B _8682_/C VGND VGND VPWR VPWR _8394_/C sky130_fd_sc_hd__or3_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4625_ _4625_/A VGND VGND VPWR VPWR _4625_/Y sky130_fd_sc_hd__clkinv_2
X_7413_ _6378_/Y _7151_/A _6371_/Y _7152_/A VGND VGND VPWR VPWR _7413_/X sky130_fd_sc_hd__o22a_1
Xhold511 hold511/A VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold500 _4497_/X VGND VGND VPWR VPWR _4498_/A sky130_fd_sc_hd__clkdlybuf4s25_1
X_4556_ _4689_/C _4708_/B _4750_/C _4750_/D VGND VGND VPWR VPWR _4865_/A sky130_fd_sc_hd__or4_4
X_7344_ _6879_/Y _7135_/X _6855_/Y _7136_/X _7343_/X VGND VGND VPWR VPWR _7363_/A
+ sky130_fd_sc_hd__o221a_1
Xhold522 _5651_/X VGND VGND VPWR VPWR _9334_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold533 _5612_/X VGND VGND VPWR VPWR _9361_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold544 _5447_/X VGND VGND VPWR VPWR _9473_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_171_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold566 _5602_/X VGND VGND VPWR VPWR _9368_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold577 hold577/A VGND VGND VPWR VPWR hold696/A sky130_fd_sc_hd__buf_12
Xhold588 _5041_/X VGND VGND VPWR VPWR _9735_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7275_ _7275_/A _7275_/B _7275_/C VGND VGND VPWR VPWR _7275_/Y sky130_fd_sc_hd__nand3_4
XFILLER_131_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold555 _5294_/X VGND VGND VPWR VPWR _9576_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4487_ _4823_/B VGND VGND VPWR VPWR _4685_/B sky130_fd_sc_hd__inv_2
Xhold599 _5603_/X VGND VGND VPWR VPWR _9367_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6226_ _9516_/Q VGND VGND VPWR VPWR _6226_/Y sky130_fd_sc_hd__clkinv_2
X_9014_ _8697_/Y _8646_/X _9017_/S VGND VGND VPWR VPWR _9014_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6157_ _9267_/Q VGND VGND VPWR VPWR _6157_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5108_ _9698_/Q _5105_/A _8965_/A1 _5105_/Y VGND VGND VPWR VPWR _9698_/D sky130_fd_sc_hd__a22o_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6088_ _9087_/Q _6085_/A _8969_/A1 _6085_/Y VGND VGND VPWR VPWR _9087_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater394 _8964_/A1 VGND VGND VPWR VPWR _6065_/B1 sky130_fd_sc_hd__buf_12
X_5039_ _9737_/Q _5038_/A hold516/X _5038_/Y VGND VGND VPWR VPWR _5039_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9778_ _9819_/CLK _9778_/D _9817_/SET_B VGND VGND VPWR VPWR _9778_/Q sky130_fd_sc_hd__dfstp_1
X_8729_ _8762_/A _8729_/B _8729_/C VGND VGND VPWR VPWR _8755_/C sky130_fd_sc_hd__or3_1
XFILLER_21_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput120 sram_ro_data[5] VGND VGND VPWR VPWR _6301_/A sky130_fd_sc_hd__clkbuf_1
Xinput131 usr2_vdd_pwrgood VGND VGND VPWR VPWR _4889_/A sky130_fd_sc_hd__clkbuf_1
Xinput153 wb_adr_i[29] VGND VGND VPWR VPWR input153/X sky130_fd_sc_hd__clkbuf_1
Xinput142 wb_adr_i[19] VGND VGND VPWR VPWR _7803_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_48_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput164 wb_cyc_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput186 wb_dat_i[29] VGND VGND VPWR VPWR _7779_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput175 wb_dat_i[19] VGND VGND VPWR VPWR _7774_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_102_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput197 wb_rstn_i VGND VGND VPWR VPWR _6177_/A sky130_fd_sc_hd__buf_12
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5390_ _5390_/A VGND VGND VPWR VPWR _5391_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7060_ _7091_/C _7127_/B VGND VGND VPWR VPWR _7061_/A sky130_fd_sc_hd__or2_4
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6011_ _9132_/Q _6011_/B _9133_/Q VGND VGND VPWR VPWR _6011_/X sky130_fd_sc_hd__and3_1
XFILLER_39_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7962_ _8709_/A _7962_/B VGND VGND VPWR VPWR _7963_/B sky130_fd_sc_hd__or2_1
X_9701_ _4471_/A1 _9701_/D _6177_/A VGND VGND VPWR VPWR _9701_/Q sky130_fd_sc_hd__dfrtp_1
X_6913_ _6910_/Y _5826_/B _7178_/A _5636_/B _6912_/Y VGND VGND VPWR VPWR _6932_/A
+ sky130_fd_sc_hd__o221a_1
X_9632_ _9651_/CLK _9632_/D _9563_/SET_B VGND VGND VPWR VPWR _9632_/Q sky130_fd_sc_hd__dfrtp_1
X_7893_ _8557_/B _8312_/B VGND VGND VPWR VPWR _8657_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6844_ _6844_/A VGND VGND VPWR VPWR _6844_/Y sky130_fd_sc_hd__inv_2
X_9563_ _9569_/CLK _9563_/D _9563_/SET_B VGND VGND VPWR VPWR _9563_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_168_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6775_ _6775_/A VGND VGND VPWR VPWR _6775_/Y sky130_fd_sc_hd__inv_2
X_9494_ _9569_/CLK _9494_/D _9563_/SET_B VGND VGND VPWR VPWR _9494_/Q sky130_fd_sc_hd__dfrtp_1
X_8514_ _8514_/A VGND VGND VPWR VPWR _8514_/Y sky130_fd_sc_hd__clkinv_2
X_5726_ _7467_/A _7471_/A _7471_/C VGND VGND VPWR VPWR _5727_/A sky130_fd_sc_hd__or3_4
XFILLER_148_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8445_ _8445_/A VGND VGND VPWR VPWR _8707_/B sky130_fd_sc_hd__inv_2
XFILLER_190_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5657_ _9328_/Q _5649_/A hold601/A _5649_/Y VGND VGND VPWR VPWR _5657_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8376_ _8243_/A _8552_/A _8702_/A _8243_/A VGND VGND VPWR VPWR _8376_/X sky130_fd_sc_hd__o22a_1
X_4608_ _9782_/Q _4600_/A _6008_/B1 _4600_/Y VGND VGND VPWR VPWR _9782_/D sky130_fd_sc_hd__a22o_1
X_5588_ _9375_/Q _5583_/A _6008_/B1 _5583_/Y VGND VGND VPWR VPWR _9375_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold330 _5692_/X VGND VGND VPWR VPWR hold331/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 hold341/A VGND VGND VPWR VPWR hold341/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold352 _4890_/B VGND VGND VPWR VPWR hold353/A sky130_fd_sc_hd__dlygate4sd3_1
X_7327_ _4924_/Y _7095_/B _4726_/Y _7157_/X VGND VGND VPWR VPWR _7327_/X sky130_fd_sc_hd__o22a_1
X_4539_ _4643_/A VGND VGND VPWR VPWR _6189_/A sky130_fd_sc_hd__buf_4
Xhold374 _5204_/X VGND VGND VPWR VPWR hold375/A sky130_fd_sc_hd__dlygate4sd3_1
X_7258_ _6329_/Y _7144_/X _6328_/Y _7145_/X _7257_/X VGND VGND VPWR VPWR _7265_/A
+ sky130_fd_sc_hd__o221a_1
Xhold385 hold385/A VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold396 _8979_/X VGND VGND VPWR VPWR hold397/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _8991_/X VGND VGND VPWR VPWR hold364/A sky130_fd_sc_hd__dlygate4sd3_1
X_6209_ _9304_/Q VGND VGND VPWR VPWR _6209_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_131_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7189_ _6695_/Y _7137_/X _6724_/Y _7138_/X _7188_/X VGND VGND VPWR VPWR _7189_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4890_ _6142_/A _4890_/B VGND VGND VPWR VPWR _4890_/X sky130_fd_sc_hd__or2_4
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6560_ _9728_/Q VGND VGND VPWR VPWR _6560_/Y sky130_fd_sc_hd__inv_2
X_5511_ _9428_/Q _5507_/A _6067_/B1 _5507_/Y VGND VGND VPWR VPWR _9428_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6491_ _8850_/B _6165_/A _6487_/Y _5979_/B _6490_/X VGND VGND VPWR VPWR _6504_/B
+ sky130_fd_sc_hd__o221a_1
X_8230_ _8230_/A _8255_/A VGND VGND VPWR VPWR _8230_/Y sky130_fd_sc_hd__nor2_1
XFILLER_145_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5442_ _9475_/Q _5438_/A _6067_/B1 _5438_/Y VGND VGND VPWR VPWR _9475_/D sky130_fd_sc_hd__a22o_1
X_8161_ _8161_/A _8161_/B VGND VGND VPWR VPWR _8439_/B sky130_fd_sc_hd__or2_4
XFILLER_160_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5373_ _9522_/Q _5369_/A _8959_/A1 _5369_/Y VGND VGND VPWR VPWR _9522_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_24_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9225_/CLK sky130_fd_sc_hd__clkbuf_16
X_8092_ _8092_/A VGND VGND VPWR VPWR _8209_/A sky130_fd_sc_hd__buf_2
X_7112_ _4753_/Y _7155_/A _4765_/Y _7156_/A _7111_/X VGND VGND VPWR VPWR _7116_/C
+ sky130_fd_sc_hd__o221a_1
X_7043_ _9668_/Q input86/X VGND VGND VPWR VPWR _7044_/A sky130_fd_sc_hd__or2b_1
XFILLER_86_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9431_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8994_ _9753_/Q _6977_/Y _8999_/S VGND VGND VPWR VPWR _8994_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7945_ _7903_/A _7924_/B _7935_/X _7941_/X _7944_/X VGND VGND VPWR VPWR _7945_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7876_ _7876_/A VGND VGND VPWR VPWR _8140_/A sky130_fd_sc_hd__inv_2
XFILLER_63_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9615_ _9731_/CLK _9615_/D _9731_/SET_B VGND VGND VPWR VPWR _9615_/Q sky130_fd_sc_hd__dfrtp_1
X_6827_ _9791_/Q VGND VGND VPWR VPWR _6827_/Y sky130_fd_sc_hd__inv_2
X_9546_ _9550_/CLK _9546_/D _9537_/SET_B VGND VGND VPWR VPWR _9546_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6758_ _6756_/Y _5255_/B _6757_/Y _4844_/X VGND VGND VPWR VPWR _6758_/X sky130_fd_sc_hd__o22a_2
X_5709_ _9305_/Q _5708_/A hold516/X _5708_/Y VGND VGND VPWR VPWR _5709_/X sky130_fd_sc_hd__a22o_1
X_6689_ _9830_/Q VGND VGND VPWR VPWR _6689_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9477_ _9483_/CLK _9477_/D _9727_/SET_B VGND VGND VPWR VPWR _9477_/Q sky130_fd_sc_hd__dfrtp_1
X_8428_ _8428_/A _8428_/B VGND VGND VPWR VPWR _8674_/B sky130_fd_sc_hd__or2_2
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8359_ _8359_/A _8359_/B VGND VGND VPWR VPWR _8639_/C sky130_fd_sc_hd__or2_1
Xhold171 hold171/A VGND VGND VPWR VPWR hold172/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 hold160/A VGND VGND VPWR VPWR _9632_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold193 hold511/X VGND VGND VPWR VPWR hold510/A sky130_fd_sc_hd__buf_12
Xhold182 _5454_/X VGND VGND VPWR VPWR hold183/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5991_ _5991_/A VGND VGND VPWR VPWR _5992_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7730_ _7730_/A _7730_/B _7730_/C _7730_/D VGND VGND VPWR VPWR _7730_/Y sky130_fd_sc_hd__nand4_2
X_4942_ _9401_/Q VGND VGND VPWR VPWR _4942_/Y sky130_fd_sc_hd__clkinv_2
X_7661_ _6971_/Y _7493_/X _6899_/Y _7494_/X VGND VGND VPWR VPWR _7661_/X sky130_fd_sc_hd__o22a_1
X_9400_ _9831_/CLK _9400_/D _9727_/SET_B VGND VGND VPWR VPWR _9400_/Q sky130_fd_sc_hd__dfrtp_1
X_4873_ _4933_/A _4920_/A VGND VGND VPWR VPWR _5378_/B sky130_fd_sc_hd__or2_4
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6612_ _9257_/Q VGND VGND VPWR VPWR _6612_/Y sky130_fd_sc_hd__inv_2
X_7592_ _6306_/Y _7502_/X _6271_/Y _7503_/X VGND VGND VPWR VPWR _7592_/X sky130_fd_sc_hd__o22a_1
X_9331_ _9391_/CLK hold89/X _9563_/SET_B VGND VGND VPWR VPWR _9331_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6543_ _6541_/Y _5698_/B _8795_/A _5805_/B VGND VGND VPWR VPWR _6543_/X sky130_fd_sc_hd__o22a_1
X_9262_ _9734_/CLK _9262_/D _9731_/SET_B VGND VGND VPWR VPWR _9262_/Q sky130_fd_sc_hd__dfrtp_1
X_6474_ _6469_/Y _4863_/X _6470_/Y _5112_/B _6473_/X VGND VGND VPWR VPWR _6474_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_173_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput210 _8798_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_118_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8213_ _8213_/A _8415_/A _8212_/X VGND VGND VPWR VPWR _8214_/B sky130_fd_sc_hd__or3b_1
X_5425_ _9486_/Q _5419_/A _8965_/A1 _5419_/Y VGND VGND VPWR VPWR _9486_/D sky130_fd_sc_hd__a22o_1
Xoutput221 _8818_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_2
Xoutput232 _8838_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_160_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9193_ _9491_/CLK _9193_/D _9731_/SET_B VGND VGND VPWR VPWR _9193_/Q sky130_fd_sc_hd__dfstp_1
Xoutput243 _8790_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_2
Xoutput265 _9047_/Z VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_2
Xoutput254 _9037_/Z VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_2
X_8144_ _8236_/A _8144_/B VGND VGND VPWR VPWR _8145_/A sky130_fd_sc_hd__or2_1
XFILLER_160_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5356_ _9533_/Q _5353_/A hold217/X _5353_/Y VGND VGND VPWR VPWR _9533_/D sky130_fd_sc_hd__a22o_1
Xoutput276 _9022_/Z VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_99_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8075_ _8666_/B _8593_/A VGND VGND VPWR VPWR _8502_/A sky130_fd_sc_hd__or2_1
Xoutput298 _9763_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_2
Xoutput287 _8880_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_2
X_5287_ _9580_/Q _5284_/A hold217/X _5284_/Y VGND VGND VPWR VPWR _9580_/D sky130_fd_sc_hd__a22o_1
X_7026_ _9290_/Q _7081_/B _7128_/A VGND VGND VPWR VPWR _7106_/B sky130_fd_sc_hd__or3_1
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8977_ _8976_/X hold368/X _9629_/Q VGND VGND VPWR VPWR _8977_/X sky130_fd_sc_hd__mux2_4
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7928_ _8567_/A _8230_/A _7942_/C _8234_/A VGND VGND VPWR VPWR _7929_/A sky130_fd_sc_hd__or4_1
XFILLER_82_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7859_ _8243_/A _8314_/A VGND VGND VPWR VPWR _8745_/A sky130_fd_sc_hd__nor2_4
XFILLER_156_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9529_ _9800_/CLK _9529_/D _9817_/SET_B VGND VGND VPWR VPWR _9529_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5210_ _9101_/Q VGND VGND VPWR VPWR _5969_/A sky130_fd_sc_hd__inv_2
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6190_ _9498_/Q VGND VGND VPWR VPWR _6190_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_89_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5141_ _9676_/Q _5135_/A _8965_/A1 _5135_/Y VGND VGND VPWR VPWR _9676_/D sky130_fd_sc_hd__a22o_1
X_5072_ _9715_/Q _5070_/A hold510/X _5070_/Y VGND VGND VPWR VPWR _9715_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8900_ _8899_/X _9210_/Q _9096_/Q VGND VGND VPWR VPWR _8900_/X sky130_fd_sc_hd__mux2_1
X_8831_ _8831_/A VGND VGND VPWR VPWR _8832_/A sky130_fd_sc_hd__clkbuf_1
X_8762_ _8762_/A _8762_/B _8762_/C VGND VGND VPWR VPWR _8763_/D sky130_fd_sc_hd__or3_1
XFILLER_64_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5974_ _9160_/Q _5973_/A _8959_/A1 _5973_/Y VGND VGND VPWR VPWR _9160_/D sky130_fd_sc_hd__a22o_1
X_7713_ _6430_/Y _7487_/A _6449_/Y _7488_/A VGND VGND VPWR VPWR _7713_/X sky130_fd_sc_hd__o22a_1
X_8693_ _8693_/A _8693_/B VGND VGND VPWR VPWR _8723_/C sky130_fd_sc_hd__or2_1
X_4925_ _4925_/A _4925_/B VGND VGND VPWR VPWR _5436_/B sky130_fd_sc_hd__or2_4
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4856_ _4913_/B _4898_/B VGND VGND VPWR VPWR _5455_/B sky130_fd_sc_hd__or2_4
X_7644_ _4733_/Y _7491_/X _4805_/Y _7492_/X _7643_/X VGND VGND VPWR VPWR _7658_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7575_ _6368_/Y _7500_/X _6433_/Y _7501_/X _7574_/X VGND VGND VPWR VPWR _7575_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9314_ _9522_/CLK _9314_/D _9537_/SET_B VGND VGND VPWR VPWR _9314_/Q sky130_fd_sc_hd__dfrtp_1
X_6526_ _9326_/Q VGND VGND VPWR VPWR _7402_/A sky130_fd_sc_hd__inv_2
X_4787_ _6142_/B _4865_/B VGND VGND VPWR VPWR _5990_/B sky130_fd_sc_hd__or2_4
XFILLER_146_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6457_ _6452_/Y _5521_/B _6453_/Y _5417_/B _6456_/X VGND VGND VPWR VPWR _6464_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9245_ _9322_/CLK _9245_/D _9797_/SET_B VGND VGND VPWR VPWR _9245_/Q sky130_fd_sc_hd__dfrtp_1
X_5408_ _5408_/A VGND VGND VPWR VPWR _5408_/Y sky130_fd_sc_hd__clkinv_2
X_6388_ _9470_/Q VGND VGND VPWR VPWR _6388_/Y sky130_fd_sc_hd__clkinv_2
X_9176_ _9679_/CLK _9176_/D _9730_/SET_B VGND VGND VPWR VPWR _9176_/Q sky130_fd_sc_hd__dfrtp_1
X_8127_ _8127_/A _8127_/B VGND VGND VPWR VPWR _8127_/Y sky130_fd_sc_hd__nand2_1
X_5339_ _9544_/Q _5331_/A hold601/X _5331_/Y VGND VGND VPWR VPWR _5339_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8058_ _8065_/A _8443_/A VGND VGND VPWR VPWR _8483_/B sky130_fd_sc_hd__or2_1
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7009_ _6268_/Y _7007_/A _9060_/Q _7007_/Y VGND VGND VPWR VPWR _9060_/D sky130_fd_sc_hd__o22a_1
XFILLER_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5690_ _9318_/Q _5689_/A hold516/X _5689_/Y VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__a22o_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _9725_/Q VGND VGND VPWR VPWR _4712_/A sky130_fd_sc_hd__clkinv_2
X_4641_ _9763_/Q _4636_/A _6008_/B1 _4636_/Y VGND VGND VPWR VPWR _4641_/X sky130_fd_sc_hd__a22o_1
X_4572_ _9107_/Q _4572_/B VGND VGND VPWR VPWR _4572_/X sky130_fd_sc_hd__or2_1
X_7360_ _6843_/Y _7182_/X _6899_/Y _7183_/X VGND VGND VPWR VPWR _7360_/X sky130_fd_sc_hd__o22a_1
Xhold704 _8886_/X VGND VGND VPWR VPWR hold704/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7291_ _6249_/Y _7171_/X _6183_/Y _7172_/X _7290_/X VGND VGND VPWR VPWR _7296_/B
+ sky130_fd_sc_hd__o221a_1
X_6311_ _6311_/A _6311_/B _6311_/C _6311_/D VGND VGND VPWR VPWR _6357_/B sky130_fd_sc_hd__and4_4
X_9030_ _9615_/Q _8795_/A VGND VGND VPWR VPWR _9030_/Z sky130_fd_sc_hd__ebufn_1
X_6242_ _6242_/A _6242_/B _6242_/C _6242_/D VGND VGND VPWR VPWR _6268_/C sky130_fd_sc_hd__and4_1
XFILLER_69_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6173_ _6171_/Y _5847_/B _6172_/Y _5598_/B VGND VGND VPWR VPWR _6173_/X sky130_fd_sc_hd__o22a_1
X_5124_ _5124_/A VGND VGND VPWR VPWR _5125_/A sky130_fd_sc_hd__clkbuf_2
X_5055_ _6017_/A VGND VGND VPWR VPWR _5056_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8814_ _8814_/A VGND VGND VPWR VPWR _8814_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9794_ _9798_/CLK _9794_/D _9821_/SET_B VGND VGND VPWR VPWR _9794_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5957_ _7806_/A _7806_/B _7806_/C _7806_/D VGND VGND VPWR VPWR _5958_/C sky130_fd_sc_hd__or4_1
X_8745_ _8745_/A _8745_/B _8745_/C _8745_/D VGND VGND VPWR VPWR _8748_/C sky130_fd_sc_hd__or4_1
XFILLER_71_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8676_ _8586_/A _8133_/Y _8629_/A _8473_/A VGND VGND VPWR VPWR _8756_/A sky130_fd_sc_hd__a211o_2
X_4908_ _4904_/Y _4525_/B _4905_/Y _5282_/B _4907_/X VGND VGND VPWR VPWR _4918_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_166_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7627_ _6103_/Y _7498_/X _6172_/Y _5727_/X VGND VGND VPWR VPWR _7627_/X sky130_fd_sc_hd__o22a_1
X_5888_ _5878_/X _8896_/X _8960_/X _9209_/Q VGND VGND VPWR VPWR _9209_/D sky130_fd_sc_hd__o22a_1
XFILLER_166_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4839_ _4933_/A _4949_/A VGND VGND VPWR VPWR _5417_/B sky130_fd_sc_hd__or2_4
XFILLER_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7558_ _7735_/A _7497_/X _7555_/X _7557_/X VGND VGND VPWR VPWR _7568_/C sky130_fd_sc_hd__o211a_1
X_6509_ _9301_/Q VGND VGND VPWR VPWR _8799_/A sky130_fd_sc_hd__inv_6
XFILLER_153_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7489_ _6896_/Y _7487_/X _6944_/Y _7488_/X VGND VGND VPWR VPWR _7489_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9228_ _9679_/CLK _9228_/D _9730_/SET_B VGND VGND VPWR VPWR _9228_/Q sky130_fd_sc_hd__dfrtp_1
X_9159_ _9730_/CLK _9159_/D _9730_/SET_B VGND VGND VPWR VPWR _9159_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold20 hold20/A VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold64 hold64/A VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__buf_12
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__buf_12
Xhold97 hold97/A VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold75 hold75/A VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_6 _4502_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6860_ _6860_/A _6860_/B _6860_/C _6860_/D VGND VGND VPWR VPWR _6861_/D sky130_fd_sc_hd__and4_1
XFILLER_179_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6791_ _9546_/Q VGND VGND VPWR VPWR _6791_/Y sky130_fd_sc_hd__inv_4
X_5811_ _9264_/Q _5807_/A _8959_/A1 _5807_/Y VGND VGND VPWR VPWR _9264_/D sky130_fd_sc_hd__a22o_1
XFILLER_62_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8530_ _8530_/A VGND VGND VPWR VPWR _8530_/X sky130_fd_sc_hd__clkbuf_1
X_5742_ _7432_/B _9097_/Q _9293_/Q _5741_/Y VGND VGND VPWR VPWR _9293_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8461_ _8594_/A _8443_/B _8457_/X _8460_/Y VGND VGND VPWR VPWR _8461_/X sky130_fd_sc_hd__o211a_1
X_5673_ _5673_/A _5685_/A _5780_/C VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__or3_1
X_8392_ _8625_/A _8625_/B _8392_/C VGND VGND VPWR VPWR _8682_/C sky130_fd_sc_hd__or3_2
X_4624_ _4624_/A VGND VGND VPWR VPWR _4625_/A sky130_fd_sc_hd__buf_2
X_7412_ _6498_/Y _7144_/A _6447_/Y _7145_/A _7411_/X VGND VGND VPWR VPWR _7419_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold501 _4832_/A VGND VGND VPWR VPWR _4913_/A sky130_fd_sc_hd__clkbuf_2
X_7343_ _6958_/Y _7137_/X _6935_/Y _7138_/X _7342_/X VGND VGND VPWR VPWR _7343_/X
+ sky130_fd_sc_hd__o221a_1
X_4555_ _9804_/Q _4547_/A _6008_/B1 _4547_/Y VGND VGND VPWR VPWR _4555_/X sky130_fd_sc_hd__a22o_1
Xhold512 _8887_/X VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold534 _5574_/X VGND VGND VPWR VPWR _9386_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold545 _5293_/X VGND VGND VPWR VPWR _9577_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold523 _6002_/X VGND VGND VPWR VPWR _9141_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold578 hold578/A VGND VGND VPWR VPWR hold578/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold567 _5850_/X VGND VGND VPWR VPWR _9239_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold556 _5690_/X VGND VGND VPWR VPWR _9318_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_131_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9013_ _8632_/Y _8555_/X _9017_/S VGND VGND VPWR VPWR _9013_/X sky130_fd_sc_hd__mux2_1
X_7274_ _7274_/A _7274_/B _7274_/C _7274_/D VGND VGND VPWR VPWR _7275_/C sky130_fd_sc_hd__and4_1
X_4486_ _9832_/Q _4485_/A hold510/X _4485_/Y VGND VGND VPWR VPWR _9832_/D sky130_fd_sc_hd__a22o_1
Xhold589 _5869_/X VGND VGND VPWR VPWR _9226_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6225_ _9225_/Q VGND VGND VPWR VPWR _6225_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_103_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6156_ _6151_/Y _5036_/B _6152_/Y _5826_/B _6155_/X VGND VGND VPWR VPWR _6175_/A
+ sky130_fd_sc_hd__o221a_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _9699_/Q _5105_/A _8964_/A1 _5105_/Y VGND VGND VPWR VPWR _9699_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6087_ _9088_/Q _6085_/A _8965_/A1 _6085_/Y VGND VGND VPWR VPWR _9088_/D sky130_fd_sc_hd__a22o_1
Xrepeater395 hold42/X VGND VGND VPWR VPWR _8964_/A1 sky130_fd_sc_hd__buf_12
X_5038_ _5038_/A VGND VGND VPWR VPWR _5038_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_167_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9777_ _9819_/CLK _9777_/D _9821_/SET_B VGND VGND VPWR VPWR _9777_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6989_ _6816_/Y _6983_/A _9072_/Q _6983_/Y VGND VGND VPWR VPWR _9072_/D sky130_fd_sc_hd__o22a_1
X_8728_ _8728_/A _8728_/B _8728_/C _8728_/D VGND VGND VPWR VPWR _8751_/D sky130_fd_sc_hd__or4_2
XFILLER_80_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8659_ _8659_/A _8659_/B VGND VGND VPWR VPWR _8749_/A sky130_fd_sc_hd__or2_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput110 sram_ro_data[25] VGND VGND VPWR VPWR _6848_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput154 wb_adr_i[2] VGND VGND VPWR VPWR _8421_/B sky130_fd_sc_hd__buf_6
Xinput143 wb_adr_i[1] VGND VGND VPWR VPWR _8436_/C sky130_fd_sc_hd__buf_4
Xinput132 wb_adr_i[0] VGND VGND VPWR VPWR _7876_/A sky130_fd_sc_hd__buf_4
XFILLER_88_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput121 sram_ro_data[6] VGND VGND VPWR VPWR _6264_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_48_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput187 wb_dat_i[2] VGND VGND VPWR VPWR _9005_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput176 wb_dat_i[1] VGND VGND VPWR VPWR _9004_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_dat_i[0] VGND VGND VPWR VPWR _9003_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput198 wb_sel_i[0] VGND VGND VPWR VPWR _5082_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6010_ _6010_/A VGND VGND VPWR VPWR _6010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7961_ _7873_/B _8341_/B _7901_/Y _7960_/Y VGND VGND VPWR VPWR _7962_/B sky130_fd_sc_hd__a31o_1
X_6912_ input47/X _8973_/S input53/X _6353_/Y VGND VGND VPWR VPWR _6912_/Y sky130_fd_sc_hd__a22oi_2
X_7892_ _8563_/B _8312_/B VGND VGND VPWR VPWR _8367_/A sky130_fd_sc_hd__or2_1
XFILLER_82_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9700_ _9833_/CLK _9700_/D _9730_/SET_B VGND VGND VPWR VPWR _9700_/Q sky130_fd_sc_hd__dfrtp_1
X_9631_ _9643_/CLK _9631_/D _9563_/SET_B VGND VGND VPWR VPWR _9631_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6843_ _9816_/Q VGND VGND VPWR VPWR _6843_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9562_ _9569_/CLK _9562_/D _9563_/SET_B VGND VGND VPWR VPWR _9562_/Q sky130_fd_sc_hd__dfstp_1
X_6774_ _9164_/Q VGND VGND VPWR VPWR _6774_/Y sky130_fd_sc_hd__clkinv_2
X_9493_ _9569_/CLK _9493_/D _9563_/SET_B VGND VGND VPWR VPWR _9493_/Q sky130_fd_sc_hd__dfstp_1
X_8513_ _8580_/C VGND VGND VPWR VPWR _8513_/Y sky130_fd_sc_hd__clkinv_2
X_5725_ _7478_/D VGND VGND VPWR VPWR _7471_/C sky130_fd_sc_hd__buf_2
X_5656_ _9329_/Q hold639/X hold593/X _5649_/Y VGND VGND VPWR VPWR _9329_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8444_ _8243_/B _8158_/A _8059_/C _8442_/X _8443_/X VGND VGND VPWR VPWR _8444_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_190_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4607_ _9783_/Q _4600_/A _6067_/B1 _4600_/Y VGND VGND VPWR VPWR _9783_/D sky130_fd_sc_hd__a22o_1
XFILLER_184_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold320 hold320/A VGND VGND VPWR VPWR _9693_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_8375_ _8762_/A _8755_/A _8375_/C VGND VGND VPWR VPWR _8377_/A sky130_fd_sc_hd__or3_1
X_5587_ _9376_/Q _5583_/A _6067_/B1 _5583_/Y VGND VGND VPWR VPWR _9376_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold331 hold331/A VGND VGND VPWR VPWR hold332/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold342 _8982_/X VGND VGND VPWR VPWR hold343/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 hold353/A VGND VGND VPWR VPWR hold354/A sky130_fd_sc_hd__dlygate4sd3_1
X_4538_ _9813_/Q _4537_/Y _6008_/B1 _4537_/A _4473_/A VGND VGND VPWR VPWR _4538_/X
+ sky130_fd_sc_hd__o221a_1
X_7326_ _4946_/Y _7149_/X _4743_/Y _7150_/X _7325_/X VGND VGND VPWR VPWR _7331_/B
+ sky130_fd_sc_hd__o221a_1
Xhold375 hold375/A VGND VGND VPWR VPWR hold376/A sky130_fd_sc_hd__dlygate4sd3_1
X_7257_ _6313_/Y _7071_/C _6335_/Y _7146_/X VGND VGND VPWR VPWR _7257_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4469_ _9626_/Q input77/X _8843_/B VGND VGND VPWR VPWR _9025_/A sky130_fd_sc_hd__mux2_1
Xhold386 _5557_/X VGND VGND VPWR VPWR hold387/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 hold364/A VGND VGND VPWR VPWR hold365/A sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ _6206_/Y _5847_/B _6207_/Y _5598_/B VGND VGND VPWR VPWR _6218_/A sky130_fd_sc_hd__o22a_1
Xhold397 hold397/A VGND VGND VPWR VPWR hold398/A sky130_fd_sc_hd__dlygate4sd3_1
X_7188_ _6744_/Y _7139_/X _6741_/Y _7140_/X VGND VGND VPWR VPWR _7188_/X sky130_fd_sc_hd__o22a_1
XFILLER_58_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6139_ _6134_/Y _5455_/B _6135_/Y _6058_/B _6138_/X VGND VGND VPWR VPWR _6150_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9829_ _9832_/CLK _9829_/D _9821_/SET_B VGND VGND VPWR VPWR _9829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_csclk clkbuf_leaf_5_csclk/A VGND VGND VPWR VPWR _9326_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5510_ _9429_/Q _5507_/A hold217/A _5507_/Y VGND VGND VPWR VPWR _9429_/D sky130_fd_sc_hd__a22o_1
X_6490_ _6488_/Y _5866_/B _6489_/Y _5990_/B VGND VGND VPWR VPWR _6490_/X sky130_fd_sc_hd__o22a_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5441_ _9476_/Q _5438_/A hold217/X _5438_/Y VGND VGND VPWR VPWR _9476_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5372_ _9523_/Q _5369_/A hold577/A _5369_/Y VGND VGND VPWR VPWR _5372_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8160_ _8160_/A VGND VGND VPWR VPWR _8588_/A sky130_fd_sc_hd__inv_2
XFILLER_160_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8091_ _8137_/B _8091_/B VGND VGND VPWR VPWR _8092_/A sky130_fd_sc_hd__or2_1
X_7111_ _4855_/Y _7056_/A _4747_/Y _7157_/A VGND VGND VPWR VPWR _7111_/X sky130_fd_sc_hd__o22a_1
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7042_ _9628_/Q _7042_/B VGND VGND VPWR VPWR _7042_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8993_ _9754_/Q _6816_/Y _8999_/S VGND VGND VPWR VPWR _8993_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7944_ _8489_/A _8042_/B _8383_/B _7935_/A _8540_/A VGND VGND VPWR VPWR _7944_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_82_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7875_ _8421_/D _7875_/B _8436_/D _7918_/A VGND VGND VPWR VPWR _8340_/A sky130_fd_sc_hd__or4_2
X_9614_ _9731_/CLK _9614_/D _9731_/SET_B VGND VGND VPWR VPWR _9614_/Q sky130_fd_sc_hd__dfrtp_1
X_6826_ _9802_/Q VGND VGND VPWR VPWR _6826_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9545_ _9577_/CLK _9545_/D _9571_/SET_B VGND VGND VPWR VPWR _9545_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6757_ _6757_/A VGND VGND VPWR VPWR _6757_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5708_ _5708_/A VGND VGND VPWR VPWR _5708_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6688_ _9476_/Q VGND VGND VPWR VPWR _6688_/Y sky130_fd_sc_hd__inv_2
X_9476_ _9483_/CLK _9476_/D _9727_/SET_B VGND VGND VPWR VPWR _9476_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8427_ _8692_/C _8427_/B VGND VGND VPWR VPWR _8478_/A sky130_fd_sc_hd__or2_1
X_5639_ _9343_/Q _5638_/A hold516/X _5638_/Y VGND VGND VPWR VPWR _5639_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8358_ _8358_/A _8540_/B VGND VGND VPWR VPWR _8532_/C sky130_fd_sc_hd__nor2_1
XFILLER_191_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold150 hold150/A VGND VGND VPWR VPWR hold151/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _5337_/X VGND VGND VPWR VPWR hold162/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7309_ _7309_/A _7309_/B _7309_/C _7309_/D VGND VGND VPWR VPWR _7319_/B sky130_fd_sc_hd__and4_1
Xhold172 hold172/A VGND VGND VPWR VPWR _9690_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold194 _6062_/X VGND VGND VPWR VPWR hold195/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/A VGND VGND VPWR VPWR hold184/A sky130_fd_sc_hd__dlygate4sd3_1
X_8289_ _8361_/A _8306_/B VGND VGND VPWR VPWR _8359_/B sky130_fd_sc_hd__nor2_1
XFILLER_132_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5990_ _5990_/A _5990_/B VGND VGND VPWR VPWR _5991_/A sky130_fd_sc_hd__or2_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4941_ _4941_/A _4953_/B VGND VGND VPWR VPWR _5505_/B sky130_fd_sc_hd__or2_4
X_4872_ _9510_/Q VGND VGND VPWR VPWR _4872_/Y sky130_fd_sc_hd__clkinv_4
X_7660_ _6832_/Y _7485_/X _6958_/Y _7486_/X _7659_/X VGND VGND VPWR VPWR _7676_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6611_ _9733_/Q VGND VGND VPWR VPWR _8787_/A sky130_fd_sc_hd__clkinv_4
XFILLER_60_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9330_ _9391_/CLK _9330_/D _9563_/SET_B VGND VGND VPWR VPWR _9330_/Q sky130_fd_sc_hd__dfrtp_1
X_7591_ _6277_/Y _7498_/X _6351_/Y _5727_/X VGND VGND VPWR VPWR _7591_/X sky130_fd_sc_hd__o22a_1
XFILLER_32_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6542_ _9263_/Q VGND VGND VPWR VPWR _8795_/A sky130_fd_sc_hd__inv_4
XFILLER_192_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9261_ _9734_/CLK _9261_/D _9731_/SET_B VGND VGND VPWR VPWR _9261_/Q sky130_fd_sc_hd__dfstp_1
X_6473_ _6471_/Y _5551_/B _6472_/Y _5927_/B VGND VGND VPWR VPWR _6473_/X sky130_fd_sc_hd__o22a_1
X_8212_ _8438_/A _8439_/B VGND VGND VPWR VPWR _8212_/X sky130_fd_sc_hd__or2_1
XFILLER_106_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5424_ _9487_/Q _5419_/A _8964_/A1 _5419_/Y VGND VGND VPWR VPWR _9487_/D sky130_fd_sc_hd__a22o_1
X_9192_ _9322_/CLK _9192_/D _9797_/SET_B VGND VGND VPWR VPWR _9192_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput233 _8840_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_2
Xoutput222 _8820_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_2
X_8143_ _8243_/B VGND VGND VPWR VPWR _8667_/A sky130_fd_sc_hd__inv_2
XFILLER_160_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput211 _8800_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput244 _8792_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_2
Xoutput266 _9048_/Z VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_2
Xoutput255 _9038_/Z VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_2
X_5355_ _9534_/Q _5353_/A _6065_/B1 _5353_/Y VGND VGND VPWR VPWR _9534_/D sky130_fd_sc_hd__a22o_1
Xoutput277 _9023_/Z VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_2
X_8074_ _8074_/A _8656_/B VGND VGND VPWR VPWR _8076_/A sky130_fd_sc_hd__nor2_1
Xoutput299 _9764_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_2
Xoutput288 _7045_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_2
X_5286_ _9581_/Q _5284_/A _6065_/B1 _5284_/Y VGND VGND VPWR VPWR _9581_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7025_ _7025_/A _9291_/Q VGND VGND VPWR VPWR _7092_/A sky130_fd_sc_hd__or2_2
XFILLER_83_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8976_ hold405/X hold672/X _9093_/Q VGND VGND VPWR VPWR _8976_/X sky130_fd_sc_hd__mux2_2
XFILLER_55_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7927_ _8489_/A _7953_/A VGND VGND VPWR VPWR _7935_/A sky130_fd_sc_hd__or2_1
X_7858_ _8436_/A _8436_/B _7875_/B VGND VGND VPWR VPWR _8314_/A sky130_fd_sc_hd__or3_4
XFILLER_130_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6809_ _6809_/A VGND VGND VPWR VPWR _6809_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7789_ _7869_/A _7789_/B _7874_/C VGND VGND VPWR VPWR _7790_/A sky130_fd_sc_hd__or3_1
XFILLER_23_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9528_ _9800_/CLK _9528_/D _9817_/SET_B VGND VGND VPWR VPWR _9528_/Q sky130_fd_sc_hd__dfstp_1
X_9459_ _9550_/CLK _9459_/D _9537_/SET_B VGND VGND VPWR VPWR _9459_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_136_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9830_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9600_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5140_ _9677_/Q _5135_/A _8964_/A1 _5135_/Y VGND VGND VPWR VPWR _9677_/D sky130_fd_sc_hd__a22o_1
X_5071_ _9716_/Q _5070_/A hold516/X _5070_/Y VGND VGND VPWR VPWR _5071_/X sky130_fd_sc_hd__a22o_1
XFILLER_111_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8830_ _8830_/A VGND VGND VPWR VPWR _8830_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8761_ _8761_/A _8761_/B _8761_/C VGND VGND VPWR VPWR _8773_/C sky130_fd_sc_hd__or3_2
X_5973_ _5973_/A VGND VGND VPWR VPWR _5973_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4924_ _9474_/Q VGND VGND VPWR VPWR _4924_/Y sky130_fd_sc_hd__inv_2
X_7712_ _7712_/A _7712_/B _7712_/C _7712_/D VGND VGND VPWR VPWR _7712_/Y sky130_fd_sc_hd__nand4_1
XFILLER_52_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8692_ _8714_/C _8692_/B _8692_/C VGND VGND VPWR VPWR _8764_/B sky130_fd_sc_hd__or3_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4855_ _9458_/Q VGND VGND VPWR VPWR _4855_/Y sky130_fd_sc_hd__clkinv_4
X_7643_ _4697_/Y _7493_/X _4831_/Y _7494_/X VGND VGND VPWR VPWR _7643_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7574_ _6377_/Y _7502_/X _6360_/Y _7503_/X VGND VGND VPWR VPWR _7574_/X sky130_fd_sc_hd__o22a_1
X_4786_ _9143_/Q VGND VGND VPWR VPWR _4786_/Y sky130_fd_sc_hd__inv_2
X_6525_ _8839_/A _6112_/B _7737_/A _4865_/X _6524_/X VGND VGND VPWR VPWR _6532_/C
+ sky130_fd_sc_hd__o221a_1
X_9313_ _9318_/CLK _9313_/D _9571_/SET_B VGND VGND VPWR VPWR _9313_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9244_ _9600_/CLK _9244_/D _9821_/SET_B VGND VGND VPWR VPWR _9244_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6456_ _6454_/Y _5474_/B _6455_/Y _5543_/B VGND VGND VPWR VPWR _6456_/X sky130_fd_sc_hd__o22a_2
X_6387_ _9332_/Q VGND VGND VPWR VPWR _6387_/Y sky130_fd_sc_hd__inv_2
X_5407_ _5407_/A VGND VGND VPWR VPWR _5408_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_133_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9175_ _9679_/CLK _9175_/D _9730_/SET_B VGND VGND VPWR VPWR _9175_/Q sky130_fd_sc_hd__dfrtp_1
X_8126_ _8126_/A _8580_/D VGND VGND VPWR VPWR _8127_/B sky130_fd_sc_hd__or2_1
X_5338_ _9545_/Q _5331_/A hold593/X _5331_/Y VGND VGND VPWR VPWR _9545_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8057_ _8068_/A _8443_/A VGND VGND VPWR VPWR _8059_/C sky130_fd_sc_hd__or2_1
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7008_ _6176_/Y _7007_/A _9061_/Q _7007_/Y VGND VGND VPWR VPWR _9061_/D sky130_fd_sc_hd__o22a_1
XFILLER_125_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5269_ _9592_/Q _5265_/A _8959_/A1 _5265_/Y VGND VGND VPWR VPWR _9592_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8959_ _9664_/Q _8959_/A1 _8973_/S VGND VGND VPWR VPWR _8959_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4640_ _9764_/Q hold673/X _6067_/B1 _4636_/Y VGND VGND VPWR VPWR _9764_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4571_ _4572_/B VGND VGND VPWR VPWR _5085_/D sky130_fd_sc_hd__clkinv_4
X_6310_ _6305_/Y _5406_/B _6306_/Y _4869_/X _6309_/X VGND VGND VPWR VPWR _6311_/D
+ sky130_fd_sc_hd__o221a_4
X_7290_ _6202_/Y _7173_/X _6236_/Y _7174_/X VGND VGND VPWR VPWR _7290_/X sky130_fd_sc_hd__o22a_1
Xhold705 _9191_/Q VGND VGND VPWR VPWR hold705/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_115_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6241_ _6236_/Y _5532_/B _6237_/Y _6117_/X _6240_/X VGND VGND VPWR VPWR _6242_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_170_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6172_ _9369_/Q VGND VGND VPWR VPWR _6172_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5123_ _5282_/A _5123_/B VGND VGND VPWR VPWR _5123_/X sky130_fd_sc_hd__or2_1
XFILLER_57_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5054_ _9725_/Q _5049_/A _6008_/B1 _5049_/Y VGND VGND VPWR VPWR _5054_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8813_ _8813_/A VGND VGND VPWR VPWR _8814_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_65_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9793_ _9798_/CLK _9793_/D _9821_/SET_B VGND VGND VPWR VPWR _9793_/Q sky130_fd_sc_hd__dfstp_1
X_5956_ _7805_/A _7805_/B _7803_/A _7803_/B VGND VGND VPWR VPWR _5966_/B sky130_fd_sc_hd__or4_1
X_8744_ _8774_/A _8777_/C VGND VGND VPWR VPWR _8744_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8675_ _8675_/A _8751_/C _8730_/C _8729_/C VGND VGND VPWR VPWR _8675_/Y sky130_fd_sc_hd__nor4_1
X_5887_ _5878_/X _8898_/X _8960_/X _9210_/Q VGND VGND VPWR VPWR _9210_/D sky130_fd_sc_hd__o22a_1
X_4907_ _6189_/A _6117_/B input34/X VGND VGND VPWR VPWR _4907_/X sky130_fd_sc_hd__or3b_1
XFILLER_166_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7626_ _6157_/Y _7491_/X _6151_/Y _7492_/X _7625_/X VGND VGND VPWR VPWR _7640_/B
+ sky130_fd_sc_hd__o221a_1
X_4838_ _9484_/Q VGND VGND VPWR VPWR _4838_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7557_ _7733_/A _7500_/X _8827_/A _7501_/X _7556_/X VGND VGND VPWR VPWR _7557_/X
+ sky130_fd_sc_hd__o221a_1
X_4769_ _4747_/Y _5687_/B _4752_/X _4757_/X _4768_/X VGND VGND VPWR VPWR _4812_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_119_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7488_ _7488_/A VGND VGND VPWR VPWR _7488_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6508_ _9271_/Q VGND VGND VPWR VPWR _6508_/Y sky130_fd_sc_hd__inv_2
X_9227_ _9679_/CLK _9227_/D _9730_/SET_B VGND VGND VPWR VPWR _9227_/Q sky130_fd_sc_hd__dfrtp_1
X_6439_ _6439_/A _6439_/B _6439_/C _6439_/D VGND VGND VPWR VPWR _6505_/A sky130_fd_sc_hd__and4_2
X_9158_ _9679_/CLK _9158_/D _9730_/SET_B VGND VGND VPWR VPWR _9158_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8109_ _8557_/A _8205_/A VGND VGND VPWR VPWR _8244_/A sky130_fd_sc_hd__or2_1
XFILLER_121_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold10 hold9/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__dlygate4sd3_1
X_9089_ _9832_/CLK _9089_/D VGND VGND VPWR VPWR _9089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold43 hold43/A VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold54 hold54/A VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold87 hold87/A VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_7 _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5810_ _9265_/Q _5807_/A hold696/X _5807_/Y VGND VGND VPWR VPWR _9265_/D sky130_fd_sc_hd__a22o_1
X_6790_ _6790_/A _6790_/B _6790_/C VGND VGND VPWR VPWR _6815_/C sky130_fd_sc_hd__and3_1
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5741_ _5741_/A VGND VGND VPWR VPWR _5741_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_175_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8460_ _8728_/A VGND VGND VPWR VPWR _8460_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5672_ _9320_/Q VGND VGND VPWR VPWR _5780_/C sky130_fd_sc_hd__inv_2
X_7411_ _6495_/Y _7067_/A _6362_/Y _7146_/A VGND VGND VPWR VPWR _7411_/X sky130_fd_sc_hd__o22a_1
X_8391_ _8682_/A _8391_/B VGND VGND VPWR VPWR _8394_/B sky130_fd_sc_hd__or2_2
X_4623_ _5201_/A _4623_/B VGND VGND VPWR VPWR _4624_/A sky130_fd_sc_hd__or2_1
X_7342_ _6904_/Y _7139_/X _6898_/Y _7140_/X VGND VGND VPWR VPWR _7342_/X sky130_fd_sc_hd__o22a_1
X_4554_ _9805_/Q _4547_/A _6067_/B1 _4547_/Y VGND VGND VPWR VPWR _9805_/D sky130_fd_sc_hd__a22o_1
Xhold502 _9131_/Q VGND VGND VPWR VPWR hold503/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _5305_/X VGND VGND VPWR VPWR _9568_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold524 _5496_/X VGND VGND VPWR VPWR _9439_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold535 _5333_/X VGND VGND VPWR VPWR _9550_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7273_ _6300_/Y _7180_/X _6342_/Y _7181_/X _7272_/X VGND VGND VPWR VPWR _7274_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6224_ _6224_/A VGND VGND VPWR VPWR _6224_/Y sky130_fd_sc_hd__inv_2
Xhold546 _5183_/X VGND VGND VPWR VPWR _9650_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold579 hold704/X VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold568 _5601_/X VGND VGND VPWR VPWR _9369_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold557 _5382_/X VGND VGND VPWR VPWR _9516_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_9012_ _8530_/X _8380_/X _9017_/S VGND VGND VPWR VPWR _9012_/X sky130_fd_sc_hd__mux2_1
X_4485_ _4485_/A VGND VGND VPWR VPWR _4485_/Y sky130_fd_sc_hd__clkinv_2
X_6155_ _6153_/Y _5786_/B _6154_/Y _5935_/B VGND VGND VPWR VPWR _6155_/X sky130_fd_sc_hd__o22a_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _9089_/Q _6085_/A _8964_/A1 _6085_/Y VGND VGND VPWR VPWR _9089_/D sky130_fd_sc_hd__a22o_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5106_ _9700_/Q _5105_/A _8959_/A1 _5105_/Y VGND VGND VPWR VPWR _9700_/D sky130_fd_sc_hd__a22o_1
X_5037_ _5037_/A VGND VGND VPWR VPWR _5038_/A sky130_fd_sc_hd__buf_4
Xrepeater396 hold136/X VGND VGND VPWR VPWR hold217/A sky130_fd_sc_hd__buf_12
XFILLER_26_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9776_ _9819_/CLK _9776_/D _9821_/SET_B VGND VGND VPWR VPWR _9776_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6988_ _6660_/Y _6983_/A _9073_/Q _6983_/Y VGND VGND VPWR VPWR _9073_/D sky130_fd_sc_hd__o22a_1
X_8727_ _8727_/A _8727_/B VGND VGND VPWR VPWR _8728_/B sky130_fd_sc_hd__or2_1
XFILLER_40_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5939_ _9173_/Q _5937_/A hold510/X _5937_/Y VGND VGND VPWR VPWR _9173_/D sky130_fd_sc_hd__a22o_1
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8658_ _8777_/A _8658_/B _8710_/D _8741_/C VGND VGND VPWR VPWR _8661_/A sky130_fd_sc_hd__or4_2
XFILLER_21_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7609_ _6231_/Y _7498_/X _6207_/Y _5727_/X VGND VGND VPWR VPWR _7609_/X sky130_fd_sc_hd__o22a_1
X_8589_ _8139_/A _8588_/Y _8440_/Y VGND VGND VPWR VPWR _8589_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput111 sram_ro_data[26] VGND VGND VPWR VPWR _6700_/A sky130_fd_sc_hd__clkbuf_1
Xinput100 sram_ro_data[16] VGND VGND VPWR VPWR _4862_/A sky130_fd_sc_hd__clkbuf_1
Xinput144 wb_adr_i[20] VGND VGND VPWR VPWR _7874_/B sky130_fd_sc_hd__buf_2
Xinput133 wb_adr_i[10] VGND VGND VPWR VPWR _7806_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_163_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput122 sram_ro_data[7] VGND VGND VPWR VPWR _6106_/A sky130_fd_sc_hd__clkbuf_1
Xinput177 wb_dat_i[20] VGND VGND VPWR VPWR _7776_/B sky130_fd_sc_hd__clkbuf_1
Xinput166 wb_dat_i[10] VGND VGND VPWR VPWR _7773_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_adr_i[30] VGND VGND VPWR VPWR _5961_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput199 wb_sel_i[1] VGND VGND VPWR VPWR _5081_/B sky130_fd_sc_hd__clkbuf_1
Xinput188 wb_dat_i[30] VGND VGND VPWR VPWR _7781_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7960_ _8118_/A _8304_/B _7959_/X VGND VGND VPWR VPWR _7960_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6911_ _9337_/Q VGND VGND VPWR VPWR _7178_/A sky130_fd_sc_hd__clkinv_2
XFILLER_94_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7891_ _7891_/A VGND VGND VPWR VPWR _8312_/B sky130_fd_sc_hd__buf_2
X_9630_ _9643_/CLK _9630_/D _9563_/SET_B VGND VGND VPWR VPWR _9630_/Q sky130_fd_sc_hd__dfrtp_1
X_6842_ _9764_/Q VGND VGND VPWR VPWR _6842_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6773_ _9676_/Q VGND VGND VPWR VPWR _6773_/Y sky130_fd_sc_hd__inv_2
X_9561_ _9561_/CLK _9561_/D _9817_/SET_B VGND VGND VPWR VPWR _9561_/Q sky130_fd_sc_hd__dfrtp_1
X_9492_ _9569_/CLK _9492_/D _9563_/SET_B VGND VGND VPWR VPWR _9492_/Q sky130_fd_sc_hd__dfstp_1
X_8512_ _8512_/A _8512_/B _8740_/A VGND VGND VPWR VPWR _8516_/A sky130_fd_sc_hd__or3_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5724_ _9297_/Q VGND VGND VPWR VPWR _7478_/D sky130_fd_sc_hd__inv_2
X_5655_ _9330_/Q _5649_/A _8965_/A1 _5649_/Y VGND VGND VPWR VPWR _5655_/X sky130_fd_sc_hd__a22o_1
X_8443_ _8443_/A _8443_/B VGND VGND VPWR VPWR _8443_/X sky130_fd_sc_hd__or2_1
XFILLER_191_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8374_ _8341_/A _8324_/C _8324_/B _8373_/X VGND VGND VPWR VPWR _8375_/C sky130_fd_sc_hd__a31o_1
X_4606_ _9784_/Q _4600_/A hold217/X _4600_/Y VGND VGND VPWR VPWR _9784_/D sky130_fd_sc_hd__a22o_1
Xhold310 hold310/A VGND VGND VPWR VPWR hold311/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7325_ _4952_/Y _7151_/X _4905_/Y _7152_/X VGND VGND VPWR VPWR _7325_/X sky130_fd_sc_hd__o22a_1
X_5586_ _9377_/Q _5583_/A hold217/X _5583_/Y VGND VGND VPWR VPWR _9377_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold321 _5537_/X VGND VGND VPWR VPWR hold322/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 hold332/A VGND VGND VPWR VPWR _9316_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold343 hold343/A VGND VGND VPWR VPWR hold344/A sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ _4537_/A VGND VGND VPWR VPWR _4537_/Y sky130_fd_sc_hd__inv_2
Xhold376 hold376/A VGND VGND VPWR VPWR _9635_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7256_ _6275_/Y _7135_/X _6287_/Y _7136_/X _7255_/X VGND VGND VPWR VPWR _7275_/A
+ sky130_fd_sc_hd__o221a_1
Xhold387 hold387/A VGND VGND VPWR VPWR hold388/A sky130_fd_sc_hd__dlygate4sd3_1
X_4468_ _9612_/Q hold23/A _9122_/Q VGND VGND VPWR VPWR _9027_/A sky130_fd_sc_hd__mux2_1
Xhold354 hold354/A VGND VGND VPWR VPWR _4920_/A sky130_fd_sc_hd__buf_2
Xhold365 hold365/A VGND VGND VPWR VPWR _4823_/B sky130_fd_sc_hd__clkbuf_2
X_6207_ _9368_/Q VGND VGND VPWR VPWR _6207_/Y sky130_fd_sc_hd__inv_2
X_7187_ _7187_/A _7187_/B _7187_/C VGND VGND VPWR VPWR _7187_/Y sky130_fd_sc_hd__nand3_4
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold398 hold398/A VGND VGND VPWR VPWR _4750_/C sky130_fd_sc_hd__buf_2
X_6138_ _6136_/Y _5133_/B _6137_/Y _4844_/X VGND VGND VPWR VPWR _6138_/X sky130_fd_sc_hd__o22a_4
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _9111_/Q _4485_/A _8964_/A1 _4485_/Y VGND VGND VPWR VPWR _9111_/D sky130_fd_sc_hd__a22o_1
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9828_ _9830_/CLK _9828_/D _9537_/SET_B VGND VGND VPWR VPWR _9828_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9759_ net399_3/A _9759_/D _4660_/X VGND VGND VPWR VPWR _9759_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_41_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5440_ _9477_/Q _5438_/A _6065_/B1 _5438_/Y VGND VGND VPWR VPWR _9477_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5371_ _9524_/Q _5369_/A hold510/X _5369_/Y VGND VGND VPWR VPWR _5371_/X sky130_fd_sc_hd__a22o_1
XFILLER_126_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8090_ _8138_/B _8596_/A _8089_/Y VGND VGND VPWR VPWR _8094_/A sky130_fd_sc_hd__o21ba_1
X_7110_ _4919_/Y _7149_/A _4800_/Y _7150_/A _7109_/X VGND VGND VPWR VPWR _7116_/B
+ sky130_fd_sc_hd__o221a_1
X_7041_ _9668_/Q _7042_/B VGND VGND VPWR VPWR _7041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_opt_1_1_wb_clk_i clkbuf_opt_1_1_wb_clk_i/A VGND VGND VPWR VPWR _9064_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_8992_ _9756_/Q _6506_/Y _8999_/S VGND VGND VPWR VPWR _8992_/X sky130_fd_sc_hd__mux2_1
X_7943_ _7943_/A VGND VGND VPWR VPWR _8540_/A sky130_fd_sc_hd__clkbuf_4
X_7874_ _7874_/A _7874_/B _7874_/C VGND VGND VPWR VPWR _7918_/A sky130_fd_sc_hd__or3_4
XFILLER_63_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _9705_/CLK sky130_fd_sc_hd__clkbuf_2
X_9613_ _9731_/CLK _9613_/D _9731_/SET_B VGND VGND VPWR VPWR _9613_/Q sky130_fd_sc_hd__dfrtp_1
X_6825_ _6825_/A VGND VGND VPWR VPWR _6825_/Y sky130_fd_sc_hd__inv_2
X_9544_ _9577_/CLK _9544_/D _9571_/SET_B VGND VGND VPWR VPWR _9544_/Q sky130_fd_sc_hd__dfstp_1
X_6756_ _9598_/Q VGND VGND VPWR VPWR _6756_/Y sky130_fd_sc_hd__inv_2
X_5707_ _5707_/A VGND VGND VPWR VPWR _5708_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9475_ _9483_/CLK _9475_/D _9727_/SET_B VGND VGND VPWR VPWR _9475_/Q sky130_fd_sc_hd__dfrtp_1
X_6687_ _9806_/Q VGND VGND VPWR VPWR _6687_/Y sky130_fd_sc_hd__inv_2
X_5638_ _5638_/A VGND VGND VPWR VPWR _5638_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8426_ _8426_/A _8693_/B VGND VGND VPWR VPWR _8427_/B sky130_fd_sc_hd__nor2_1
X_5569_ _9388_/Q _5561_/A hold601/X _5561_/Y VGND VGND VPWR VPWR _5569_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8357_ _8280_/A _8540_/B _8346_/Y _8355_/X _8356_/X VGND VGND VPWR VPWR _8360_/A
+ sky130_fd_sc_hd__o2111ai_4
Xhold151 hold151/A VGND VGND VPWR VPWR _9390_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold140 _5375_/X VGND VGND VPWR VPWR hold141/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 hold162/A VGND VGND VPWR VPWR hold163/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7308_ _6152_/Y _7160_/X _6093_/Y _7071_/B _7307_/X VGND VGND VPWR VPWR _7309_/D
+ sky130_fd_sc_hd__o221a_1
Xhold173 _9701_/Q VGND VGND VPWR VPWR hold174/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 hold195/A VGND VGND VPWR VPWR hold196/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 hold184/A VGND VGND VPWR VPWR _9466_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_78_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8288_ _8288_/A _8288_/B VGND VGND VPWR VPWR _8532_/B sky130_fd_sc_hd__nor2_1
XFILLER_132_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7239_ _6459_/Y _7095_/B _6408_/Y _7157_/X VGND VGND VPWR VPWR _7239_/X sky130_fd_sc_hd__o22a_1
XFILLER_77_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4940_ _9427_/Q VGND VGND VPWR VPWR _4940_/Y sky130_fd_sc_hd__clkinv_2
X_4871_ _6142_/B _4951_/B VGND VGND VPWR VPWR _5466_/B sky130_fd_sc_hd__or2_4
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7590_ _6332_/Y _7491_/X _6328_/Y _7492_/X _7589_/X VGND VGND VPWR VPWR _7604_/B
+ sky130_fd_sc_hd__o221a_1
X_6610_ _6605_/Y _5321_/B _8809_/A _5521_/B _6609_/X VGND VGND VPWR VPWR _6617_/B
+ sky130_fd_sc_hd__o221a_1
X_6541_ _9309_/Q VGND VGND VPWR VPWR _6541_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_32_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9260_ _9734_/CLK _9260_/D _9731_/SET_B VGND VGND VPWR VPWR _9260_/Q sky130_fd_sc_hd__dfstp_1
X_6472_ _9179_/Q VGND VGND VPWR VPWR _6472_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8211_ _8211_/A _8431_/A VGND VGND VPWR VPWR _8438_/A sky130_fd_sc_hd__or2_1
X_5423_ _9488_/Q _5419_/A _8959_/A1 _5419_/Y VGND VGND VPWR VPWR _9488_/D sky130_fd_sc_hd__a22o_1
X_9191_ _9319_/CLK _9191_/D _9797_/SET_B VGND VGND VPWR VPWR _9191_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput234 _8842_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_2
Xoutput223 _8822_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_2
X_8142_ _8255_/A VGND VGND VPWR VPWR _8243_/B sky130_fd_sc_hd__buf_8
Xoutput212 _8802_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_2
X_5354_ _9535_/Q _5353_/A _6064_/B1 _5353_/Y VGND VGND VPWR VPWR _9535_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput245 _8866_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_2
Xoutput256 _8869_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_2
Xoutput267 _9021_/Z VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_141_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8073_ _8563_/A _8593_/A VGND VGND VPWR VPWR _8656_/B sky130_fd_sc_hd__nor2_1
Xoutput278 _9024_/Z VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_2
Xoutput289 _7045_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_2
X_5285_ _9582_/Q _5284_/A _6064_/B1 _5284_/Y VGND VGND VPWR VPWR _9582_/D sky130_fd_sc_hd__a22o_1
X_7024_ _9096_/Q _8861_/X _9096_/Q _7028_/C _9097_/Q VGND VGND VPWR VPWR _9096_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_59_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8975_ _9644_/Q _8975_/A1 _8975_/S VGND VGND VPWR VPWR _8975_/X sky130_fd_sc_hd__mux2_1
X_7926_ _7873_/B _7918_/Y _7925_/X VGND VGND VPWR VPWR _7926_/Y sky130_fd_sc_hd__o21ai_2
X_7857_ _8702_/B VGND VGND VPWR VPWR _8324_/B sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_4_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9728_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6808_ _6803_/Y _5971_/B _6804_/Y _5112_/B _6807_/X VGND VGND VPWR VPWR _6814_/C
+ sky130_fd_sc_hd__o221a_1
X_7788_ _8702_/A VGND VGND VPWR VPWR _8341_/A sky130_fd_sc_hd__inv_2
X_6739_ _6737_/Y _4892_/X _6738_/Y _5628_/B VGND VGND VPWR VPWR _6739_/X sky130_fd_sc_hd__o22a_1
X_9527_ _9800_/CLK _9527_/D _9817_/SET_B VGND VGND VPWR VPWR _9527_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9458_ _9516_/CLK _9458_/D _9571_/SET_B VGND VGND VPWR VPWR _9458_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_136_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8409_ _8409_/A _8409_/B VGND VGND VPWR VPWR _8620_/C sky130_fd_sc_hd__or2_1
XFILLER_3_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9389_ _9391_/CLK _9389_/D _9689_/SET_B VGND VGND VPWR VPWR _9389_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_136_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5070_ _5070_/A VGND VGND VPWR VPWR _5070_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8760_ _8389_/X _8759_/X _8265_/B _8354_/D VGND VGND VPWR VPWR _8761_/B sky130_fd_sc_hd__o211ai_1
XFILLER_92_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5972_ _5972_/A VGND VGND VPWR VPWR _5973_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4923_ _4923_/A VGND VGND VPWR VPWR _4923_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7711_ _7711_/A _7711_/B _7711_/C _7711_/D VGND VGND VPWR VPWR _7712_/D sky130_fd_sc_hd__and4_1
XFILLER_52_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8691_ _8764_/A _8723_/B _8762_/B VGND VGND VPWR VPWR _8691_/Y sky130_fd_sc_hd__nor3_1
XFILLER_33_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4854_ _4883_/A _6117_/B VGND VGND VPWR VPWR _4854_/X sky130_fd_sc_hd__or2_4
X_7642_ _4942_/Y _7485_/X _4752_/A _7486_/X _7641_/X VGND VGND VPWR VPWR _7658_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7573_ _6453_/Y _7498_/X _6391_/Y _5727_/X VGND VGND VPWR VPWR _7573_/X sky130_fd_sc_hd__o22a_1
X_4785_ _4808_/A _6142_/B VGND VGND VPWR VPWR _5589_/B sky130_fd_sc_hd__or2_4
X_9312_ _9318_/CLK _9312_/D _9571_/SET_B VGND VGND VPWR VPWR _9312_/Q sky130_fd_sc_hd__dfstp_1
X_6524_ _6522_/Y _5570_/B _8793_/A _5826_/B VGND VGND VPWR VPWR _6524_/X sky130_fd_sc_hd__o22a_1
XFILLER_118_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9243_ _9600_/CLK _9243_/D _9797_/SET_B VGND VGND VPWR VPWR _9243_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6455_ _9405_/Q VGND VGND VPWR VPWR _6455_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_161_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9174_ _9830_/CLK _9174_/D _9537_/SET_B VGND VGND VPWR VPWR _9174_/Q sky130_fd_sc_hd__dfrtp_1
X_5406_ _5570_/A _5406_/B VGND VGND VPWR VPWR _5407_/A sky130_fd_sc_hd__or2_2
X_6386_ _6385_/Y _5144_/B _4866_/X _6189_/X VGND VGND VPWR VPWR _6386_/X sky130_fd_sc_hd__o211a_1
X_5337_ _9546_/Q _5331_/A hold136/X _5331_/Y VGND VGND VPWR VPWR _5337_/X sky130_fd_sc_hd__a22o_1
X_8125_ _8125_/A _8563_/B VGND VGND VPWR VPWR _8580_/D sky130_fd_sc_hd__or2_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8056_ _8056_/A _8056_/B _8056_/C _8056_/D VGND VGND VPWR VPWR _8056_/X sky130_fd_sc_hd__or4_1
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5268_ _9593_/Q _5265_/A hold696/A _5265_/Y VGND VGND VPWR VPWR _9593_/D sky130_fd_sc_hd__a22o_1
X_7007_ _7007_/A VGND VGND VPWR VPWR _7007_/Y sky130_fd_sc_hd__inv_2
X_5199_ _9637_/Q _5192_/A hold593/X _5192_/Y VGND VGND VPWR VPWR _9637_/D sky130_fd_sc_hd__a22o_1
X_8958_ _9651_/Q hold516/X _8975_/S VGND VGND VPWR VPWR _8958_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7909_ _7909_/A VGND VGND VPWR VPWR _8288_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8889_ _7053_/Y _9682_/Q _9629_/Q VGND VGND VPWR VPWR _8889_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4570_ _8853_/A _9017_/S VGND VGND VPWR VPWR _4572_/B sky130_fd_sc_hd__nand2_8
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold706 _9213_/Q VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6240_ _6238_/Y _4844_/X _6239_/Y _4929_/X VGND VGND VPWR VPWR _6240_/X sky130_fd_sc_hd__o22a_4
XFILLER_170_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6171_ _9239_/Q VGND VGND VPWR VPWR _6171_/Y sky130_fd_sc_hd__clkinv_2
X_5122_ _9688_/Q _5114_/A _8975_/A1 _5114_/Y VGND VGND VPWR VPWR _9688_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5053_ _9726_/Q _5049_/A _6067_/B1 _5049_/Y VGND VGND VPWR VPWR _9726_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8812_ _8812_/A VGND VGND VPWR VPWR _8812_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9792_ _9798_/CLK _9792_/D _9821_/SET_B VGND VGND VPWR VPWR _9792_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5955_ _7803_/C _7803_/D _5955_/C input149/X VGND VGND VPWR VPWR _5966_/A sky130_fd_sc_hd__or4b_1
X_8743_ _8105_/C _8742_/Y _8056_/C _8569_/C _8655_/B VGND VGND VPWR VPWR _8777_/C
+ sky130_fd_sc_hd__a2111o_2
X_8674_ _8674_/A _8674_/B VGND VGND VPWR VPWR _8729_/C sky130_fd_sc_hd__nor2_1
X_5886_ _5878_/X _8900_/X _8960_/X _9211_/Q VGND VGND VPWR VPWR _9211_/D sky130_fd_sc_hd__o22a_1
X_4906_ _4933_/A _6142_/B VGND VGND VPWR VPWR _5282_/B sky130_fd_sc_hd__or2_4
XFILLER_33_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7625_ _6160_/Y _7493_/X _6147_/Y _7494_/X VGND VGND VPWR VPWR _7625_/X sky130_fd_sc_hd__o22a_1
X_4837_ _4913_/B _6189_/B VGND VGND VPWR VPWR _6058_/B sky130_fd_sc_hd__or2_4
XFILLER_193_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7556_ _8821_/A _7502_/X _8819_/A _7503_/X VGND VGND VPWR VPWR _7556_/X sky130_fd_sc_hd__o22a_1
X_4768_ _4758_/Y _6165_/A _4761_/Y _5847_/B _4767_/X VGND VGND VPWR VPWR _4768_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6507_ _6180_/A _6506_/Y _9082_/Q _6180_/Y VGND VGND VPWR VPWR _9082_/D sky130_fd_sc_hd__o22a_2
XFILLER_174_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4699_ _4803_/A _4947_/A VGND VGND VPWR VPWR _5201_/B sky130_fd_sc_hd__or2_4
X_7487_ _7487_/A VGND VGND VPWR VPWR _7487_/X sky130_fd_sc_hd__clkbuf_8
X_9226_ _9421_/CLK _9226_/D _9537_/SET_B VGND VGND VPWR VPWR _9226_/Q sky130_fd_sc_hd__dfrtp_1
X_6438_ _6433_/Y _5263_/B _6434_/Y _4511_/B _6437_/X VGND VGND VPWR VPWR _6439_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_106_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9157_ _9730_/CLK _9157_/D _9730_/SET_B VGND VGND VPWR VPWR _9157_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_22_csclk clkbuf_opt_4_0_csclk/X VGND VGND VPWR VPWR _9651_/CLK sky130_fd_sc_hd__clkbuf_16
X_8108_ _8108_/A _8581_/A VGND VGND VPWR VPWR _8110_/A sky130_fd_sc_hd__nor2_1
XFILLER_121_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6369_ _6367_/Y _4915_/X _6368_/Y _5935_/B VGND VGND VPWR VPWR _6369_/X sky130_fd_sc_hd__o22a_1
XFILLER_102_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 hold11/A VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_9088_ _9832_/CLK _9088_/D VGND VGND VPWR VPWR _9088_/Q sky130_fd_sc_hd__dfxtp_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__dlygate4sd3_1
X_8039_ _8157_/B _8091_/B VGND VGND VPWR VPWR _8040_/A sky130_fd_sc_hd__or2_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9827_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_8 _4772_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5740_ _5723_/A _5732_/Y _5738_/Y _9294_/Q _5741_/A VGND VGND VPWR VPWR _9294_/D
+ sky130_fd_sc_hd__o32a_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _7028_/A _5669_/Y _5752_/B _9096_/Q _8861_/X VGND VGND VPWR VPWR _5685_/A
+ sky130_fd_sc_hd__a32o_1
X_7410_ _6428_/Y _7135_/A _6418_/Y _7136_/A _7409_/X VGND VGND VPWR VPWR _7429_/A
+ sky130_fd_sc_hd__o221a_1
X_8390_ _8420_/B _8389_/X _8258_/X VGND VGND VPWR VPWR _8391_/B sky130_fd_sc_hd__o21a_1
X_4622_ _6142_/A _4943_/A VGND VGND VPWR VPWR _4623_/B sky130_fd_sc_hd__or2_4
XFILLER_156_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4553_ _9806_/Q _4547_/A hold217/X _4547_/Y VGND VGND VPWR VPWR _9806_/D sky130_fd_sc_hd__a22o_1
X_7341_ _7341_/A _7341_/B _7341_/C VGND VGND VPWR VPWR _7341_/Y sky130_fd_sc_hd__nand3_2
Xhold525 _5535_/X VGND VGND VPWR VPWR _9413_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold514 _9708_/Q VGND VGND VPWR VPWR hold515/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 _5458_/X VGND VGND VPWR VPWR _9465_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7272_ _6322_/Y _7182_/X _6272_/Y _7183_/X VGND VGND VPWR VPWR _7272_/X sky130_fd_sc_hd__o22a_1
X_4484_ _4484_/A VGND VGND VPWR VPWR _4485_/A sky130_fd_sc_hd__buf_2
Xhold503 hold503/A VGND VGND VPWR VPWR hold504/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 _8957_/X VGND VGND VPWR VPWR hold569/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_9011_ _8338_/Y _7983_/X _9017_/S VGND VGND VPWR VPWR _9011_/X sky130_fd_sc_hd__mux2_1
Xhold547 _5332_/X VGND VGND VPWR VPWR _9551_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold558 _6061_/X VGND VGND VPWR VPWR _9119_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6223_ _6219_/Y _6058_/B _6220_/Y _4511_/B _6222_/X VGND VGND VPWR VPWR _6242_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_103_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6154_ _9174_/Q VGND VGND VPWR VPWR _6154_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5105_ _5105_/A VGND VGND VPWR VPWR _5105_/Y sky130_fd_sc_hd__inv_2
X_6085_ _6085_/A VGND VGND VPWR VPWR _6085_/Y sky130_fd_sc_hd__inv_2
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5201_/A _5036_/B VGND VGND VPWR VPWR _5037_/A sky130_fd_sc_hd__or2_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater397 hold136/X VGND VGND VPWR VPWR _8965_/A1 sky130_fd_sc_hd__buf_12
X_6987_ _6506_/Y _6983_/A _9074_/Q _6983_/Y VGND VGND VPWR VPWR _9074_/D sky130_fd_sc_hd__o22a_2
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9775_ _9817_/CLK _9775_/D _9817_/SET_B VGND VGND VPWR VPWR _9775_/Q sky130_fd_sc_hd__dfstp_1
X_5938_ _9174_/Q _5937_/A hold516/X _5937_/Y VGND VGND VPWR VPWR _5938_/X sky130_fd_sc_hd__a22o_1
X_8726_ _8156_/Y _8667_/B _8447_/A _8725_/X _8671_/B VGND VGND VPWR VPWR _8731_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5869_ _9226_/Q _5868_/A hold516/X _5868_/Y VGND VGND VPWR VPWR _5869_/X sky130_fd_sc_hd__a22o_1
X_8657_ _8657_/A _8657_/B _8657_/C _8657_/D VGND VGND VPWR VPWR _8741_/C sky130_fd_sc_hd__or4_1
X_8588_ _8588_/A _8608_/B VGND VGND VPWR VPWR _8588_/Y sky130_fd_sc_hd__nor2_1
X_7608_ _6213_/Y _7491_/X _6246_/Y _7492_/X _7607_/X VGND VGND VPWR VPWR _7622_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7539_ _6785_/Y _7500_/X _6792_/Y _7501_/X _7538_/X VGND VGND VPWR VPWR _7539_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9209_ _9212_/CLK _9209_/D _9797_/SET_B VGND VGND VPWR VPWR _9209_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput101 sram_ro_data[17] VGND VGND VPWR VPWR _6837_/A sky130_fd_sc_hd__clkbuf_1
Xinput145 wb_adr_i[21] VGND VGND VPWR VPWR _7869_/A sky130_fd_sc_hd__buf_2
Xinput134 wb_adr_i[11] VGND VGND VPWR VPWR _7806_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_163_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput112 sram_ro_data[27] VGND VGND VPWR VPWR _6592_/A sky130_fd_sc_hd__clkbuf_1
Xinput123 sram_ro_data[8] VGND VGND VPWR VPWR _4914_/A sky130_fd_sc_hd__clkbuf_1
Xinput178 wb_dat_i[21] VGND VGND VPWR VPWR _7778_/B sky130_fd_sc_hd__clkbuf_1
Xinput167 wb_dat_i[11] VGND VGND VPWR VPWR _7775_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput156 wb_adr_i[31] VGND VGND VPWR VPWR _5961_/A sky130_fd_sc_hd__clkbuf_1
Xinput189 wb_dat_i[31] VGND VGND VPWR VPWR _7783_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6910_ _9247_/Q VGND VGND VPWR VPWR _6910_/Y sky130_fd_sc_hd__clkinv_2
X_7890_ _8366_/A _8489_/A VGND VGND VPWR VPWR _7891_/A sky130_fd_sc_hd__or2_1
XFILLER_54_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6841_ _6836_/Y _5255_/B _6837_/Y _4863_/X _6840_/X VGND VGND VPWR VPWR _6860_/A
+ sky130_fd_sc_hd__o221a_1
X_9560_ _9686_/CLK _9560_/D _7042_/B VGND VGND VPWR VPWR _9560_/Q sky130_fd_sc_hd__dfrtp_1
X_8511_ _7887_/A _8229_/A _8138_/B _8596_/A VGND VGND VPWR VPWR _8740_/A sky130_fd_sc_hd__o22ai_1
X_6772_ _6772_/A _6772_/B _6772_/C _6772_/D VGND VGND VPWR VPWR _6815_/B sky130_fd_sc_hd__and4_1
XFILLER_188_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9491_ _9491_/CLK _9491_/D _9731_/SET_B VGND VGND VPWR VPWR _9491_/Q sky130_fd_sc_hd__dfrtp_1
X_5723_ _5723_/A _7471_/A _7467_/A VGND VGND VPWR VPWR _5723_/Y sky130_fd_sc_hd__nor3_1
X_5654_ _9331_/Q _5649_/A hold42/X _5649_/Y VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__a22o_1
XFILLER_148_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8442_ _8563_/A _8158_/A _8435_/Y _8443_/B _8441_/X VGND VGND VPWR VPWR _8442_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_175_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8373_ _8373_/A _8373_/B VGND VGND VPWR VPWR _8373_/X sky130_fd_sc_hd__or2_1
X_4605_ _9785_/Q _4600_/A _6065_/B1 _4600_/Y VGND VGND VPWR VPWR _9785_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold300 _5372_/X VGND VGND VPWR VPWR hold301/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 hold311/A VGND VGND VPWR VPWR _9278_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7324_ _4782_/Y _7144_/X _4805_/Y _7145_/X _7323_/X VGND VGND VPWR VPWR _7331_/A
+ sky130_fd_sc_hd__o221a_1
X_5585_ _9378_/Q _5583_/A _6065_/B1 _5583_/Y VGND VGND VPWR VPWR _9378_/D sky130_fd_sc_hd__a22o_1
Xhold322 hold322/A VGND VGND VPWR VPWR hold323/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _5526_/X VGND VGND VPWR VPWR hold334/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold344 hold344/A VGND VGND VPWR VPWR _4473_/A sky130_fd_sc_hd__buf_6
X_4536_ _4920_/A _4643_/A VGND VGND VPWR VPWR _4536_/X sky130_fd_sc_hd__or2_2
Xhold377 _8956_/X VGND VGND VPWR VPWR hold378/A sky130_fd_sc_hd__dlygate4sd3_1
X_7255_ _6340_/Y _7137_/X _6318_/Y _7138_/X _7254_/X VGND VGND VPWR VPWR _7255_/X
+ sky130_fd_sc_hd__o221a_1
Xhold366 _9719_/Q VGND VGND VPWR VPWR hold367/A sky130_fd_sc_hd__dlygate4sd3_1
X_4467_ _9613_/Q _4467_/A1 _9724_/Q VGND VGND VPWR VPWR _9028_/A sky130_fd_sc_hd__mux2_1
Xhold355 _8987_/X VGND VGND VPWR VPWR hold625/A sky130_fd_sc_hd__dlygate4sd3_1
X_6206_ _9238_/Q VGND VGND VPWR VPWR _6206_/Y sky130_fd_sc_hd__clkinv_2
X_7186_ _7186_/A _7186_/B _7186_/C _7186_/D VGND VGND VPWR VPWR _7187_/C sky130_fd_sc_hd__and4_1
Xhold388 hold388/A VGND VGND VPWR VPWR _9397_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold399 _4866_/A VGND VGND VPWR VPWR hold400/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6137_ _6137_/A VGND VGND VPWR VPWR _6137_/Y sky130_fd_sc_hd__inv_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6068_ _9112_/Q _6060_/A hold601/A _6060_/Y VGND VGND VPWR VPWR _6068_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5019_ _8954_/X _9741_/Q _5024_/S VGND VGND VPWR VPWR _5020_/A sky130_fd_sc_hd__mux2_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9827_ _9827_/CLK _9827_/D _9797_/SET_B VGND VGND VPWR VPWR _9827_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_26_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9758_ net399_3/A _9758_/D _4663_/X VGND VGND VPWR VPWR _9758_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_186_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9689_ _9694_/CLK _9689_/D _9689_/SET_B VGND VGND VPWR VPWR _9689_/Q sky130_fd_sc_hd__dfstp_1
X_8709_ _8709_/A _8709_/B VGND VGND VPWR VPWR _8710_/B sky130_fd_sc_hd__or2_1
XFILLER_41_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5370_ _9525_/Q _5369_/A hold516/A _5369_/Y VGND VGND VPWR VPWR _5370_/X sky130_fd_sc_hd__a22o_1
XFILLER_126_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7040_ _9093_/Q _6024_/B _9092_/Q _7039_/X VGND VGND VPWR VPWR _9092_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8991_ _8990_/X hold359/X _9629_/Q VGND VGND VPWR VPWR _8991_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7942_ _8005_/A _8230_/A _7942_/C _8234_/A VGND VGND VPWR VPWR _7943_/A sky130_fd_sc_hd__or4_1
XFILLER_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7873_ _7873_/A _7873_/B _7873_/C VGND VGND VPWR VPWR _8704_/A sky130_fd_sc_hd__and3_1
X_9612_ _9731_/CLK _9612_/D _9731_/SET_B VGND VGND VPWR VPWR _9612_/Q sky130_fd_sc_hd__dfrtp_1
X_6824_ _9389_/Q VGND VGND VPWR VPWR _6824_/Y sky130_fd_sc_hd__inv_6
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9543_ _9576_/CLK _9543_/D _9537_/SET_B VGND VGND VPWR VPWR _9543_/Q sky130_fd_sc_hd__dfrtp_1
X_6755_ _9416_/Q VGND VGND VPWR VPWR _6755_/Y sky130_fd_sc_hd__inv_2
X_5706_ _5847_/A _5706_/B VGND VGND VPWR VPWR _5707_/A sky130_fd_sc_hd__or2_1
X_9474_ _9483_/CLK _9474_/D _9727_/SET_B VGND VGND VPWR VPWR _9474_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8425_ _8678_/A _8556_/A VGND VGND VPWR VPWR _8693_/B sky130_fd_sc_hd__or2_1
XFILLER_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6686_ _6681_/Y _6058_/B _6682_/Y _4623_/B _6685_/X VGND VGND VPWR VPWR _6722_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5637_ _5637_/A VGND VGND VPWR VPWR _5638_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5568_ _9389_/Q _5561_/A hold593/X _5561_/Y VGND VGND VPWR VPWR _9389_/D sky130_fd_sc_hd__a22o_1
X_8356_ _8358_/A _8306_/B _8496_/A VGND VGND VPWR VPWR _8356_/X sky130_fd_sc_hd__o21a_1
XFILLER_191_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold130 _9744_/Q VGND VGND VPWR VPWR hold131/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _5617_/X VGND VGND VPWR VPWR hold153/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 hold141/A VGND VGND VPWR VPWR hold142/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7307_ _6157_/Y _7161_/X _6114_/Y _7162_/X VGND VGND VPWR VPWR _7307_/X sky130_fd_sc_hd__o22a_1
XFILLER_132_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8287_ _8287_/A _8404_/B _8617_/B VGND VGND VPWR VPWR _8290_/A sky130_fd_sc_hd__or3_1
X_4519_ _9822_/Q _4513_/A _8965_/A1 _4513_/Y VGND VGND VPWR VPWR _9822_/D sky130_fd_sc_hd__a22o_1
Xhold174 hold174/A VGND VGND VPWR VPWR hold175/A sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _9436_/Q hold632/X _8959_/A1 _5495_/Y VGND VGND VPWR VPWR _5499_/X sky130_fd_sc_hd__a22o_1
Xhold163 hold163/A VGND VGND VPWR VPWR _9546_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold185 _5388_/X VGND VGND VPWR VPWR hold186/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7238_ _6427_/Y _7149_/X _6399_/Y _7150_/X _7237_/X VGND VGND VPWR VPWR _7243_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_78_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold196 hold196/A VGND VGND VPWR VPWR _9118_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7169_ _6926_/Y _7167_/X _6920_/Y _7168_/X VGND VGND VPWR VPWR _7169_/X sky130_fd_sc_hd__o22a_1
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4870_ _9453_/Q VGND VGND VPWR VPWR _4870_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6540_ _9365_/Q VGND VGND VPWR VPWR _8805_/A sky130_fd_sc_hd__inv_4
XFILLER_146_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6471_ _9400_/Q VGND VGND VPWR VPWR _6471_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_173_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8210_ _8210_/A VGND VGND VPWR VPWR _8415_/A sky130_fd_sc_hd__inv_2
X_5422_ _9489_/Q _5419_/A hold696/X _5419_/Y VGND VGND VPWR VPWR _9489_/D sky130_fd_sc_hd__a22o_1
X_9190_ _9297_/CLK _9190_/D _9797_/SET_B VGND VGND VPWR VPWR _9190_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput235 _8875_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_2
Xoutput224 _8824_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_2
X_8141_ _8141_/A VGND VGND VPWR VPWR _8255_/A sky130_fd_sc_hd__buf_4
Xoutput213 _8804_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_2
X_5353_ _5353_/A VGND VGND VPWR VPWR _5353_/Y sky130_fd_sc_hd__inv_2
Xoutput268 _9049_/Z VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_2
Xoutput257 _9039_/Z VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_2
Xoutput246 _9029_/Z VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_2
XFILLER_114_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8072_ _8053_/A _8592_/A _8071_/X VGND VGND VPWR VPWR _8074_/A sky130_fd_sc_hd__o21ai_1
Xoutput279 _9025_/Z VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_2
X_5284_ _5284_/A VGND VGND VPWR VPWR _5284_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7023_ _5669_/Y _5782_/B _9095_/Q _7022_/Y VGND VGND VPWR VPWR _9095_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8974_ _9645_/Q hold593/X _8975_/S VGND VGND VPWR VPWR _8974_/X sky130_fd_sc_hd__mux2_1
X_7925_ _8608_/A _7925_/B _7918_/B _7924_/X VGND VGND VPWR VPWR _7925_/X sky130_fd_sc_hd__or4bb_1
XFILLER_43_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7856_ _7856_/A VGND VGND VPWR VPWR _8702_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_63_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6807_ _6805_/Y _5144_/B _6806_/Y _5979_/B VGND VGND VPWR VPWR _6807_/X sky130_fd_sc_hd__o22a_1
X_4999_ hold46/A _4989_/A hold36/A _4989_/Y VGND VGND VPWR VPWR _9746_/D sky130_fd_sc_hd__a22o_1
X_7787_ _8421_/D _8436_/B _7875_/B VGND VGND VPWR VPWR _8702_/A sky130_fd_sc_hd__or3_4
XFILLER_23_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9526_ _9800_/CLK _9526_/D _9817_/SET_B VGND VGND VPWR VPWR _9526_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6738_ _9346_/Q VGND VGND VPWR VPWR _6738_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6669_ _9270_/Q VGND VGND VPWR VPWR _6669_/Y sky130_fd_sc_hd__inv_2
X_9457_ _9579_/CLK _9457_/D _7042_/B VGND VGND VPWR VPWR _9457_/Q sky130_fd_sc_hd__dfrtp_1
X_9388_ _9694_/CLK _9388_/D _9689_/SET_B VGND VGND VPWR VPWR _9388_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_191_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8408_ _8727_/B _8535_/B VGND VGND VPWR VPWR _8717_/A sky130_fd_sc_hd__or2_1
X_8339_ _8693_/A _8648_/B VGND VGND VPWR VPWR _8715_/A sky130_fd_sc_hd__or2_2
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5971_ _5990_/A _5971_/B VGND VGND VPWR VPWR _5972_/A sky130_fd_sc_hd__or2_1
X_8690_ _8608_/B _8256_/Y _8382_/C VGND VGND VPWR VPWR _8723_/B sky130_fd_sc_hd__o21a_1
X_4922_ _4951_/B _4922_/B VGND VGND VPWR VPWR _5428_/B sky130_fd_sc_hd__or2_4
X_7710_ _6559_/Y _7525_/A _7402_/A _7526_/A _7709_/X VGND VGND VPWR VPWR _7711_/D
+ sky130_fd_sc_hd__o221a_1
X_7641_ _4946_/Y _7487_/X _4712_/A _7488_/X VGND VGND VPWR VPWR _7641_/X sky130_fd_sc_hd__o22a_1
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4853_ _4853_/A VGND VGND VPWR VPWR _4853_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7572_ _6403_/Y _7491_/X _6493_/Y _7492_/X _7571_/X VGND VGND VPWR VPWR _7586_/B
+ sky130_fd_sc_hd__o221a_1
X_4784_ _9370_/Q VGND VGND VPWR VPWR _4784_/Y sky130_fd_sc_hd__inv_2
X_6523_ _9249_/Q VGND VGND VPWR VPWR _8793_/A sky130_fd_sc_hd__clkinv_4
X_9311_ _9574_/CLK _9311_/D _9571_/SET_B VGND VGND VPWR VPWR _9311_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_20_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_opt_2_0_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_146_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9242_ _9600_/CLK _9242_/D _9821_/SET_B VGND VGND VPWR VPWR _9242_/Q sky130_fd_sc_hd__dfstp_1
X_6454_ _9452_/Q VGND VGND VPWR VPWR _6454_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5405_ _5770_/A VGND VGND VPWR VPWR _5570_/A sky130_fd_sc_hd__buf_8
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9173_ _9225_/CLK _9173_/D _9731_/SET_B VGND VGND VPWR VPWR _9173_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6385_ _9673_/Q VGND VGND VPWR VPWR _6385_/Y sky130_fd_sc_hd__clkinv_2
X_5336_ _9547_/Q _5331_/A _8964_/A1 _5331_/Y VGND VGND VPWR VPWR _9547_/D sky130_fd_sc_hd__a22o_1
X_8124_ _8226_/A _8228_/A _8124_/C VGND VGND VPWR VPWR _8127_/A sky130_fd_sc_hd__and3_1
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8055_ _7941_/B _8053_/B _8134_/A VGND VGND VPWR VPWR _8056_/D sky130_fd_sc_hd__a21oi_1
X_5267_ _9594_/Q _5265_/A hold510/X _5265_/Y VGND VGND VPWR VPWR _9594_/D sky130_fd_sc_hd__a22o_1
X_7006_ _7006_/A VGND VGND VPWR VPWR _7007_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5198_ _9638_/Q _5192_/A hold136/X _5192_/Y VGND VGND VPWR VPWR _5198_/X sky130_fd_sc_hd__a22o_1
X_8957_ _9650_/Q hold510/X _8975_/S VGND VGND VPWR VPWR _8957_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7908_ _8268_/C _8358_/A VGND VGND VPWR VPWR _7909_/A sky130_fd_sc_hd__or2_1
XFILLER_43_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8888_ hold245/X hold515/X _8987_/S VGND VGND VPWR VPWR _8888_/X sky130_fd_sc_hd__mux2_8
XFILLER_169_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7839_ _8229_/B _8666_/B VGND VGND VPWR VPWR _8604_/A sky130_fd_sc_hd__nor2_2
XFILLER_34_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9509_ _9800_/CLK _9509_/D _9817_/SET_B VGND VGND VPWR VPWR _9509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold707 _9216_/Q VGND VGND VPWR VPWR hold707/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6170_ _9305_/Q VGND VGND VPWR VPWR _6170_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5121_ _9689_/Q _5114_/A hold593/X _5114_/Y VGND VGND VPWR VPWR _9689_/D sky130_fd_sc_hd__a22o_1
XFILLER_170_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_3_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9729_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5052_ _9727_/Q _5049_/A hold217/X _5049_/Y VGND VGND VPWR VPWR _9727_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8811_ _8811_/A VGND VGND VPWR VPWR _8812_/A sky130_fd_sc_hd__clkbuf_1
X_9791_ _9791_/CLK _9791_/D _9821_/SET_B VGND VGND VPWR VPWR _9791_/Q sky130_fd_sc_hd__dfstp_1
X_8742_ _8557_/B _8229_/A _8383_/B VGND VGND VPWR VPWR _8742_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5954_ _9107_/D VGND VGND VPWR VPWR _6178_/B sky130_fd_sc_hd__inv_2
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8673_ _8673_/A _8673_/B VGND VGND VPWR VPWR _8730_/C sky130_fd_sc_hd__or2_1
X_5885_ _5878_/X _8902_/X _8960_/X _9212_/Q VGND VGND VPWR VPWR _9212_/D sky130_fd_sc_hd__o22a_1
X_4905_ _9578_/Q VGND VGND VPWR VPWR _4905_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_52_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7624_ _6122_/Y _7485_/X _6170_/Y _7486_/X _7623_/X VGND VGND VPWR VPWR _7640_/A
+ sky130_fd_sc_hd__o221a_1
X_4836_ _9112_/Q VGND VGND VPWR VPWR _4836_/Y sky130_fd_sc_hd__inv_4
XFILLER_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7555_ _8835_/A _7498_/X _8805_/A _5727_/X VGND VGND VPWR VPWR _7555_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6506_ _6506_/A _6506_/B _6506_/C _6506_/D VGND VGND VPWR VPWR _6506_/Y sky130_fd_sc_hd__nand4_2
X_4767_ _4763_/Y _5598_/B _4765_/Y _6112_/B VGND VGND VPWR VPWR _4767_/X sky130_fd_sc_hd__o22a_1
X_7486_ _7486_/A VGND VGND VPWR VPWR _7486_/X sky130_fd_sc_hd__buf_6
X_4698_ _4808_/B _4865_/B VGND VGND VPWR VPWR _5103_/B sky130_fd_sc_hd__or2_4
XFILLER_161_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9225_ _9225_/CLK _9225_/D _9537_/SET_B VGND VGND VPWR VPWR _9225_/Q sky130_fd_sc_hd__dfrtp_1
X_6437_ _6435_/Y _5505_/B _6436_/Y _4598_/B VGND VGND VPWR VPWR _6437_/X sky130_fd_sc_hd__o22a_1
XFILLER_161_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6368_ _9171_/Q VGND VGND VPWR VPWR _6368_/Y sky130_fd_sc_hd__clkinv_2
X_9156_ _9678_/CLK _9156_/D _9730_/SET_B VGND VGND VPWR VPWR _9156_/Q sky130_fd_sc_hd__dfrtp_1
X_8107_ _8324_/B _8560_/A _8324_/C VGND VGND VPWR VPWR _8581_/A sky130_fd_sc_hd__and3_2
XFILLER_121_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5319_ _9558_/Q _5315_/A _6067_/B1 _5315_/Y VGND VGND VPWR VPWR _9558_/D sky130_fd_sc_hd__a22o_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9087_ _9832_/CLK _9087_/D VGND VGND VPWR VPWR _9087_/Q sky130_fd_sc_hd__dfxtp_1
X_6299_ _9809_/Q VGND VGND VPWR VPWR _6299_/Y sky130_fd_sc_hd__inv_2
Xhold23 hold23/A VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_8038_ _8038_/A VGND VGND VPWR VPWR _8443_/A sky130_fd_sc_hd__clkbuf_4
Xhold34 hold34/A VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold67 hold67/A VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 _4792_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _9097_/Q VGND VGND VPWR VPWR _5752_/B sky130_fd_sc_hd__inv_2
X_4621_ _9774_/Q _4613_/A _6008_/B1 _4613_/Y VGND VGND VPWR VPWR _9774_/D sky130_fd_sc_hd__a22o_1
XFILLER_156_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7340_ _7340_/A _7340_/B _7340_/C _7340_/D VGND VGND VPWR VPWR _7341_/C sky130_fd_sc_hd__and4_1
X_4552_ _9807_/Q _4547_/A _6065_/B1 _4547_/Y VGND VGND VPWR VPWR _9807_/D sky130_fd_sc_hd__a22o_1
Xhold515 hold515/A VGND VGND VPWR VPWR hold515/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold526 _5573_/X VGND VGND VPWR VPWR _9387_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7271_ _6277_/Y _5756_/X _6334_/Y _7071_/A _7270_/X VGND VGND VPWR VPWR _7274_/C
+ sky130_fd_sc_hd__o221a_1
X_4483_ _5201_/A _6282_/A VGND VGND VPWR VPWR _4484_/A sky130_fd_sc_hd__or2_1
Xhold504 hold504/A VGND VGND VPWR VPWR hold504/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_9010_ _7783_/X _9010_/A1 _9017_/S VGND VGND VPWR VPWR _9010_/X sky130_fd_sc_hd__mux2_1
Xhold537 _5182_/X VGND VGND VPWR VPWR _9651_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold548 _5790_/X VGND VGND VPWR VPWR _9279_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold559 _5459_/X VGND VGND VPWR VPWR _9464_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6222_ input41/X _8971_/S _6221_/Y _5455_/B VGND VGND VPWR VPWR _6222_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_143_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6153_ _9280_/Q VGND VGND VPWR VPWR _6153_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6084_ _6084_/A VGND VGND VPWR VPWR _6085_/A sky130_fd_sc_hd__clkbuf_2
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5104_ _5104_/A VGND VGND VPWR VPWR _5105_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _9090_/Q _8999_/S _4971_/A _9738_/Q _5034_/X VGND VGND VPWR VPWR _9738_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_72_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater398 hold593/A VGND VGND VPWR VPWR _8969_/A1 sky130_fd_sc_hd__buf_12
X_6986_ _6357_/Y _6983_/A _9075_/Q _6983_/Y VGND VGND VPWR VPWR _9075_/D sky130_fd_sc_hd__o22a_1
X_9774_ _9819_/CLK _9774_/D _9821_/SET_B VGND VGND VPWR VPWR _9774_/Q sky130_fd_sc_hd__dfstp_1
X_5937_ _5937_/A VGND VGND VPWR VPWR _5937_/Y sky130_fd_sc_hd__inv_2
X_8725_ _8725_/A _8725_/B VGND VGND VPWR VPWR _8725_/X sky130_fd_sc_hd__or2_1
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8656_ _8656_/A _8656_/B _8656_/C _8656_/D VGND VGND VPWR VPWR _8710_/D sky130_fd_sc_hd__or4_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5868_ _5868_/A VGND VGND VPWR VPWR _5868_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7607_ _6263_/Y _7493_/X _6220_/Y _7494_/X VGND VGND VPWR VPWR _7607_/X sky130_fd_sc_hd__o22a_1
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8587_ _8667_/B VGND VGND VPWR VPWR _8596_/B sky130_fd_sc_hd__clkinv_4
X_4819_ _9763_/Q VGND VGND VPWR VPWR _4819_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5799_ _5799_/A VGND VGND VPWR VPWR _5799_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7538_ _6725_/Y _7502_/X _6791_/Y _7503_/X VGND VGND VPWR VPWR _7538_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7469_ _4761_/Y _7513_/A _4938_/Y _7514_/A _7468_/X VGND VGND VPWR VPWR _7482_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9208_ _9212_/CLK _9208_/D _9797_/SET_B VGND VGND VPWR VPWR _9208_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9139_ _9574_/CLK _9139_/D _9571_/SET_B VGND VGND VPWR VPWR _9139_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput102 sram_ro_data[18] VGND VGND VPWR VPWR _6775_/A sky130_fd_sc_hd__clkbuf_1
Xinput135 wb_adr_i[12] VGND VGND VPWR VPWR _7806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput113 sram_ro_data[28] VGND VGND VPWR VPWR _6475_/A sky130_fd_sc_hd__clkbuf_1
Xinput124 sram_ro_data[9] VGND VGND VPWR VPWR _6839_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput168 wb_dat_i[12] VGND VGND VPWR VPWR _7777_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput146 wb_adr_i[22] VGND VGND VPWR VPWR _7816_/B sky130_fd_sc_hd__clkbuf_1
Xinput157 wb_adr_i[3] VGND VGND VPWR VPWR _8421_/D sky130_fd_sc_hd__buf_4
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput179 wb_dat_i[22] VGND VGND VPWR VPWR _7780_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6840_ _6838_/Y _4502_/B _6839_/Y _4915_/X VGND VGND VPWR VPWR _6840_/X sky130_fd_sc_hd__o22a_1
X_6771_ _6766_/Y _5301_/B _6767_/Y _5367_/B _6770_/X VGND VGND VPWR VPWR _6772_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_90_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8510_ _8510_/A _8672_/A VGND VGND VPWR VPWR _8512_/B sky130_fd_sc_hd__or2_1
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5722_ _9296_/Q _9295_/Q VGND VGND VPWR VPWR _7467_/A sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_21_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9643_/CLK sky130_fd_sc_hd__clkbuf_16
X_9490_ _9491_/CLK _9490_/D _9731_/SET_B VGND VGND VPWR VPWR _9490_/Q sky130_fd_sc_hd__dfrtp_1
X_5653_ _9332_/Q _5649_/A hold53/X _5649_/Y VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__a22o_1
X_8441_ _8243_/B _8158_/B _8437_/X _8440_/Y VGND VGND VPWR VPWR _8441_/X sky130_fd_sc_hd__o211a_1
X_8372_ _8418_/A _8372_/B VGND VGND VPWR VPWR _8373_/B sky130_fd_sc_hd__or2_1
XFILLER_148_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4604_ _9786_/Q _4600_/A _6064_/B1 _4600_/Y VGND VGND VPWR VPWR _9786_/D sky130_fd_sc_hd__a22o_1
X_5584_ _9379_/Q _5583_/A _6064_/B1 _5583_/Y VGND VGND VPWR VPWR _9379_/D sky130_fd_sc_hd__a22o_1
Xhold301 hold301/A VGND VGND VPWR VPWR hold302/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4535_ _8981_/X _4823_/B _4685_/C VGND VGND VPWR VPWR _6117_/A sky130_fd_sc_hd__or3_4
X_7323_ _4697_/Y _7071_/C _4796_/Y _7146_/X VGND VGND VPWR VPWR _7323_/X sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_36_csclk clkbuf_opt_2_0_csclk/X VGND VGND VPWR VPWR _9832_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold323 hold323/A VGND VGND VPWR VPWR _9411_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold334 hold334/A VGND VGND VPWR VPWR hold335/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _5345_/X VGND VGND VPWR VPWR hold313/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold378 hold378/A VGND VGND VPWR VPWR hold379/A sky130_fd_sc_hd__dlygate4sd3_1
X_7254_ _6305_/Y _7139_/X _6270_/Y _7140_/X VGND VGND VPWR VPWR _7254_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4466_ _9614_/Q _4971_/A _9724_/Q VGND VGND VPWR VPWR _9029_/A sky130_fd_sc_hd__mux2_1
Xhold367 hold367/A VGND VGND VPWR VPWR hold368/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 hold625/X VGND VGND VPWR VPWR _4534_/D sky130_fd_sc_hd__buf_2
Xhold345 _4538_/X VGND VGND VPWR VPWR hold346/A sky130_fd_sc_hd__dlygate4sd3_1
X_6205_ _6205_/A _6205_/B _6205_/C _6205_/D VGND VGND VPWR VPWR _6268_/A sky130_fd_sc_hd__and4_1
X_7185_ _6902_/Y _7180_/X _6915_/Y _7181_/X _7184_/X VGND VGND VPWR VPWR _7186_/D
+ sky130_fd_sc_hd__o221a_1
Xhold389 _5552_/X VGND VGND VPWR VPWR hold390/A sky130_fd_sc_hd__dlygate4sd3_1
X_6136_ _9681_/Q VGND VGND VPWR VPWR _6136_/Y sky130_fd_sc_hd__inv_2
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _9113_/Q _6060_/A _6067_/B1 _6060_/Y VGND VGND VPWR VPWR _6067_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5018_ _5018_/A VGND VGND VPWR VPWR _5018_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9826_ _9827_/CLK _9826_/D _9797_/SET_B VGND VGND VPWR VPWR _9826_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6969_ _9350_/Q VGND VGND VPWR VPWR _6969_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9757_ _8879_/A1 _9757_/D _4666_/X VGND VGND VPWR VPWR _9757_/Q sky130_fd_sc_hd__dfrtn_1
X_9688_ _9695_/CLK _9688_/D _9689_/SET_B VGND VGND VPWR VPWR _9688_/Q sky130_fd_sc_hd__dfstp_1
X_8708_ _8708_/A _8708_/B _8708_/C _8708_/D VGND VGND VPWR VPWR _8777_/D sky130_fd_sc_hd__or4_2
XFILLER_139_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8639_ _8639_/A _8639_/B _8639_/C _8639_/D VGND VGND VPWR VPWR _8699_/D sky130_fd_sc_hd__or4_4
XFILLER_166_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8990_ _9129_/Q _9128_/Q _9093_/Q VGND VGND VPWR VPWR _8990_/X sky130_fd_sc_hd__mux2_1
X_7941_ _8042_/B _7941_/B VGND VGND VPWR VPWR _7941_/X sky130_fd_sc_hd__or2_1
XFILLER_82_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7872_ _8489_/A VGND VGND VPWR VPWR _7873_/B sky130_fd_sc_hd__inv_4
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9611_ _9751_/CLK _9611_/D _5236_/X VGND VGND VPWR VPWR _9611_/Q sky130_fd_sc_hd__dfrtp_4
X_6823_ _6818_/Y _5378_/B _6819_/Y _4869_/X _6822_/X VGND VGND VPWR VPWR _6861_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_149_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9542_ _9576_/CLK _9542_/D _9537_/SET_B VGND VGND VPWR VPWR _9542_/Q sky130_fd_sc_hd__dfrtp_1
X_6754_ _9481_/Q VGND VGND VPWR VPWR _6754_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_148_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9473_ _9577_/CLK _9473_/D _9571_/SET_B VGND VGND VPWR VPWR _9473_/Q sky130_fd_sc_hd__dfrtp_1
X_6685_ _6683_/Y _4525_/B _6684_/Y _5201_/B VGND VGND VPWR VPWR _6685_/X sky130_fd_sc_hd__o22a_1
X_5705_ _9306_/Q _5700_/A _6008_/B1 _5700_/Y VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8424_ _8747_/A _8424_/B VGND VGND VPWR VPWR _8426_/A sky130_fd_sc_hd__or2_1
X_5636_ _5847_/A _5636_/B VGND VGND VPWR VPWR _5637_/A sky130_fd_sc_hd__or2_1
XFILLER_148_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5567_ _9390_/Q _5561_/A hold136/X _5561_/Y VGND VGND VPWR VPWR _5567_/X sky130_fd_sc_hd__a22o_1
X_8355_ _8538_/A _8348_/X _8272_/A _8540_/B _8354_/X VGND VGND VPWR VPWR _8355_/X
+ sky130_fd_sc_hd__o221a_2
Xhold131 hold131/A VGND VGND VPWR VPWR hold132/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 hold120/A VGND VGND VPWR VPWR hold120/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold153 hold153/A VGND VGND VPWR VPWR hold154/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 hold142/A VGND VGND VPWR VPWR _9520_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_5498_ _9437_/Q _5495_/A hold577/A _5495_/Y VGND VGND VPWR VPWR _5498_/X sky130_fd_sc_hd__a22o_1
X_7306_ _6098_/Y _7155_/X _6112_/A _7156_/X _7305_/X VGND VGND VPWR VPWR _7309_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8286_ _8358_/A _8302_/B VGND VGND VPWR VPWR _8617_/B sky130_fd_sc_hd__nor2_1
X_4518_ _9823_/Q hold648/X _8964_/A1 _4513_/Y VGND VGND VPWR VPWR _9823_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold175 hold175/A VGND VGND VPWR VPWR hold176/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _5463_/X VGND VGND VPWR VPWR hold165/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold186 hold186/A VGND VGND VPWR VPWR hold187/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7237_ _6360_/Y _7151_/X _6380_/Y _7152_/X VGND VGND VPWR VPWR _7237_/X sky130_fd_sc_hd__o22a_1
Xhold197 _8970_/X VGND VGND VPWR VPWR hold198/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7168_ _7168_/A VGND VGND VPWR VPWR _7168_/X sky130_fd_sc_hd__buf_4
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _6116_/Y _6117_/X _6118_/Y _4892_/X VGND VGND VPWR VPWR _6119_/X sky130_fd_sc_hd__o22a_1
X_7099_ _7127_/A _7099_/B VGND VGND VPWR VPWR _7139_/A sky130_fd_sc_hd__or2_2
XFILLER_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9809_ _9817_/CLK _9809_/D _9817_/SET_B VGND VGND VPWR VPWR _9809_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_186_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6470_ _9692_/Q VGND VGND VPWR VPWR _6470_/Y sky130_fd_sc_hd__inv_4
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5421_ _9490_/Q _5419_/A hold510/X _5419_/Y VGND VGND VPWR VPWR _9490_/D sky130_fd_sc_hd__a22o_1
Xoutput225 _8826_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_2
X_8140_ _8140_/A _8140_/B VGND VGND VPWR VPWR _8141_/A sky130_fd_sc_hd__or2_1
Xoutput214 _8806_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_2
Xoutput203 _8848_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_2
X_5352_ _5352_/A VGND VGND VPWR VPWR _5353_/A sky130_fd_sc_hd__clkbuf_2
Xoutput236 _8876_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_2
Xoutput258 _9040_/Z VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_2
XFILLER_126_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput247 _9030_/Z VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_99_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8071_ _8429_/A _8592_/A _8067_/X _8452_/A _8070_/X VGND VGND VPWR VPWR _8071_/X
+ sky130_fd_sc_hd__o2111a_1
Xoutput269 _9050_/Z VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_141_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7022_ _9833_/Q VGND VGND VPWR VPWR _7022_/Y sky130_fd_sc_hd__inv_2
X_5283_ _5283_/A VGND VGND VPWR VPWR _5284_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8973_ _9666_/Q hold510/X _8973_/S VGND VGND VPWR VPWR _8973_/X sky130_fd_sc_hd__mux2_1
X_7924_ _7957_/A _7924_/B VGND VGND VPWR VPWR _7924_/X sky130_fd_sc_hd__or2_1
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7855_ _7942_/C _8570_/A _8625_/A _7933_/B VGND VGND VPWR VPWR _7856_/A sky130_fd_sc_hd__or4_1
X_6806_ _9150_/Q VGND VGND VPWR VPWR _6806_/Y sky130_fd_sc_hd__inv_2
X_4998_ _4998_/A VGND VGND VPWR VPWR _4998_/X sky130_fd_sc_hd__clkbuf_1
X_9525_ _9569_/CLK _9525_/D _9563_/SET_B VGND VGND VPWR VPWR _9525_/Q sky130_fd_sc_hd__dfrtp_1
X_7786_ _8436_/C _7876_/A VGND VGND VPWR VPWR _7875_/B sky130_fd_sc_hd__or2_2
XFILLER_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6737_ _6737_/A VGND VGND VPWR VPWR _6737_/Y sky130_fd_sc_hd__clkinv_2
X_6668_ _9248_/Q VGND VGND VPWR VPWR _6668_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_149_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9456_ _9579_/CLK _9456_/D _9727_/SET_B VGND VGND VPWR VPWR _9456_/Q sky130_fd_sc_hd__dfrtp_1
X_5619_ _9354_/Q _5611_/A hold601/A _5611_/Y VGND VGND VPWR VPWR _5619_/X sky130_fd_sc_hd__a22o_1
X_9387_ _9522_/CLK _9387_/D _9563_/SET_B VGND VGND VPWR VPWR _9387_/Q sky130_fd_sc_hd__dfrtp_1
X_6599_ _9539_/Q VGND VGND VPWR VPWR _8831_/A sky130_fd_sc_hd__clkinv_8
X_8407_ _8593_/A _8420_/B _8292_/A VGND VGND VPWR VPWR _8619_/C sky130_fd_sc_hd__o21ai_1
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8338_ _8338_/A _8338_/B VGND VGND VPWR VPWR _8338_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8269_ _8637_/B _8269_/B _8613_/B _8541_/B VGND VGND VPWR VPWR _8273_/A sky130_fd_sc_hd__or4_1
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5970_ _9101_/Q _7763_/A _9161_/Q _5968_/Y _5969_/X VGND VGND VPWR VPWR _9161_/D
+ sky130_fd_sc_hd__o221a_1
X_4921_ _9479_/Q VGND VGND VPWR VPWR _4921_/Y sky130_fd_sc_hd__clkinv_2
X_7640_ _7640_/A _7640_/B _7640_/C _7640_/D VGND VGND VPWR VPWR _7640_/Y sky130_fd_sc_hd__nand4_4
X_4852_ _4852_/A _4852_/B _4852_/C _4852_/D VGND VGND VPWR VPWR _4957_/A sky130_fd_sc_hd__and4_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7571_ _6494_/Y _7493_/X _6434_/Y _7494_/X VGND VGND VPWR VPWR _7571_/X sky130_fd_sc_hd__o22a_1
X_4783_ _4913_/A _4865_/B VGND VGND VPWR VPWR _5858_/B sky130_fd_sc_hd__or2_4
XFILLER_186_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6522_ _9383_/Q VGND VGND VPWR VPWR _6522_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_158_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9310_ _9831_/CLK _9310_/D _9727_/SET_B VGND VGND VPWR VPWR _9310_/Q sky130_fd_sc_hd__dfrtp_1
X_6453_ _9488_/Q VGND VGND VPWR VPWR _6453_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9241_ _9600_/CLK _9241_/D _9821_/SET_B VGND VGND VPWR VPWR _9241_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9172_ _9225_/CLK _9172_/D _9731_/SET_B VGND VGND VPWR VPWR _9172_/Q sky130_fd_sc_hd__dfrtp_1
X_5404_ _9500_/Q _5399_/A _6008_/B1 _5399_/Y VGND VGND VPWR VPWR _9500_/D sky130_fd_sc_hd__a22o_1
X_6384_ _9236_/Q VGND VGND VPWR VPWR _6384_/Y sky130_fd_sc_hd__clkinv_4
X_8123_ _8123_/A _8227_/A VGND VGND VPWR VPWR _8124_/C sky130_fd_sc_hd__and2_1
X_5335_ _9548_/Q _5331_/A _8959_/A1 _5331_/Y VGND VGND VPWR VPWR _9548_/D sky130_fd_sc_hd__a22o_1
X_8054_ _8068_/A _8158_/A _8053_/X VGND VGND VPWR VPWR _8056_/C sky130_fd_sc_hd__o21ai_1
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5266_ _9595_/Q _5265_/A hold516/X _5265_/Y VGND VGND VPWR VPWR _9595_/D sky130_fd_sc_hd__a22o_1
X_7005_ _7005_/A _7005_/B VGND VGND VPWR VPWR _7006_/A sky130_fd_sc_hd__or2_1
XFILLER_102_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5197_ _9639_/Q _5192_/A hold612/X _5192_/Y VGND VGND VPWR VPWR _9639_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8956_ _9649_/Q hold577/A _8975_/S VGND VGND VPWR VPWR _8956_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7907_ _7907_/A VGND VGND VPWR VPWR _8358_/A sky130_fd_sc_hd__buf_2
X_8887_ hold191/X hold509/X _8987_/S VGND VGND VPWR VPWR _8887_/X sky130_fd_sc_hd__mux2_8
X_7838_ _8065_/A VGND VGND VPWR VPWR _8666_/B sky130_fd_sc_hd__buf_6
XFILLER_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7769_ _9110_/Q _7769_/A2 _9109_/Q _7769_/B2 _7768_/X VGND VGND VPWR VPWR _7769_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_184_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9508_ _9800_/CLK _9508_/D _9817_/SET_B VGND VGND VPWR VPWR _9508_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9439_ _9522_/CLK _9439_/D _9563_/SET_B VGND VGND VPWR VPWR _9439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold708 _9753_/Q VGND VGND VPWR VPWR hold708/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5120_ _9690_/Q _5114_/A hold136/X _5114_/Y VGND VGND VPWR VPWR _5120_/X sky130_fd_sc_hd__a22o_1
XFILLER_151_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5051_ _9728_/Q _5049_/A _6065_/B1 _5049_/Y VGND VGND VPWR VPWR _9728_/D sky130_fd_sc_hd__a22o_1
XFILLER_111_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8810_ _8810_/A VGND VGND VPWR VPWR _8810_/X sky130_fd_sc_hd__clkbuf_1
X_9790_ _9791_/CLK _9790_/D _9821_/SET_B VGND VGND VPWR VPWR _9790_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_37_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8741_ _8741_/A _8741_/B _8741_/C _8741_/D VGND VGND VPWR VPWR _8774_/A sky130_fd_sc_hd__or4_1
XFILLER_92_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5953_ _9162_/Q _5948_/A _8975_/A1 _5948_/Y VGND VGND VPWR VPWR _9162_/D sky130_fd_sc_hd__a22o_1
X_8672_ _8672_/A _8672_/B _8672_/C _8672_/D VGND VGND VPWR VPWR _8751_/C sky130_fd_sc_hd__or4_2
XFILLER_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4904_ _9815_/Q VGND VGND VPWR VPWR _4904_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_33_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5884_ _5878_/X _8904_/X _8960_/X _9213_/Q VGND VGND VPWR VPWR _9213_/D sky130_fd_sc_hd__o22a_1
X_7623_ _6109_/Y _7487_/X _6090_/Y _7488_/X VGND VGND VPWR VPWR _7623_/X sky130_fd_sc_hd__o22a_1
X_4835_ _9803_/Q VGND VGND VPWR VPWR _4835_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_21_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7554_ _8795_/A _7491_/X _8787_/A _7492_/X _7553_/X VGND VGND VPWR VPWR _7568_/B
+ sky130_fd_sc_hd__o221a_1
X_4766_ _4803_/A _4827_/A VGND VGND VPWR VPWR _6112_/B sky130_fd_sc_hd__or2_4
X_6505_ _6505_/A _6505_/B _6505_/C _6505_/D VGND VGND VPWR VPWR _6506_/D sky130_fd_sc_hd__and4_1
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7485_ _7485_/A VGND VGND VPWR VPWR _7485_/X sky130_fd_sc_hd__buf_6
X_4697_ _9696_/Q VGND VGND VPWR VPWR _4697_/Y sky130_fd_sc_hd__clkinv_2
X_9224_ _9420_/CLK _9224_/D _9537_/SET_B VGND VGND VPWR VPWR _9224_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6436_ _9786_/Q VGND VGND VPWR VPWR _6436_/Y sky130_fd_sc_hd__inv_2
X_9155_ _9225_/CLK _9155_/D _9731_/SET_B VGND VGND VPWR VPWR _9155_/Q sky130_fd_sc_hd__dfrtp_1
X_6367_ _6367_/A VGND VGND VPWR VPWR _6367_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_130_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8106_ _8106_/A _8745_/C VGND VGND VPWR VPWR _8108_/A sky130_fd_sc_hd__or2_1
XFILLER_88_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5318_ _9559_/Q _5315_/A hold217/X _5315_/Y VGND VGND VPWR VPWR _9559_/D sky130_fd_sc_hd__a22o_1
Xhold13 hold13/A VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9086_ _9832_/CLK _9086_/D VGND VGND VPWR VPWR _9086_/Q sky130_fd_sc_hd__dfxtp_1
X_6298_ _6293_/Y _4929_/X _6294_/Y _5263_/B _6297_/X VGND VGND VPWR VPWR _6311_/B
+ sky130_fd_sc_hd__o221a_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ _9603_/Q _5241_/Y hold650/X _5241_/A VGND VGND VPWR VPWR _5249_/X sky130_fd_sc_hd__o22a_1
XFILLER_152_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8037_ _8157_/B _8037_/B VGND VGND VPWR VPWR _8038_/A sky130_fd_sc_hd__or2_1
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold24 hold24/A VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold79 hold79/A VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8939_ _9656_/Q _8959_/A1 _8971_/S VGND VGND VPWR VPWR _8939_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _9775_/Q _4613_/A _6067_/B1 _4613_/Y VGND VGND VPWR VPWR _9775_/D sky130_fd_sc_hd__a22o_1
X_4551_ _9808_/Q _4547_/A _6064_/B1 _4547_/Y VGND VGND VPWR VPWR _9808_/D sky130_fd_sc_hd__a22o_1
Xhold516 hold516/A VGND VGND VPWR VPWR hold516/X sky130_fd_sc_hd__buf_12
Xhold527 _5497_/X VGND VGND VPWR VPWR _9438_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7270_ _7270_/A _7380_/B VGND VGND VPWR VPWR _7270_/X sky130_fd_sc_hd__or2_1
Xhold505 hold690/X VGND VGND VPWR VPWR hold506/A sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ _4482_/A _4941_/A VGND VGND VPWR VPWR _6282_/A sky130_fd_sc_hd__or2_4
Xhold549 _5709_/X VGND VGND VPWR VPWR _9305_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6221_ _9464_/Q VGND VGND VPWR VPWR _6221_/Y sky130_fd_sc_hd__inv_2
Xhold538 _5381_/X VGND VGND VPWR VPWR _9517_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6152_ _9253_/Q VGND VGND VPWR VPWR _6152_/Y sky130_fd_sc_hd__clkinv_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5282_/A _5103_/B VGND VGND VPWR VPWR _5104_/A sky130_fd_sc_hd__or2_1
XFILLER_111_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6083_/A _6083_/B _6083_/C VGND VGND VPWR VPWR _6084_/A sky130_fd_sc_hd__or3_2
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5034_ _6053_/B _7034_/C VGND VGND VPWR VPWR _5034_/X sky130_fd_sc_hd__or2_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater399 hold593/X VGND VGND VPWR VPWR _6067_/B1 sky130_fd_sc_hd__buf_12
X_6985_ _6268_/Y _6983_/A _9076_/Q _6983_/Y VGND VGND VPWR VPWR _9076_/D sky130_fd_sc_hd__o22a_1
XFILLER_80_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9773_ _9817_/CLK _9773_/D _9821_/SET_B VGND VGND VPWR VPWR _9773_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8724_ _8762_/B _8764_/A _8764_/B _8765_/A VGND VGND VPWR VPWR _8724_/X sky130_fd_sc_hd__or4_2
X_5936_ _5936_/A VGND VGND VPWR VPWR _5937_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8655_ _8708_/C _8655_/B _8708_/D VGND VGND VPWR VPWR _8658_/B sky130_fd_sc_hd__or3_1
XFILLER_80_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5867_ _5867_/A VGND VGND VPWR VPWR _5868_/A sky130_fd_sc_hd__clkbuf_4
X_7606_ _6183_/Y _7485_/X _6209_/Y _7486_/X _7605_/X VGND VGND VPWR VPWR _7622_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_166_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8586_ _8586_/A _8586_/B _8586_/C VGND VGND VPWR VPWR _8667_/B sky130_fd_sc_hd__or3_2
X_4818_ _4883_/A _4818_/B VGND VGND VPWR VPWR _5144_/B sky130_fd_sc_hd__or2_4
X_5798_ _5798_/A VGND VGND VPWR VPWR _5799_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7537_ _6794_/Y _7498_/X _6692_/Y _5727_/X VGND VGND VPWR VPWR _7537_/X sky130_fd_sc_hd__o22a_1
X_4749_ _9282_/Q VGND VGND VPWR VPWR _4752_/A sky130_fd_sc_hd__inv_2
XFILLER_147_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7468_ _4826_/Y _7515_/A _4790_/Y _7516_/A VGND VGND VPWR VPWR _7468_/X sky130_fd_sc_hd__o22a_1
XFILLER_134_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9207_ _9212_/CLK _9207_/D _9797_/SET_B VGND VGND VPWR VPWR _9207_/Q sky130_fd_sc_hd__dfrtp_1
X_6419_ _6417_/Y _6117_/X _6418_/Y _5359_/B VGND VGND VPWR VPWR _6419_/X sky130_fd_sc_hd__o22a_1
XFILLER_163_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7399_ _6517_/Y _7070_/A _6539_/Y _7166_/A _7398_/X VGND VGND VPWR VPWR _7406_/A
+ sky130_fd_sc_hd__o221a_1
X_9138_ _9514_/CLK _9138_/D _9571_/SET_B VGND VGND VPWR VPWR _9138_/Q sky130_fd_sc_hd__dfrtp_2
Xinput136 wb_adr_i[13] VGND VGND VPWR VPWR _7806_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9069_ _9723_/CLK _9069_/D VGND VGND VPWR VPWR _9069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput125 trap VGND VGND VPWR VPWR _4923_/A sky130_fd_sc_hd__buf_6
XFILLER_76_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput114 sram_ro_data[29] VGND VGND VPWR VPWR _6280_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput103 sram_ro_data[19] VGND VGND VPWR VPWR _6589_/A sky130_fd_sc_hd__clkbuf_1
Xinput169 wb_dat_i[13] VGND VGND VPWR VPWR _7779_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput147 wb_adr_i[23] VGND VGND VPWR VPWR _7816_/A sky130_fd_sc_hd__clkbuf_1
Xinput158 wb_adr_i[4] VGND VGND VPWR VPWR _7933_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9831_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6770_ _6768_/Y _5559_/B _6769_/Y _5609_/B VGND VGND VPWR VPWR _6770_/X sky130_fd_sc_hd__o22a_1
XFILLER_90_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5721_ _7460_/A VGND VGND VPWR VPWR _7471_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5652_ _9333_/Q _5649_/A hold577/A _5649_/Y VGND VGND VPWR VPWR _5652_/X sky130_fd_sc_hd__a22o_1
X_8440_ _8438_/Y _8439_/Y _8162_/Y VGND VGND VPWR VPWR _8440_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8371_ _8704_/A _8642_/A _8371_/C VGND VGND VPWR VPWR _8373_/A sky130_fd_sc_hd__or3_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4603_ _9787_/Q _4600_/A hold696/A _4600_/Y VGND VGND VPWR VPWR _4603_/X sky130_fd_sc_hd__a22o_1
X_5583_ _5583_/A VGND VGND VPWR VPWR _5583_/Y sky130_fd_sc_hd__inv_2
Xhold302 hold302/A VGND VGND VPWR VPWR _9523_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4534_ _4689_/A _4642_/B _4750_/A _4534_/D VGND VGND VPWR VPWR _4890_/B sky130_fd_sc_hd__or4_4
X_7322_ _4910_/Y _7135_/X _4887_/Y _7136_/X _7321_/X VGND VGND VPWR VPWR _7341_/A
+ sky130_fd_sc_hd__o221a_1
Xhold324 _5831_/X VGND VGND VPWR VPWR hold325/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 hold335/A VGND VGND VPWR VPWR _9419_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold313 hold313/A VGND VGND VPWR VPWR hold314/A sky130_fd_sc_hd__dlygate4sd3_1
X_4465_ _9631_/Q input78/X _8875_/S VGND VGND VPWR VPWR _9052_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold368 hold368/A VGND VGND VPWR VPWR hold368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _9722_/Q VGND VGND VPWR VPWR hold358/A sky130_fd_sc_hd__dlygate4sd3_1
X_7253_ _7253_/A _7253_/B _7253_/C VGND VGND VPWR VPWR _7253_/Y sky130_fd_sc_hd__nand3_2
Xhold346 hold346/A VGND VGND VPWR VPWR hold347/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 hold379/A VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_6204_ _6199_/Y _5301_/B _6200_/Y _5329_/B _6203_/X VGND VGND VPWR VPWR _6205_/D
+ sky130_fd_sc_hd__o221a_1
X_7184_ _6854_/Y _7182_/X _6875_/Y _7183_/X VGND VGND VPWR VPWR _7184_/X sky130_fd_sc_hd__o22a_1
X_6135_ _9119_/Q VGND VGND VPWR VPWR _6135_/Y sky130_fd_sc_hd__clkinv_2
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6066_ _9114_/Q _6060_/A hold217/X _6060_/Y VGND VGND VPWR VPWR _6066_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _5017_/A VGND VGND VPWR VPWR _5018_/A sky130_fd_sc_hd__clkbuf_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9825_ _9832_/CLK _9825_/D _9821_/SET_B VGND VGND VPWR VPWR _9825_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9756_ _9751_/CLK _9756_/D _4669_/X VGND VGND VPWR VPWR _9756_/Q sky130_fd_sc_hd__dfrtn_1
X_8707_ _8707_/A _8707_/B _7916_/X VGND VGND VPWR VPWR _8708_/B sky130_fd_sc_hd__or3b_1
X_6968_ _6963_/Y _5818_/B _6964_/Y _5847_/B _6967_/X VGND VGND VPWR VPWR _6975_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_13_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5919_ _5889_/X _8926_/X _8960_/X _9186_/Q VGND VGND VPWR VPWR _9186_/D sky130_fd_sc_hd__o22a_1
X_6899_ _9584_/Q VGND VGND VPWR VPWR _6899_/Y sky130_fd_sc_hd__clkinv_4
X_9687_ _9791_/CLK _9687_/D _9817_/SET_B VGND VGND VPWR VPWR _9687_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_42_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8638_ _8118_/A _8281_/B _8278_/A _8346_/Y _8546_/B VGND VGND VPWR VPWR _8769_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_154_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8569_ _8654_/B _8569_/B _8569_/C _8708_/A VGND VGND VPWR VPWR _8573_/B sky130_fd_sc_hd__or4_1
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7940_ _8514_/A _8559_/A VGND VGND VPWR VPWR _7941_/B sky130_fd_sc_hd__or2_1
XFILLER_55_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7871_ _8268_/C VGND VGND VPWR VPWR _8489_/A sky130_fd_sc_hd__buf_4
X_9610_ _9651_/CLK _9610_/D _9563_/SET_B VGND VGND VPWR VPWR _9610_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6822_ _6820_/Y _4623_/B _6821_/Y _4545_/B VGND VGND VPWR VPWR _6822_/X sky130_fd_sc_hd__o22a_4
XFILLER_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9541_ _9576_/CLK _9541_/D _9571_/SET_B VGND VGND VPWR VPWR _9541_/Q sky130_fd_sc_hd__dfrtp_1
X_6753_ _6748_/Y _5340_/B _6749_/Y _5543_/B _6752_/X VGND VGND VPWR VPWR _6772_/A
+ sky130_fd_sc_hd__o221a_1
X_9472_ _9577_/CLK _9472_/D _9571_/SET_B VGND VGND VPWR VPWR _9472_/Q sky130_fd_sc_hd__dfrtp_1
X_6684_ _8845_/A VGND VGND VPWR VPWR _6684_/Y sky130_fd_sc_hd__inv_2
X_5704_ _9307_/Q _5700_/A _6067_/B1 _5700_/Y VGND VGND VPWR VPWR _9307_/D sky130_fd_sc_hd__a22o_1
XFILLER_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8423_ _8764_/A _8423_/B VGND VGND VPWR VPWR _8424_/B sky130_fd_sc_hd__or2_1
X_5635_ _9344_/Q _5630_/A _6008_/B1 _5630_/Y VGND VGND VPWR VPWR _9344_/D sky130_fd_sc_hd__a22o_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5566_ _9391_/Q _5561_/A hold42/X _5561_/Y VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__a22o_1
Xhold110 hold110/A VGND VGND VPWR VPWR _9648_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_151_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8354_ _8352_/X _8718_/B _8634_/A _8354_/D VGND VGND VPWR VPWR _8354_/X sky130_fd_sc_hd__and4bb_1
XFILLER_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold143 _5540_/X VGND VGND VPWR VPWR hold144/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 hold132/A VGND VGND VPWR VPWR hold133/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _8882_/X VGND VGND VPWR VPWR hold595/A sky130_fd_sc_hd__dlygate4sd3_1
X_5497_ _9438_/Q _5495_/A hold510/X _5495_/Y VGND VGND VPWR VPWR _5497_/X sky130_fd_sc_hd__a22o_1
X_7305_ _6134_/Y _7095_/B _6097_/Y _7157_/X VGND VGND VPWR VPWR _7305_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8285_ _8285_/A VGND VGND VPWR VPWR _8404_/B sky130_fd_sc_hd__inv_2
X_4517_ _9824_/Q _4513_/A _8959_/A1 _4513_/Y VGND VGND VPWR VPWR _9824_/D sky130_fd_sc_hd__a22o_1
Xhold176 hold176/A VGND VGND VPWR VPWR hold176/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold154 hold154/A VGND VGND VPWR VPWR _9356_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_171_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold165 hold165/A VGND VGND VPWR VPWR hold166/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7236_ _6384_/Y _7144_/X _6493_/Y _7145_/X _7235_/X VGND VGND VPWR VPWR _7243_/A
+ sky130_fd_sc_hd__o221a_1
Xhold198 hold198/A VGND VGND VPWR VPWR hold199/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold187 hold187/A VGND VGND VPWR VPWR _9510_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7167_ _7167_/A VGND VGND VPWR VPWR _7167_/X sky130_fd_sc_hd__buf_4
XFILLER_112_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6118_/A VGND VGND VPWR VPWR _6118_/Y sky130_fd_sc_hd__inv_2
X_7098_ _7108_/C _7128_/A _7127_/A VGND VGND VPWR VPWR _7136_/A sky130_fd_sc_hd__or3_2
XFILLER_58_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6049_ _8975_/A1 _9123_/Q _6049_/S VGND VGND VPWR VPWR _6050_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9808_ _9817_/CLK _9808_/D _9817_/SET_B VGND VGND VPWR VPWR _9808_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9739_ _9751_/CLK _9739_/D _5027_/X VGND VGND VPWR VPWR _9739_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9421_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_35_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9673_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5420_ _9491_/Q _5419_/A hold516/X _5419_/Y VGND VGND VPWR VPWR _5420_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput226 _8828_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_2
Xoutput215 _8808_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_133_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput204 _9813_/Q VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_2
X_5351_ _5474_/A _5351_/B VGND VGND VPWR VPWR _5352_/A sky130_fd_sc_hd__or2_1
Xoutput259 _9041_/Z VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_2
Xoutput237 _8877_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_2
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput248 _9031_/Z VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_2
X_8070_ _8666_/B _8592_/A VGND VGND VPWR VPWR _8070_/X sky130_fd_sc_hd__or2_1
X_5282_ _5282_/A _5282_/B VGND VGND VPWR VPWR _5283_/A sky130_fd_sc_hd__or2_1
X_7021_ _9751_/Q _6054_/Y _4975_/Y _9091_/Q VGND VGND VPWR VPWR _9091_/D sky130_fd_sc_hd__a31o_1
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8972_ _9660_/Q _8975_/A1 _8973_/S VGND VGND VPWR VPWR _8972_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7923_ _7942_/C _8234_/A _8625_/A VGND VGND VPWR VPWR _7924_/B sky130_fd_sc_hd__or3_2
X_7854_ _8383_/A VGND VGND VPWR VPWR _7873_/C sky130_fd_sc_hd__inv_2
XFILLER_23_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7785_ _7996_/C VGND VGND VPWR VPWR _8436_/B sky130_fd_sc_hd__buf_4
X_6805_ _9671_/Q VGND VGND VPWR VPWR _6805_/Y sky130_fd_sc_hd__inv_2
X_4997_ _5017_/A VGND VGND VPWR VPWR _4998_/A sky130_fd_sc_hd__clkbuf_1
X_9524_ _9550_/CLK _9524_/D _9537_/SET_B VGND VGND VPWR VPWR _9524_/Q sky130_fd_sc_hd__dfrtp_1
X_6736_ _9528_/Q VGND VGND VPWR VPWR _6736_/Y sky130_fd_sc_hd__clkinv_2
X_6667_ _7204_/A _5636_/B _6663_/Y _5620_/B _6666_/X VGND VGND VPWR VPWR _6680_/A
+ sky130_fd_sc_hd__o221a_1
X_9455_ _9579_/CLK _9455_/D _9727_/SET_B VGND VGND VPWR VPWR _9455_/Q sky130_fd_sc_hd__dfstp_1
X_5618_ _9355_/Q _5611_/A hold593/X _5611_/Y VGND VGND VPWR VPWR _9355_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9386_ _9522_/CLK _9386_/D _9537_/SET_B VGND VGND VPWR VPWR _9386_/Q sky130_fd_sc_hd__dfrtp_1
X_8406_ _8406_/A _8772_/C _8617_/C _8406_/D VGND VGND VPWR VPWR _8410_/A sky130_fd_sc_hd__or4_1
X_6598_ _6598_/A _6598_/B _6598_/C _6598_/D VGND VGND VPWR VPWR _6659_/A sky130_fd_sc_hd__and4_1
XFILLER_191_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8337_ _8337_/A _8337_/B VGND VGND VPWR VPWR _8338_/B sky130_fd_sc_hd__and2_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5549_ _9402_/Q _5545_/A _6067_/B1 _5545_/Y VGND VGND VPWR VPWR _9402_/D sky130_fd_sc_hd__a22o_1
XFILLER_191_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8268_ _8288_/A _8347_/B _8268_/C VGND VGND VPWR VPWR _8541_/B sky130_fd_sc_hd__nor3_1
XFILLER_105_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7219_ _8795_/A _7161_/X _8827_/A _7162_/X VGND VGND VPWR VPWR _7219_/X sky130_fd_sc_hd__o22a_1
X_8199_ _8199_/A _8672_/B VGND VGND VPWR VPWR _8201_/A sky130_fd_sc_hd__or2_1
XFILLER_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _4471_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_123_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4920_ _4920_/A _4953_/B VGND VGND VPWR VPWR _5367_/B sky130_fd_sc_hd__or2_4
X_4851_ _4843_/Y _4844_/X _4845_/Y _5123_/B _4850_/X VGND VGND VPWR VPWR _4852_/D
+ sky130_fd_sc_hd__o221a_1
X_7570_ _6452_/Y _7485_/X _6402_/Y _7486_/X _7569_/X VGND VGND VPWR VPWR _7586_/A
+ sky130_fd_sc_hd__o221a_1
X_4782_ _9227_/Q VGND VGND VPWR VPWR _4782_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6521_ _9138_/Q VGND VGND VPWR VPWR _7737_/A sky130_fd_sc_hd__inv_6
XFILLER_146_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6452_ _9418_/Q VGND VGND VPWR VPWR _6452_/Y sky130_fd_sc_hd__inv_2
X_9240_ _9431_/CLK _9240_/D _9797_/SET_B VGND VGND VPWR VPWR _9240_/Q sky130_fd_sc_hd__dfrtp_1
X_9171_ _9491_/CLK _9171_/D _9731_/SET_B VGND VGND VPWR VPWR _9171_/Q sky130_fd_sc_hd__dfrtp_1
X_5403_ _9501_/Q _5399_/A _6067_/B1 _5399_/Y VGND VGND VPWR VPWR _9501_/D sky130_fd_sc_hd__a22o_1
X_8122_ _8229_/B _8682_/B VGND VGND VPWR VPWR _8227_/A sky130_fd_sc_hd__or2_1
X_6383_ _6383_/A _6383_/B _6383_/C _6383_/D VGND VGND VPWR VPWR _6506_/A sky130_fd_sc_hd__and4_1
X_5334_ _9549_/Q _5331_/A hold577/A _5331_/Y VGND VGND VPWR VPWR _5334_/X sky130_fd_sc_hd__a22o_1
XFILLER_126_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8053_ _8053_/A _8053_/B VGND VGND VPWR VPWR _8053_/X sky130_fd_sc_hd__or2_1
XFILLER_125_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5265_ _5265_/A VGND VGND VPWR VPWR _5265_/Y sky130_fd_sc_hd__inv_2
X_5196_ _9640_/Q _5192_/A hold53/X _5192_/Y VGND VGND VPWR VPWR _9640_/D sky130_fd_sc_hd__a22o_1
X_7004_ _9103_/Q VGND VGND VPWR VPWR _7005_/A sky130_fd_sc_hd__inv_2
XFILLER_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8955_ _7762_/Y _9741_/Q _9090_/Q VGND VGND VPWR VPWR _8955_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8886_ hold261/X hold576/X _9629_/Q VGND VGND VPWR VPWR _8886_/X sky130_fd_sc_hd__mux2_8
X_7906_ _7999_/A _8570_/A _8625_/A _7933_/B VGND VGND VPWR VPWR _7907_/A sky130_fd_sc_hd__or4_4
X_7837_ _8436_/B _8134_/A VGND VGND VPWR VPWR _8065_/A sky130_fd_sc_hd__or2_4
XFILLER_70_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7768_ _9108_/Q _7768_/B VGND VGND VPWR VPWR _7768_/X sky130_fd_sc_hd__and2_1
XFILLER_177_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6719_ input45/X _8975_/S _6718_/Y _5866_/B VGND VGND VPWR VPWR _6719_/X sky130_fd_sc_hd__o2bb2a_2
X_9507_ _9561_/CLK _9507_/D _9817_/SET_B VGND VGND VPWR VPWR _9507_/Q sky130_fd_sc_hd__dfstp_1
X_7699_ _6574_/Y _7498_/A _6515_/Y _5727_/A VGND VGND VPWR VPWR _7699_/X sky130_fd_sc_hd__o22a_1
X_9438_ _9522_/CLK _9438_/D _9537_/SET_B VGND VGND VPWR VPWR _9438_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9369_ _9421_/CLK _9369_/D _9537_/SET_B VGND VGND VPWR VPWR _9369_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold709 _9187_/Q VGND VGND VPWR VPWR hold709/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5050_ _9729_/Q _5049_/A _6064_/B1 _5049_/Y VGND VGND VPWR VPWR _9729_/D sky130_fd_sc_hd__a22o_1
XFILLER_111_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8740_ _8740_/A _8750_/A _7970_/A VGND VGND VPWR VPWR _8741_/B sky130_fd_sc_hd__or3b_1
XFILLER_92_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5952_ _9163_/Q _5948_/A _8969_/A1 _5948_/Y VGND VGND VPWR VPWR _9163_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4903_ _4896_/Y _4623_/B _4897_/Y _5133_/B _4902_/X VGND VGND VPWR VPWR _4918_/B
+ sky130_fd_sc_hd__o221a_1
X_8671_ _8752_/A _8671_/B _8728_/D _8670_/X VGND VGND VPWR VPWR _8675_/A sky130_fd_sc_hd__or4b_1
XFILLER_21_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5883_ _5878_/X _8906_/X _8960_/X _9214_/Q VGND VGND VPWR VPWR _9214_/D sky130_fd_sc_hd__o22a_1
X_7622_ _7622_/A _7622_/B _7622_/C _7622_/D VGND VGND VPWR VPWR _7622_/Y sky130_fd_sc_hd__nand4_4
XFILLER_21_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4834_ _4822_/Y _5313_/B _4826_/Y _5559_/B _4833_/X VGND VGND VPWR VPWR _4852_/B
+ sky130_fd_sc_hd__o221a_1
X_4765_ _9432_/Q VGND VGND VPWR VPWR _4765_/Y sky130_fd_sc_hd__clkinv_4
X_7553_ _8785_/A _7493_/X _8823_/A _7494_/X VGND VGND VPWR VPWR _7553_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6504_ _6504_/A _6504_/B _6504_/C _6504_/D VGND VGND VPWR VPWR _6505_/D sky130_fd_sc_hd__and4_1
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9223_ _9420_/CLK _9223_/D _9537_/SET_B VGND VGND VPWR VPWR _9223_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4696_ _4808_/A _4900_/A VGND VGND VPWR VPWR _5532_/B sky130_fd_sc_hd__or2_4
X_7484_ _7484_/A VGND VGND VPWR VPWR _7484_/X sky130_fd_sc_hd__clkbuf_1
X_6435_ _9431_/Q VGND VGND VPWR VPWR _6435_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_161_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9154_ _9736_/CLK _9154_/D _9731_/SET_B VGND VGND VPWR VPWR _9154_/Q sky130_fd_sc_hd__dfrtp_1
X_6366_ _9426_/Q VGND VGND VPWR VPWR _6366_/Y sky130_fd_sc_hd__inv_2
X_9085_ _9705_/CLK _9085_/D VGND VGND VPWR VPWR _9085_/Q sky130_fd_sc_hd__dfxtp_1
X_8105_ _8560_/A _8105_/B _8105_/C VGND VGND VPWR VPWR _8745_/C sky130_fd_sc_hd__and3_1
XFILLER_0_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5317_ _9560_/Q _5315_/A _6065_/B1 _5315_/Y VGND VGND VPWR VPWR _9560_/D sky130_fd_sc_hd__a22o_1
X_8036_ _8169_/A VGND VGND VPWR VPWR _8171_/B sky130_fd_sc_hd__buf_2
Xhold14 hold14/A VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6297_ _6295_/Y _5455_/B _6296_/Y _4623_/B VGND VGND VPWR VPWR _6297_/X sky130_fd_sc_hd__o22a_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _9604_/Q _5241_/Y _8974_/X hold689/X VGND VGND VPWR VPWR _9604_/D sky130_fd_sc_hd__o22a_1
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold25 hold25/A VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5179_ _6166_/A _5179_/B VGND VGND VPWR VPWR _5180_/A sky130_fd_sc_hd__or2_2
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8938_ _8937_/X hold705/X _9096_/Q VGND VGND VPWR VPWR _8938_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8869_ _8868_/X _7051_/B _9628_/Q VGND VGND VPWR VPWR _8869_/X sky130_fd_sc_hd__mux2_4
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4550_ _9809_/Q _4547_/A hold696/X _4547_/Y VGND VGND VPWR VPWR _9809_/D sky130_fd_sc_hd__a22o_1
XFILLER_183_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold517 hold517/A VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__clkbuf_2
X_4481_ _4750_/A _4750_/B _4750_/C _4642_/B VGND VGND VPWR VPWR _4866_/A sky130_fd_sc_hd__or4_4
Xhold506 hold506/A VGND VGND VPWR VPWR hold507/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold539 _5371_/X VGND VGND VPWR VPWR _9524_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold528 _5691_/X VGND VGND VPWR VPWR _9317_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6220_ _9826_/Q VGND VGND VPWR VPWR _6220_/Y sky130_fd_sc_hd__inv_4
X_6151_ _9737_/Q VGND VGND VPWR VPWR _6151_/Y sky130_fd_sc_hd__clkinv_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A VGND VGND VPWR VPWR _9701_/D sky130_fd_sc_hd__clkbuf_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6082_/A VGND VGND VPWR VPWR _6082_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A VGND VGND VPWR VPWR _5033_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6984_ _6176_/Y _6983_/A _9077_/Q _6983_/Y VGND VGND VPWR VPWR _9077_/D sky130_fd_sc_hd__o22a_1
X_9772_ _9817_/CLK _9772_/D _9817_/SET_B VGND VGND VPWR VPWR _9772_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8723_ _8723_/A _8723_/B _8723_/C VGND VGND VPWR VPWR _8765_/A sky130_fd_sc_hd__or3_1
X_5935_ _6083_/A _5935_/B VGND VGND VPWR VPWR _5936_/A sky130_fd_sc_hd__or2_1
X_5866_ _6083_/A _5866_/B VGND VGND VPWR VPWR _5867_/A sky130_fd_sc_hd__or2_1
X_8654_ _8654_/A _8654_/B VGND VGND VPWR VPWR _8708_/D sky130_fd_sc_hd__or2_1
XFILLER_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7605_ _6227_/Y _7487_/X _6261_/Y _7488_/X VGND VGND VPWR VPWR _7605_/X sky130_fd_sc_hd__o22a_1
X_4817_ _9669_/Q VGND VGND VPWR VPWR _4817_/Y sky130_fd_sc_hd__inv_2
X_8585_ _8585_/A VGND VGND VPWR VPWR _8585_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5797_ _5990_/A _5797_/B VGND VGND VPWR VPWR _5798_/A sky130_fd_sc_hd__or2_1
XFILLER_193_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7536_ _6670_/Y _7491_/X _6712_/Y _7492_/X _7535_/X VGND VGND VPWR VPWR _7550_/B
+ sky130_fd_sc_hd__o221a_1
X_4748_ _4920_/A _4801_/B VGND VGND VPWR VPWR _5687_/B sky130_fd_sc_hd__or2_4
XFILLER_174_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4679_ _9133_/Q _9132_/Q _9134_/Q VGND VGND VPWR VPWR _7034_/C sky130_fd_sc_hd__or3_2
X_7467_ _7467_/A _7473_/A _9297_/Q VGND VGND VPWR VPWR _7516_/A sky130_fd_sc_hd__or3_2
X_6418_ _9530_/Q VGND VGND VPWR VPWR _6418_/Y sky130_fd_sc_hd__clkinv_2
X_9206_ _9319_/CLK _9206_/D _9797_/SET_B VGND VGND VPWR VPWR _9206_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9137_ _9574_/CLK _9137_/D _9571_/SET_B VGND VGND VPWR VPWR _9137_/Q sky130_fd_sc_hd__dfrtp_1
X_7398_ _6515_/Y _7167_/A _6559_/Y _7168_/A VGND VGND VPWR VPWR _7398_/X sky130_fd_sc_hd__o22a_1
XFILLER_163_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6349_ _6347_/Y _5687_/B _6348_/Y _6165_/A VGND VGND VPWR VPWR _6349_/X sky130_fd_sc_hd__o22a_1
XFILLER_103_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9068_ _9723_/CLK _9068_/D VGND VGND VPWR VPWR _9068_/Q sky130_fd_sc_hd__dfxtp_1
Xinput126 uart_enabled VGND VGND VPWR VPWR _8843_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput104 sram_ro_data[1] VGND VGND VPWR VPWR _6851_/A sky130_fd_sc_hd__clkbuf_1
Xinput115 sram_ro_data[2] VGND VGND VPWR VPWR _6710_/A sky130_fd_sc_hd__clkbuf_1
Xinput148 wb_adr_i[24] VGND VGND VPWR VPWR _5955_/C sky130_fd_sc_hd__clkbuf_1
Xinput137 wb_adr_i[14] VGND VGND VPWR VPWR _7805_/B sky130_fd_sc_hd__clkbuf_1
Xinput159 wb_adr_i[5] VGND VGND VPWR VPWR _8567_/A sky130_fd_sc_hd__buf_6
X_8019_ _8019_/A VGND VGND VPWR VPWR _8034_/A sky130_fd_sc_hd__inv_2
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5720_ _9294_/Q _9293_/Q VGND VGND VPWR VPWR _7460_/A sky130_fd_sc_hd__or2_1
XFILLER_50_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5651_ _9334_/Q _5649_/A hold510/X _5649_/Y VGND VGND VPWR VPWR _5651_/X sky130_fd_sc_hd__a22o_1
X_8370_ _7887_/A _8342_/B _8369_/Y VGND VGND VPWR VPWR _8371_/C sky130_fd_sc_hd__o21ai_1
X_4602_ _9788_/Q _4600_/A hold510/X _4600_/Y VGND VGND VPWR VPWR _9788_/D sky130_fd_sc_hd__a22o_1
X_5582_ _5582_/A VGND VGND VPWR VPWR _5583_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4533_ _9814_/Q _4485_/A _8959_/A1 _4485_/Y VGND VGND VPWR VPWR _9814_/D sky130_fd_sc_hd__a22o_1
X_7321_ _4752_/A _7137_/X _4691_/Y _7138_/X _7320_/X VGND VGND VPWR VPWR _7321_/X
+ sky130_fd_sc_hd__o221a_1
Xhold325 hold325/A VGND VGND VPWR VPWR hold326/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 hold314/A VGND VGND VPWR VPWR _9541_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold303 _5449_/X VGND VGND VPWR VPWR hold304/A sky130_fd_sc_hd__dlygate4sd3_1
X_7252_ _7252_/A _7252_/B _7252_/C _7252_/D VGND VGND VPWR VPWR _7253_/C sky130_fd_sc_hd__and4_1
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4464_ _9630_/Q input80/X _8875_/S VGND VGND VPWR VPWR _9051_/A sky130_fd_sc_hd__mux2_1
Xhold336 _5871_/X VGND VGND VPWR VPWR hold337/A sky130_fd_sc_hd__dlygate4sd3_1
X_6203_ _6201_/Y _5647_/B _6202_/Y _4869_/X VGND VGND VPWR VPWR _6203_/X sky130_fd_sc_hd__o22a_1
Xhold358 hold358/A VGND VGND VPWR VPWR hold359/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _8977_/X VGND VGND VPWR VPWR hold370/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 hold347/A VGND VGND VPWR VPWR _9813_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7183_ _7183_/A VGND VGND VPWR VPWR _7183_/X sky130_fd_sc_hd__buf_6
X_6134_ _9465_/Q VGND VGND VPWR VPWR _6134_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _9115_/Q _6060_/A _6065_/B1 _6060_/Y VGND VGND VPWR VPWR _9115_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5016_/A VGND VGND VPWR VPWR _9742_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9824_ _9827_/CLK _9824_/D _9797_/SET_B VGND VGND VPWR VPWR _9824_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _7358_/A _5658_/B _6966_/Y _5797_/B VGND VGND VPWR VPWR _6967_/X sky130_fd_sc_hd__o22a_1
X_9755_ net399_3/A _9755_/D _4672_/X VGND VGND VPWR VPWR _9755_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8706_ _8706_/A VGND VGND VPWR VPWR _8706_/X sky130_fd_sc_hd__clkbuf_1
X_5918_ _5889_/X _8928_/X _8960_/X _9187_/Q VGND VGND VPWR VPWR _9187_/D sky130_fd_sc_hd__o22a_1
X_9686_ _9686_/CLK _9686_/D _9817_/SET_B VGND VGND VPWR VPWR _9686_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6898_ _9454_/Q VGND VGND VPWR VPWR _6898_/Y sky130_fd_sc_hd__clkinv_2
X_5849_ _5849_/A VGND VGND VPWR VPWR _5849_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8637_ _8637_/A _8637_/B _8637_/C _7941_/X VGND VGND VPWR VPWR _8701_/C sky130_fd_sc_hd__or4b_1
XFILLER_42_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8568_ _8567_/Y _8559_/Y _8560_/X _8491_/A VGND VGND VPWR VPWR _8708_/A sky130_fd_sc_hd__a31o_1
XFILLER_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7519_ _7519_/A VGND VGND VPWR VPWR _7519_/X sky130_fd_sc_hd__buf_6
X_8499_ _8563_/B _8288_/B _8070_/X VGND VGND VPWR VPWR _8501_/C sky130_fd_sc_hd__o21ai_1
XFILLER_162_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7870_ _7870_/A VGND VGND VPWR VPWR _8268_/C sky130_fd_sc_hd__buf_6
X_6821_ _9805_/Q VGND VGND VPWR VPWR _6821_/Y sky130_fd_sc_hd__inv_2
X_9540_ _9576_/CLK _9540_/D _9537_/SET_B VGND VGND VPWR VPWR _9540_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6752_ _6750_/Y _5474_/B _6751_/Y _5455_/B VGND VGND VPWR VPWR _6752_/X sky130_fd_sc_hd__o22a_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9471_ _9577_/CLK _9471_/D _9571_/SET_B VGND VGND VPWR VPWR _9471_/Q sky130_fd_sc_hd__dfrtp_1
X_5703_ _9308_/Q _5700_/A hold217/X _5700_/Y VGND VGND VPWR VPWR _9308_/D sky130_fd_sc_hd__a22o_1
X_6683_ _9817_/Q VGND VGND VPWR VPWR _6683_/Y sky130_fd_sc_hd__clkinv_4
X_8422_ _8422_/A _8422_/B _8762_/C _8627_/A VGND VGND VPWR VPWR _8423_/B sky130_fd_sc_hd__or4_1
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5634_ _9345_/Q _5630_/A _6067_/B1 _5630_/Y VGND VGND VPWR VPWR _9345_/D sky130_fd_sc_hd__a22o_1
XFILLER_191_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8353_ _8682_/A _8353_/B VGND VGND VPWR VPWR _8634_/A sky130_fd_sc_hd__or2_2
XFILLER_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold100 hold99/X VGND VGND VPWR VPWR hold101/A sky130_fd_sc_hd__dlygate4sd3_1
X_5565_ _9392_/Q _5561_/A hold53/X _5561_/Y VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__a22o_1
X_7304_ _6109_/Y _7149_/X _6153_/Y _7150_/X _7303_/X VGND VGND VPWR VPWR _7309_/B
+ sky130_fd_sc_hd__o221a_1
Xhold144 hold144/A VGND VGND VPWR VPWR hold145/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 hold133/A VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold122 hold595/X VGND VGND VPWR VPWR hold594/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _5853_/X VGND VGND VPWR VPWR hold112/A sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ _9439_/Q _5495_/A hold516/X _5495_/Y VGND VGND VPWR VPWR _5496_/X sky130_fd_sc_hd__a22o_1
X_8284_ _8552_/A _8288_/B VGND VGND VPWR VPWR _8285_/A sky130_fd_sc_hd__or2_2
X_4516_ _9825_/Q _4513_/A hold696/A _4513_/Y VGND VGND VPWR VPWR _4516_/X sky130_fd_sc_hd__a22o_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold177 hold603/X VGND VGND VPWR VPWR hold602/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _5187_/X VGND VGND VPWR VPWR hold156/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 hold166/A VGND VGND VPWR VPWR _9460_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7235_ _6494_/Y _7071_/C _6368_/Y _7146_/X VGND VGND VPWR VPWR _7235_/X sky130_fd_sc_hd__o22a_1
Xhold199 hold199/A VGND VGND VPWR VPWR hold199/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold188 _9748_/Q VGND VGND VPWR VPWR hold189/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7166_ _7166_/A VGND VGND VPWR VPWR _7166_/X sky130_fd_sc_hd__buf_4
XFILLER_100_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6117_ _6117_/A _6117_/B VGND VGND VPWR VPWR _6117_/X sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_1_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9483_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7108_/C _7129_/A _7127_/A VGND VGND VPWR VPWR _7135_/A sky130_fd_sc_hd__or3_2
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6048_ _9124_/Q _6026_/A _8949_/X _6026_/Y VGND VGND VPWR VPWR _9124_/D sky130_fd_sc_hd__a22o_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9807_ _9810_/CLK _9807_/D _7042_/B VGND VGND VPWR VPWR _9807_/Q sky130_fd_sc_hd__dfrtp_4
X_7999_ _7999_/A _8005_/A _8006_/B VGND VGND VPWR VPWR _8234_/B sky130_fd_sc_hd__or3_2
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9738_ _9751_/CLK _9738_/D _5033_/X VGND VGND VPWR VPWR _9738_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9669_ _9832_/CLK _9669_/D _9797_/SET_B VGND VGND VPWR VPWR _9669_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _8879_/A1
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput216 _8810_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_2
X_5350_ _9536_/Q _5342_/A hold601/X _5342_/Y VGND VGND VPWR VPWR _5350_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput205 _8849_/Y VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput227 _8830_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_141_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput249 _9032_/Z VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_2
X_5281_ _9583_/Q _5276_/A _8975_/A1 _5276_/Y VGND VGND VPWR VPWR _9583_/D sky130_fd_sc_hd__a22o_1
Xoutput238 _7738_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_2
X_7020_ _8855_/A _8851_/A _6981_/B VGND VGND VPWR VPWR _7020_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_141_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8971_ _9659_/Q hold516/X _8971_/S VGND VGND VPWR VPWR _8971_/X sky130_fd_sc_hd__mux2_1
X_7922_ _8439_/A VGND VGND VPWR VPWR _7925_/B sky130_fd_sc_hd__inv_2
XFILLER_82_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7853_ _8243_/A _8138_/B VGND VGND VPWR VPWR _8135_/A sky130_fd_sc_hd__or2_1
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6804_ _9690_/Q VGND VGND VPWR VPWR _6804_/Y sky130_fd_sc_hd__inv_4
X_4996_ _9747_/Q _4989_/A hold46/A _4989_/Y VGND VGND VPWR VPWR _9747_/D sky130_fd_sc_hd__a22o_1
XFILLER_168_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7784_ _8421_/B VGND VGND VPWR VPWR _7996_/C sky130_fd_sc_hd__inv_2
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9523_ _9550_/CLK _9523_/D _9563_/SET_B VGND VGND VPWR VPWR _9523_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6735_ _9512_/Q VGND VGND VPWR VPWR _6735_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9454_ _9579_/CLK _9454_/D _9727_/SET_B VGND VGND VPWR VPWR _9454_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6666_ _6664_/Y _5687_/B _6665_/Y _5698_/B VGND VGND VPWR VPWR _6666_/X sky130_fd_sc_hd__o22a_1
XFILLER_191_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5617_ _9356_/Q _5611_/A hold136/X _5611_/Y VGND VGND VPWR VPWR _5617_/X sky130_fd_sc_hd__a22o_1
X_9385_ _9522_/CLK _9385_/D _9537_/SET_B VGND VGND VPWR VPWR _9385_/Q sky130_fd_sc_hd__dfrtp_1
X_8405_ _8669_/B _8532_/B VGND VGND VPWR VPWR _8406_/D sky130_fd_sc_hd__or2_1
X_6597_ _6592_/Y _4854_/X _8833_/A _5378_/B _6596_/X VGND VGND VPWR VPWR _6598_/D
+ sky130_fd_sc_hd__o221a_1
X_8336_ _8336_/A _8692_/C VGND VGND VPWR VPWR _8337_/B sky130_fd_sc_hd__or2_1
XFILLER_151_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5548_ _9403_/Q _5545_/A hold217/X _5545_/Y VGND VGND VPWR VPWR _9403_/D sky130_fd_sc_hd__a22o_1
XFILLER_151_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8267_ _8347_/B _8302_/B VGND VGND VPWR VPWR _8613_/B sky130_fd_sc_hd__nor2_2
XFILLER_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7218_ _6613_/Y _7155_/X _8839_/A _7156_/X _7217_/X VGND VGND VPWR VPWR _7221_/C
+ sky130_fd_sc_hd__o221a_1
X_5479_ _9450_/Q _5476_/A hold217/X _5476_/Y VGND VGND VPWR VPWR _9450_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8198_ _8205_/A _8596_/A VGND VGND VPWR VPWR _8672_/B sky130_fd_sc_hd__nor2_1
XFILLER_48_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7149_ _7149_/A VGND VGND VPWR VPWR _7149_/X sky130_fd_sc_hd__buf_6
XFILLER_171_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4850_ _8849_/A _4848_/X _4849_/Y _6282_/A VGND VGND VPWR VPWR _4850_/X sky130_fd_sc_hd__o22a_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6520_ _9435_/Q VGND VGND VPWR VPWR _8839_/A sky130_fd_sc_hd__inv_4
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4781_ _4949_/A _4801_/B VGND VGND VPWR VPWR _5636_/B sky130_fd_sc_hd__or2_4
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6451_ _6446_/Y _5406_/B _6447_/Y _5971_/B _6450_/X VGND VGND VPWR VPWR _6464_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_173_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9170_ _9491_/CLK _9170_/D _9731_/SET_B VGND VGND VPWR VPWR _9170_/Q sky130_fd_sc_hd__dfrtp_1
X_5402_ _9502_/Q _5399_/A hold217/X _5399_/Y VGND VGND VPWR VPWR _9502_/D sky130_fd_sc_hd__a22o_1
X_6382_ _6377_/Y _4869_/X _6378_/Y _5351_/B _6381_/X VGND VGND VPWR VPWR _6383_/D
+ sky130_fd_sc_hd__o221a_1
X_8121_ _8153_/A VGND VGND VPWR VPWR _8682_/B sky130_fd_sc_hd__buf_8
X_5333_ _9550_/Q _5331_/A hold510/X _5331_/Y VGND VGND VPWR VPWR _5333_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8052_ _8565_/A _8559_/A VGND VGND VPWR VPWR _8053_/B sky130_fd_sc_hd__or2_1
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5264_ _5264_/A VGND VGND VPWR VPWR _5265_/A sky130_fd_sc_hd__clkbuf_4
X_5195_ _9641_/Q _5192_/A hold577/A _5192_/Y VGND VGND VPWR VPWR _5195_/X sky130_fd_sc_hd__a22o_1
X_7003_ _4958_/Y _6995_/A _9062_/Q _6995_/Y VGND VGND VPWR VPWR _9062_/D sky130_fd_sc_hd__o22a_1
XFILLER_83_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8954_ _7760_/X _9740_/Q _9090_/Q VGND VGND VPWR VPWR _8954_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8885_ hold49/X hold656/X _9629_/Q VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__mux2_8
X_7905_ _7905_/A VGND VGND VPWR VPWR _8361_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7836_ _8421_/C _7876_/A _8421_/D VGND VGND VPWR VPWR _8134_/A sky130_fd_sc_hd__or3_4
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7767_ _9109_/Q _5081_/X _7765_/X _7766_/X VGND VGND VPWR VPWR _7767_/X sky130_fd_sc_hd__a211o_1
X_4979_ _5017_/A VGND VGND VPWR VPWR _4980_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6718_ _9221_/Q VGND VGND VPWR VPWR _6718_/Y sky130_fd_sc_hd__clkinv_2
X_9506_ _9561_/CLK _9506_/D _9817_/SET_B VGND VGND VPWR VPWR _9506_/Q sky130_fd_sc_hd__dfrtp_1
X_7698_ _6612_/Y _7491_/A _6570_/Y _7492_/A _7697_/X VGND VGND VPWR VPWR _7712_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_164_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9437_ _9522_/CLK _9437_/D _9537_/SET_B VGND VGND VPWR VPWR _9437_/Q sky130_fd_sc_hd__dfrtp_1
X_6649_ _6649_/A VGND VGND VPWR VPWR _6649_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9368_ _9643_/CLK _9368_/D _9563_/SET_B VGND VGND VPWR VPWR _9368_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_34_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9833_/CLK sky130_fd_sc_hd__clkbuf_16
X_9299_ _9392_/CLK _9299_/D _9689_/SET_B VGND VGND VPWR VPWR _9299_/Q sky130_fd_sc_hd__dfstp_1
X_8319_ _8567_/A _7904_/D _8243_/B _8625_/A _8230_/Y VGND VGND VPWR VPWR _8387_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_145_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_49_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9582_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_1_mgmt_gpio_in[4] clkbuf_1_0_1_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR clkbuf_2_1_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_2
X_5951_ _9164_/Q _5948_/A _8965_/A1 _5948_/Y VGND VGND VPWR VPWR _9164_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8670_ _8171_/B _8596_/B _8496_/B _8174_/A _8450_/Y VGND VGND VPWR VPWR _8670_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_92_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4902_ _4899_/Y _5521_/B _4901_/Y _4536_/X VGND VGND VPWR VPWR _4902_/X sky130_fd_sc_hd__o22a_1
X_5882_ _5878_/X _8908_/X _8960_/X _9215_/Q VGND VGND VPWR VPWR _9215_/D sky130_fd_sc_hd__o22a_1
X_7621_ _7621_/A _7621_/B _7621_/C _7621_/D VGND VGND VPWR VPWR _7622_/D sky130_fd_sc_hd__and4_2
XFILLER_21_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4833_ _4953_/A _6189_/A _4830_/Y _4831_/Y _5274_/B VGND VGND VPWR VPWR _4833_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_119_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7552_ _8817_/A _7487_/X _7737_/A _7488_/X _7551_/X VGND VGND VPWR VPWR _7568_/A
+ sky130_fd_sc_hd__o221a_1
X_4764_ _4898_/B _4764_/B VGND VGND VPWR VPWR _5598_/B sky130_fd_sc_hd__or2_4
XFILLER_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6503_ _6498_/Y _5858_/B _6499_/Y _5902_/B _6502_/X VGND VGND VPWR VPWR _6504_/D
+ sky130_fd_sc_hd__o221a_1
X_7483_ _7483_/A _7483_/B _7483_/C _7483_/D VGND VGND VPWR VPWR _7484_/A sky130_fd_sc_hd__and4_1
X_4695_ _9406_/Q VGND VGND VPWR VPWR _4695_/Y sky130_fd_sc_hd__clkinv_4
X_9222_ _9421_/CLK _9222_/D _9537_/SET_B VGND VGND VPWR VPWR _9222_/Q sky130_fd_sc_hd__dfrtp_1
X_6434_ _9824_/Q VGND VGND VPWR VPWR _6434_/Y sky130_fd_sc_hd__inv_4
XFILLER_161_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9153_ _9736_/CLK _9153_/D _9731_/SET_B VGND VGND VPWR VPWR _9153_/Q sky130_fd_sc_hd__dfrtp_1
X_6365_ _9139_/Q VGND VGND VPWR VPWR _6365_/Y sky130_fd_sc_hd__inv_2
X_9084_ _9705_/CLK _9084_/D VGND VGND VPWR VPWR _9084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8104_ _8118_/A VGND VGND VPWR VPWR _8560_/A sky130_fd_sc_hd__inv_2
X_6296_ _9773_/Q VGND VGND VPWR VPWR _6296_/Y sky130_fd_sc_hd__inv_2
X_5316_ _9561_/Q _5315_/A _6064_/B1 _5315_/Y VGND VGND VPWR VPWR _9561_/D sky130_fd_sc_hd__a22o_1
X_5247_ _9605_/Q _5241_/Y hold199/X _5241_/A VGND VGND VPWR VPWR _5247_/X sky130_fd_sc_hd__o22a_1
X_8035_ _8157_/B _8035_/B VGND VGND VPWR VPWR _8169_/A sky130_fd_sc_hd__or2_1
XFILLER_102_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold37 hold37/A VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold26 hold26/A VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5178_ _9652_/Q _5170_/A _8975_/A1 _5170_/Y VGND VGND VPWR VPWR _9652_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8937_ _7429_/Y _9673_/Q _9001_/S VGND VGND VPWR VPWR _8937_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8868_ _8867_/X _6536_/A _9724_/Q VGND VGND VPWR VPWR _8868_/X sky130_fd_sc_hd__mux2_1
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7819_ _7936_/A _7937_/B VGND VGND VPWR VPWR _8125_/A sky130_fd_sc_hd__or2_2
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8799_ _8799_/A VGND VGND VPWR VPWR _8800_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold518 _8888_/X VGND VGND VPWR VPWR hold518/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_167_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4480_ _4708_/B VGND VGND VPWR VPWR _4750_/B sky130_fd_sc_hd__clkinv_2
Xhold507 hold507/A VGND VGND VPWR VPWR _4823_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_7_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold529 _5830_/X VGND VGND VPWR VPWR _9252_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6150_ _6150_/A _6150_/B _6150_/C _6150_/D VGND VGND VPWR VPWR _6176_/C sky130_fd_sc_hd__and4_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _9003_/X _9701_/Q _5101_/S VGND VGND VPWR VPWR _5102_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6081_/A VGND VGND VPWR VPWR _6082_/A sky130_fd_sc_hd__clkbuf_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _6017_/A VGND VGND VPWR VPWR _5033_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_122_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6983_ _6983_/A VGND VGND VPWR VPWR _6983_/Y sky130_fd_sc_hd__clkinv_2
X_9771_ _9817_/CLK _9771_/D _9821_/SET_B VGND VGND VPWR VPWR _9771_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8722_ _8758_/D _8773_/D _8722_/C _8762_/A VGND VGND VPWR VPWR _8722_/Y sky130_fd_sc_hd__nor4_1
X_5934_ _9175_/Q _5929_/A _8975_/A1 _5929_/Y VGND VGND VPWR VPWR _9175_/D sky130_fd_sc_hd__a22o_1
X_8653_ _8105_/C _8652_/Y _8056_/A _8569_/B VGND VGND VPWR VPWR _8655_/B sky130_fd_sc_hd__a211o_1
X_5865_ _9227_/Q _5860_/A _8975_/A1 _5860_/Y VGND VGND VPWR VPWR _9227_/D sky130_fd_sc_hd__a22o_1
XFILLER_178_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7604_ _7604_/A _7604_/B _7604_/C _7604_/D VGND VGND VPWR VPWR _7604_/Y sky130_fd_sc_hd__nand4_4
X_4816_ _4933_/A _4951_/A VGND VGND VPWR VPWR _5263_/B sky130_fd_sc_hd__or2_4
XFILLER_193_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5796_ _9273_/Q _5788_/A _8975_/A1 _5788_/Y VGND VGND VPWR VPWR _9273_/D sky130_fd_sc_hd__a22o_1
X_8584_ _8745_/B _8647_/A _8747_/A _8583_/Y VGND VGND VPWR VPWR _8585_/A sky130_fd_sc_hd__or4b_1
XFILLER_119_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4747_ _9311_/Q VGND VGND VPWR VPWR _4747_/Y sky130_fd_sc_hd__inv_2
X_7535_ _6698_/Y _7493_/X _6723_/Y _7494_/X VGND VGND VPWR VPWR _7535_/X sky130_fd_sc_hd__o22a_1
XFILLER_31_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4678_ _4678_/A VGND VGND VPWR VPWR _4678_/X sky130_fd_sc_hd__clkbuf_1
X_7466_ _7467_/A _7473_/A _7478_/D VGND VGND VPWR VPWR _7515_/A sky130_fd_sc_hd__or3_2
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9205_ _9574_/CLK _9205_/D _9571_/SET_B VGND VGND VPWR VPWR _9205_/Q sky130_fd_sc_hd__dfrtp_1
X_6417_ input7/X VGND VGND VPWR VPWR _6417_/Y sky130_fd_sc_hd__inv_2
X_7397_ _7397_/A _7397_/B _7397_/C _7397_/D VGND VGND VPWR VPWR _7407_/B sky130_fd_sc_hd__and4_1
X_6348_ _6348_/A VGND VGND VPWR VPWR _6348_/Y sky130_fd_sc_hd__inv_2
X_9136_ _9574_/CLK _9136_/D _9571_/SET_B VGND VGND VPWR VPWR _9136_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_88_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput127 user_clock VGND VGND VPWR VPWR _4470_/A1 sky130_fd_sc_hd__buf_2
X_9067_ _9723_/CLK _9067_/D VGND VGND VPWR VPWR _9067_/Q sky130_fd_sc_hd__dfxtp_1
X_6279_ _6274_/Y _4598_/B _6275_/Y _5340_/B _6278_/X VGND VGND VPWR VPWR _6279_/X
+ sky130_fd_sc_hd__o221a_2
Xinput116 sram_ro_data[30] VGND VGND VPWR VPWR _6258_/A sky130_fd_sc_hd__clkbuf_1
Xinput105 sram_ro_data[20] VGND VGND VPWR VPWR _6469_/A sky130_fd_sc_hd__clkbuf_1
Xinput149 wb_adr_i[25] VGND VGND VPWR VPWR input149/X sky130_fd_sc_hd__clkbuf_1
Xinput138 wb_adr_i[15] VGND VGND VPWR VPWR _7805_/A sky130_fd_sc_hd__clkbuf_1
X_8018_ _8137_/A _8139_/A VGND VGND VPWR VPWR _8035_/B sky130_fd_sc_hd__or2_1
X_8857__412 VGND VGND VPWR VPWR _9099_/D _8857__412/LO sky130_fd_sc_hd__conb_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5650_ _9335_/Q _5649_/A hold516/X _5649_/Y VGND VGND VPWR VPWR _5650_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4601_ _9789_/Q _4600_/A hold516/X _4600_/Y VGND VGND VPWR VPWR _9789_/D sky130_fd_sc_hd__a22o_1
X_5581_ _5698_/A _5581_/B VGND VGND VPWR VPWR _5582_/A sky130_fd_sc_hd__or2_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4532_ _9815_/Q _4527_/A _6008_/B1 _4527_/Y VGND VGND VPWR VPWR _4532_/X sky130_fd_sc_hd__a22o_1
X_7320_ _4921_/Y _7139_/X _4870_/Y _7140_/X VGND VGND VPWR VPWR _7320_/X sky130_fd_sc_hd__o22a_1
Xhold326 hold326/A VGND VGND VPWR VPWR _9251_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold304 hold304/A VGND VGND VPWR VPWR hold305/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 _5295_/X VGND VGND VPWR VPWR hold316/A sky130_fd_sc_hd__dlygate4sd3_1
X_7251_ _6359_/Y _7180_/X _6441_/Y _7181_/X _7250_/X VGND VGND VPWR VPWR _7252_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold337 hold337/A VGND VGND VPWR VPWR hold338/A sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _9576_/Q VGND VGND VPWR VPWR _6202_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold348 _9717_/Q VGND VGND VPWR VPWR hold349/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold359 hold359/A VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_131_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7182_ _7182_/A VGND VGND VPWR VPWR _7182_/X sky130_fd_sc_hd__buf_6
XFILLER_97_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6133_ _6128_/Y _4854_/X _6129_/Y _5559_/B _6132_/X VGND VGND VPWR VPWR _6150_/A
+ sky130_fd_sc_hd__o221a_2
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6064_ _9116_/Q _6060_/A _6064_/B1 _6060_/Y VGND VGND VPWR VPWR _6064_/X sky130_fd_sc_hd__a22o_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _8955_/X _9742_/Q _5024_/S VGND VGND VPWR VPWR _5016_/A sky130_fd_sc_hd__mux2_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9823_ _9832_/CLK _9823_/D _9821_/SET_B VGND VGND VPWR VPWR _9823_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9754_ net399_3/A _9754_/D _4675_/X VGND VGND VPWR VPWR _9754_/Q sky130_fd_sc_hd__dfrtn_1
X_6966_ _9269_/Q VGND VGND VPWR VPWR _6966_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8705_ _8738_/C _8769_/C _8705_/C _8763_/A VGND VGND VPWR VPWR _8706_/A sky130_fd_sc_hd__or4_1
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5917_ _5889_/X _8930_/X _8960_/X _9188_/Q VGND VGND VPWR VPWR _9188_/D sky130_fd_sc_hd__o22a_1
X_9685_ _9819_/CLK _9685_/D _9817_/SET_B VGND VGND VPWR VPWR _9685_/Q sky130_fd_sc_hd__dfrtp_1
X_6897_ _9506_/Q VGND VGND VPWR VPWR _6897_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5848_ _5848_/A VGND VGND VPWR VPWR _5849_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_139_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8636_ _8636_/A _8636_/B _7935_/X VGND VGND VPWR VPWR _8637_/A sky130_fd_sc_hd__or3b_1
X_8567_ _8567_/A _8580_/B _8567_/C VGND VGND VPWR VPWR _8567_/Y sky130_fd_sc_hd__nor3_4
X_5779_ _9098_/Q _8861_/X VGND VGND VPWR VPWR _5779_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7518_ _6964_/Y _7513_/X _6884_/Y _7514_/X _7517_/X VGND VGND VPWR VPWR _7531_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8498_ _7903_/X _8358_/A _8138_/B _8178_/B VGND VGND VPWR VPWR _8776_/C sky130_fd_sc_hd__o22ai_1
X_7449_ _7477_/A _7479_/C _7471_/C VGND VGND VPWR VPWR _7498_/A sky130_fd_sc_hd__or3_2
XFILLER_174_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9119_ _9516_/CLK _9119_/D _9571_/SET_B VGND VGND VPWR VPWR _9119_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6820_ _9769_/Q VGND VGND VPWR VPWR _6820_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6751_ _9460_/Q VGND VGND VPWR VPWR _6751_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_50_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9470_ _9514_/CLK _9470_/D _9571_/SET_B VGND VGND VPWR VPWR _9470_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_5702_ _9309_/Q _5700_/A _6065_/B1 _5700_/Y VGND VGND VPWR VPWR _9309_/D sky130_fd_sc_hd__a22o_1
X_6682_ _9770_/Q VGND VGND VPWR VPWR _6682_/Y sky130_fd_sc_hd__inv_2
X_8421_ _8243_/A _8421_/B _8421_/C _8421_/D VGND VGND VPWR VPWR _8627_/A sky130_fd_sc_hd__and4b_1
X_5633_ _9346_/Q _5630_/A hold217/X _5630_/Y VGND VGND VPWR VPWR _9346_/D sky130_fd_sc_hd__a22o_1
X_5564_ _9393_/Q _5561_/A hold577/A _5561_/Y VGND VGND VPWR VPWR _5564_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8352_ _8613_/B _8352_/B _8539_/A _8351_/X VGND VGND VPWR VPWR _8352_/X sky130_fd_sc_hd__or4b_1
XFILLER_117_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold101 hold101/A VGND VGND VPWR VPWR _9391_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7303_ _6141_/Y _7151_/X _6110_/Y _7152_/X VGND VGND VPWR VPWR _7303_/X sky130_fd_sc_hd__o22a_1
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4515_ _9826_/Q _4513_/A hold510/X _4513_/Y VGND VGND VPWR VPWR _9826_/D sky130_fd_sc_hd__a22o_1
Xhold134 _8883_/X VGND VGND VPWR VPWR hold135/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 hold594/X VGND VGND VPWR VPWR hold593/A sky130_fd_sc_hd__buf_12
Xhold112 hold112/A VGND VGND VPWR VPWR hold113/A sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ _5495_/A VGND VGND VPWR VPWR _5495_/Y sky130_fd_sc_hd__inv_2
X_8283_ _8283_/A _8616_/B _8403_/B _8772_/B VGND VGND VPWR VPWR _8287_/A sky130_fd_sc_hd__or4_1
Xhold145 hold145/A VGND VGND VPWR VPWR _9408_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold156 hold156/A VGND VGND VPWR VPWR hold157/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _5348_/X VGND VGND VPWR VPWR hold168/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7234_ _6458_/Y _7135_/X _6421_/Y _7136_/X _7233_/X VGND VGND VPWR VPWR _7253_/A
+ sky130_fd_sc_hd__o221a_1
Xhold189 hold189/A VGND VGND VPWR VPWR hold190/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 hold602/X VGND VGND VPWR VPWR hold601/A sky130_fd_sc_hd__buf_12
X_7165_ _7165_/A _7165_/B _7165_/C _7165_/D VGND VGND VPWR VPWR _7187_/B sky130_fd_sc_hd__and4_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6116_/A VGND VGND VPWR VPWR _6116_/Y sky130_fd_sc_hd__inv_2
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7096_/A VGND VGND VPWR VPWR _9001_/S sky130_fd_sc_hd__buf_6
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6047_ _6047_/A VGND VGND VPWR VPWR _6047_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9806_ _9812_/CLK _9806_/D _7042_/B VGND VGND VPWR VPWR _9806_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7998_ _8230_/A _8140_/B VGND VGND VPWR VPWR _8006_/B sky130_fd_sc_hd__or2_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9737_ _9830_/CLK _9737_/D _9537_/SET_B VGND VGND VPWR VPWR _9737_/Q sky130_fd_sc_hd__dfrtp_1
X_6949_ _6944_/Y _4865_/X _6945_/Y _5647_/B _6948_/X VGND VGND VPWR VPWR _6956_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_14_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9668_ _9751_/CLK _9668_/D _5153_/X VGND VGND VPWR VPWR _9668_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8619_ _8619_/A _8619_/B _8619_/C VGND VGND VPWR VPWR _8717_/C sky130_fd_sc_hd__or3_1
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9599_ _9600_/CLK _9599_/D _9821_/SET_B VGND VGND VPWR VPWR _9599_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold690 _4488_/X VGND VGND VPWR VPWR hold690/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput217 _8812_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput206 _8850_/Y VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_2
Xoutput228 _8832_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_141_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5280_ _9584_/Q _5276_/A _8969_/A1 _5276_/Y VGND VGND VPWR VPWR _9584_/D sky130_fd_sc_hd__a22o_1
Xoutput239 _7736_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_4_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8970_ _9646_/Q hold136/X _8975_/S VGND VGND VPWR VPWR _8970_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7921_ _8436_/D _8053_/A VGND VGND VPWR VPWR _8439_/A sky130_fd_sc_hd__or2_4
XFILLER_82_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7852_ _8053_/A VGND VGND VPWR VPWR _8138_/B sky130_fd_sc_hd__buf_6
XFILLER_63_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7783_ _9110_/Q _7783_/A2 _9109_/Q _7783_/B2 _7782_/X VGND VGND VPWR VPWR _7783_/X
+ sky130_fd_sc_hd__a221o_1
X_4995_ _4995_/A VGND VGND VPWR VPWR _4995_/X sky130_fd_sc_hd__clkbuf_1
X_6803_ _9158_/Q VGND VGND VPWR VPWR _6803_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_189_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9522_ _9522_/CLK _9522_/D _9563_/SET_B VGND VGND VPWR VPWR _9522_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6734_ _6729_/Y _6282_/A _6730_/Y _4598_/B _6733_/X VGND VGND VPWR VPWR _6747_/B
+ sky130_fd_sc_hd__o221a_2
X_9453_ _9579_/CLK _9453_/D _9727_/SET_B VGND VGND VPWR VPWR _9453_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6665_ _9308_/Q VGND VGND VPWR VPWR _6665_/Y sky130_fd_sc_hd__inv_2
X_8404_ _8404_/A _8404_/B VGND VGND VPWR VPWR _8617_/C sky130_fd_sc_hd__or2_1
X_5616_ _9357_/Q _5611_/A hold42/X _5611_/Y VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__a22o_1
X_9384_ _9522_/CLK _9384_/D _9537_/SET_B VGND VGND VPWR VPWR _9384_/Q sky130_fd_sc_hd__dfrtp_1
X_6596_ _8825_/A _6058_/B _6595_/Y _4883_/X VGND VGND VPWR VPWR _6596_/X sky130_fd_sc_hd__o22a_1
X_8335_ _8419_/C _8246_/A _9109_/Q VGND VGND VPWR VPWR _8692_/C sky130_fd_sc_hd__o21ai_2
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5547_ _9404_/Q _5545_/A _6065_/B1 _5545_/Y VGND VGND VPWR VPWR _9404_/D sky130_fd_sc_hd__a22o_1
X_8266_ _8637_/C _8266_/B _8266_/C _8265_/X VGND VGND VPWR VPWR _8269_/B sky130_fd_sc_hd__or4b_2
X_5478_ _9451_/Q _5475_/X _6065_/B1 _5476_/Y VGND VGND VPWR VPWR _5478_/X sky130_fd_sc_hd__a22o_1
X_7217_ _8837_/A _7095_/B _8801_/A _7157_/X VGND VGND VPWR VPWR _7217_/X sky130_fd_sc_hd__o22a_1
X_8197_ _8197_/A _8620_/A VGND VGND VPWR VPWR _8199_/A sky130_fd_sc_hd__or2_1
X_7148_ _6964_/Y _7144_/X _6952_/Y _7145_/X _7147_/X VGND VGND VPWR VPWR _7165_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7079_ _7092_/A _7099_/B VGND VGND VPWR VPWR _7155_/A sky130_fd_sc_hd__or2_4
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4780_ _9336_/Q VGND VGND VPWR VPWR _7125_/A sky130_fd_sc_hd__clkinv_4
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_0_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9579_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6450_ _6448_/Y _5436_/B _6449_/Y _5047_/B VGND VGND VPWR VPWR _6450_/X sky130_fd_sc_hd__o22a_1
XFILLER_118_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6381_ _6379_/Y _5428_/B _6380_/Y _5301_/B VGND VGND VPWR VPWR _6381_/X sky130_fd_sc_hd__o22a_1
X_5401_ _9503_/Q _5399_/A _6065_/B1 _5399_/Y VGND VGND VPWR VPWR _9503_/D sky130_fd_sc_hd__a22o_1
XFILLER_173_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8120_ _8421_/D _8436_/B _8120_/C VGND VGND VPWR VPWR _8153_/A sky130_fd_sc_hd__or3_2
X_5332_ _9551_/Q _5331_/A hold516/X _5331_/Y VGND VGND VPWR VPWR _5332_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8051_ _8625_/A _8580_/B _8567_/C VGND VGND VPWR VPWR _8565_/A sky130_fd_sc_hd__or3_2
XFILLER_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5263_ _5378_/A _5263_/B VGND VGND VPWR VPWR _5264_/A sky130_fd_sc_hd__or2_1
X_5194_ _9642_/Q _5192_/A hold510/X _5192_/Y VGND VGND VPWR VPWR _5194_/X sky130_fd_sc_hd__a22o_1
XFILLER_141_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7002_ _6977_/Y _6995_/A _9063_/Q _6995_/Y VGND VGND VPWR VPWR _9063_/D sky130_fd_sc_hd__o22a_1
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8953_ _7758_/Y _4971_/A _9090_/Q VGND VGND VPWR VPWR _8953_/X sky130_fd_sc_hd__mux2_1
X_8884_ hold39/X hold611/X _8987_/S VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__mux2_8
X_7904_ _7999_/A _8570_/A _8567_/A _7904_/D VGND VGND VPWR VPWR _7905_/A sky130_fd_sc_hd__or4_4
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7835_ _8436_/C VGND VGND VPWR VPWR _8421_/C sky130_fd_sc_hd__inv_6
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7766_ _7766_/A _7766_/B _9110_/Q VGND VGND VPWR VPWR _7766_/X sky130_fd_sc_hd__and3_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9505_ _9561_/CLK _9505_/D _9817_/SET_B VGND VGND VPWR VPWR _9505_/Q sky130_fd_sc_hd__dfrtp_1
X_4978_ _6081_/A VGND VGND VPWR VPWR _5017_/A sky130_fd_sc_hd__buf_8
X_6717_ _9408_/Q VGND VGND VPWR VPWR _6717_/Y sky130_fd_sc_hd__inv_2
X_7697_ _6564_/Y _7493_/A _6640_/Y _7494_/A VGND VGND VPWR VPWR _7697_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9436_ _9522_/CLK _9436_/D _9563_/SET_B VGND VGND VPWR VPWR _9436_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6648_ _9672_/Q VGND VGND VPWR VPWR _6648_/Y sky130_fd_sc_hd__inv_2
X_9367_ _9421_/CLK _9367_/D _9537_/SET_B VGND VGND VPWR VPWR _9367_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8318_ _8702_/A _8702_/B _8538_/A VGND VGND VPWR VPWR _8322_/B sky130_fd_sc_hd__or3_1
XFILLER_105_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6579_ _6574_/Y _5397_/B _6575_/Y _5133_/B _6578_/X VGND VGND VPWR VPWR _6598_/A
+ sky130_fd_sc_hd__o221a_1
X_9298_ _9694_/CLK _9298_/D _9689_/SET_B VGND VGND VPWR VPWR _9298_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_117_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8249_ _8249_/A VGND VGND VPWR VPWR _8306_/B sky130_fd_sc_hd__buf_4
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5950_ _9165_/Q _5948_/A _8964_/A1 _5948_/Y VGND VGND VPWR VPWR _9165_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4901_ _9813_/Q VGND VGND VPWR VPWR _4901_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7620_ _6243_/Y _7525_/X _7292_/A _7526_/X _7619_/X VGND VGND VPWR VPWR _7621_/D
+ sky130_fd_sc_hd__o221a_1
X_5881_ _5878_/X _8910_/X _8960_/X _9216_/Q VGND VGND VPWR VPWR _9216_/D sky130_fd_sc_hd__o22a_1
X_4832_ _4832_/A _4953_/B VGND VGND VPWR VPWR _5274_/B sky130_fd_sc_hd__or2_4
XFILLER_60_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_190 _4826_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4763_ _9362_/Q VGND VGND VPWR VPWR _4763_/Y sky130_fd_sc_hd__clkinv_4
X_7551_ _8809_/A _7485_/A _8799_/A _7486_/A VGND VGND VPWR VPWR _7551_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4694_ _4681_/Y _5581_/B _4684_/Y _5935_/B _4693_/X VGND VGND VPWR VPWR _4725_/A
+ sky130_fd_sc_hd__o221a_1
X_6502_ _6500_/Y _4545_/B _6501_/Y _4892_/X VGND VGND VPWR VPWR _6502_/X sky130_fd_sc_hd__o22a_4
X_7482_ _7482_/A _7482_/B _7482_/C _7482_/D VGND VGND VPWR VPWR _7483_/D sky130_fd_sc_hd__and4_1
XFILLER_174_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9221_ _9225_/CLK _9221_/D _9537_/SET_B VGND VGND VPWR VPWR _9221_/Q sky130_fd_sc_hd__dfrtp_1
X_6433_ _9592_/Q VGND VGND VPWR VPWR _6433_/Y sky130_fd_sc_hd__inv_4
XFILLER_134_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9152_ _9734_/CLK _9152_/D _9731_/SET_B VGND VGND VPWR VPWR _9152_/Q sky130_fd_sc_hd__dfrtp_1
X_6364_ _6359_/Y _5482_/B _6360_/Y _5329_/B _6363_/X VGND VGND VPWR VPWR _6383_/A
+ sky130_fd_sc_hd__o221a_1
X_9083_ _9705_/CLK _9083_/D VGND VGND VPWR VPWR _9083_/Q sky130_fd_sc_hd__dfxtp_1
X_6295_ _9463_/Q VGND VGND VPWR VPWR _6295_/Y sky130_fd_sc_hd__inv_6
X_8103_ _8103_/A _8103_/B VGND VGND VPWR VPWR _8106_/A sky130_fd_sc_hd__or2_1
X_5315_ _5315_/A VGND VGND VPWR VPWR _5315_/Y sky130_fd_sc_hd__inv_2
X_5246_ _9606_/Q _5241_/Y hold613/X _5241_/A VGND VGND VPWR VPWR _5246_/X sky130_fd_sc_hd__o22a_1
X_8034_ _8034_/A _8034_/B VGND VGND VPWR VPWR _8157_/B sky130_fd_sc_hd__nand2_4
XFILLER_142_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold27 hold27/A VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_5177_ _9653_/Q _5170_/A _8969_/A1 _5170_/Y VGND VGND VPWR VPWR _9653_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8936_ _8935_/X _9190_/Q _9096_/Q VGND VGND VPWR VPWR _8936_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8867_ _9621_/Q _9760_/Q _9019_/S VGND VGND VPWR VPWR _8867_/X sky130_fd_sc_hd__mux2_1
X_7818_ _8009_/A _7812_/Y _7869_/A _7812_/A _8260_/A VGND VGND VPWR VPWR _7937_/B
+ sky130_fd_sc_hd__a221o_1
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8798_ _8798_/A VGND VGND VPWR VPWR _8798_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7749_ _9128_/Q _7748_/B _7750_/A VGND VGND VPWR VPWR _7749_/X sky130_fd_sc_hd__o21a_1
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9419_ _9420_/CLK _9419_/D _9537_/SET_B VGND VGND VPWR VPWR _9419_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold508 _9707_/Q VGND VGND VPWR VPWR hold509/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 _5650_/X VGND VGND VPWR VPWR _9335_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5100_ _5100_/A VGND VGND VPWR VPWR _9702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6080_ _6080_/A VGND VGND VPWR VPWR _6080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A VGND VGND VPWR VPWR _9739_/D sky130_fd_sc_hd__clkbuf_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9770_ _9817_/CLK _9770_/D _9821_/SET_B VGND VGND VPWR VPWR _9770_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6982_ _6982_/A VGND VGND VPWR VPWR _6983_/A sky130_fd_sc_hd__clkbuf_4
X_8721_ _8763_/A _8762_/C _8763_/C _8765_/C VGND VGND VPWR VPWR _8722_/C sky130_fd_sc_hd__or4_2
Xclkbuf_leaf_33_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9730_/CLK sky130_fd_sc_hd__clkbuf_16
X_5933_ _9176_/Q _5929_/A _8969_/A1 _5929_/Y VGND VGND VPWR VPWR _9176_/D sky130_fd_sc_hd__a22o_1
X_8652_ _7904_/D _7924_/X _7920_/A VGND VGND VPWR VPWR _8652_/Y sky130_fd_sc_hd__o21ai_1
X_5864_ _9228_/Q _5860_/A _8969_/A1 _5860_/Y VGND VGND VPWR VPWR _9228_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7603_ _7603_/A _7603_/B _7603_/C _7603_/D VGND VGND VPWR VPWR _7604_/D sky130_fd_sc_hd__and4_1
X_8583_ _8583_/A _8659_/B _8747_/D _8661_/D VGND VGND VPWR VPWR _8583_/Y sky130_fd_sc_hd__nor4_1
X_4815_ _4913_/B VGND VGND VPWR VPWR _4933_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_193_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5795_ _9274_/Q _5788_/A _8969_/A1 _5788_/Y VGND VGND VPWR VPWR _9274_/D sky130_fd_sc_hd__a22o_1
X_7534_ _6755_/Y _7485_/X _6695_/Y _7486_/X _7533_/X VGND VGND VPWR VPWR _7550_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4746_ _4737_/Y _5866_/B _4739_/Y _5620_/B _4745_/X VGND VGND VPWR VPWR _4812_/B
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_48_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9812_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4677_ _4969_/A VGND VGND VPWR VPWR _4678_/A sky130_fd_sc_hd__clkbuf_1
X_7465_ _7473_/A _7476_/B _7471_/C VGND VGND VPWR VPWR _7514_/A sky130_fd_sc_hd__or3_2
X_9204_ _9326_/CLK _9204_/D _9571_/SET_B VGND VGND VPWR VPWR _9204_/Q sky130_fd_sc_hd__dfrtp_1
X_6416_ _6416_/A VGND VGND VPWR VPWR _6416_/Y sky130_fd_sc_hd__inv_2
X_7396_ _6529_/Y _7160_/A _6582_/Y _7064_/A _7395_/X VGND VGND VPWR VPWR _7397_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6347_ _9316_/Q VGND VGND VPWR VPWR _6347_/Y sky130_fd_sc_hd__inv_2
X_9135_ _9574_/CLK _9135_/D _9571_/SET_B VGND VGND VPWR VPWR _9135_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9066_ _9723_/CLK _9066_/D VGND VGND VPWR VPWR _9066_/Q sky130_fd_sc_hd__dfxtp_1
X_6278_ _6276_/Y _4844_/X _6277_/Y _5417_/B VGND VGND VPWR VPWR _6278_/X sky130_fd_sc_hd__o22a_1
Xinput117 sram_ro_data[31] VGND VGND VPWR VPWR _6128_/A sky130_fd_sc_hd__clkbuf_1
Xinput106 sram_ro_data[21] VGND VGND VPWR VPWR _6283_/A sky130_fd_sc_hd__clkbuf_1
Xinput128 usr1_vcc_pwrgood VGND VGND VPWR VPWR _6624_/A sky130_fd_sc_hd__clkbuf_1
Xinput139 wb_adr_i[16] VGND VGND VPWR VPWR _7803_/B sky130_fd_sc_hd__clkbuf_1
X_8017_ _8132_/B _8028_/A VGND VGND VPWR VPWR _8137_/A sky130_fd_sc_hd__nand2_4
X_5229_ _9617_/Q _5226_/Y _8890_/X _5226_/A VGND VGND VPWR VPWR _9617_/D sky130_fd_sc_hd__o22a_1
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8919_ _7231_/Y _9677_/Q _9001_/S VGND VGND VPWR VPWR _8919_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_90 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_140_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4600_ _4600_/A VGND VGND VPWR VPWR _4600_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_175_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5580_ _9380_/Q _5572_/A hold601/A _5572_/Y VGND VGND VPWR VPWR _5580_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4531_ _9816_/Q _4527_/A _6067_/B1 _4527_/Y VGND VGND VPWR VPWR _9816_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold316 hold316/A VGND VGND VPWR VPWR hold317/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold305 hold305/A VGND VGND VPWR VPWR _9471_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7250_ _6461_/Y _7182_/X _6434_/Y _7183_/X VGND VGND VPWR VPWR _7250_/X sky130_fd_sc_hd__o22a_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6201_ _9334_/Q VGND VGND VPWR VPWR _6201_/Y sky130_fd_sc_hd__clkinv_2
Xhold338 hold338/A VGND VGND VPWR VPWR _9224_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold327 _5383_/X VGND VGND VPWR VPWR hold328/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold349 hold349/A VGND VGND VPWR VPWR hold350/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7181_ _7181_/A VGND VGND VPWR VPWR _7181_/X sky130_fd_sc_hd__buf_6
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _6130_/Y _4915_/X _6131_/Y _4863_/X VGND VGND VPWR VPWR _6132_/X sky130_fd_sc_hd__o22a_1
X_6063_ _9117_/Q _6059_/X hold577/A _6060_/Y VGND VGND VPWR VPWR _6063_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5014_/A _8999_/X VGND VGND VPWR VPWR _5024_/S sky130_fd_sc_hd__or2b_1
X_9822_ _9827_/CLK _9822_/D _9821_/SET_B VGND VGND VPWR VPWR _9822_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _9324_/Q VGND VGND VPWR VPWR _7358_/A sky130_fd_sc_hd__inv_2
X_9753_ net399_3/A _9753_/D _4678_/X VGND VGND VPWR VPWR _9753_/Q sky130_fd_sc_hd__dfrtn_1
X_8704_ _8704_/A _8704_/B _8704_/C _8703_/X VGND VGND VPWR VPWR _8705_/C sky130_fd_sc_hd__or4b_1
X_9684_ _9819_/CLK _9684_/D _9817_/SET_B VGND VGND VPWR VPWR _9684_/Q sky130_fd_sc_hd__dfrtp_1
X_5916_ _5889_/X _8932_/X _8960_/X _9189_/Q VGND VGND VPWR VPWR _9189_/D sky130_fd_sc_hd__o22a_1
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6896_ _9519_/Q VGND VGND VPWR VPWR _6896_/Y sky130_fd_sc_hd__inv_4
X_8635_ _7873_/B _8633_/Y _8683_/A _8543_/C VGND VGND VPWR VPWR _8737_/D sky130_fd_sc_hd__a211o_1
XFILLER_166_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5847_ _5847_/A _5847_/B VGND VGND VPWR VPWR _5848_/A sky130_fd_sc_hd__or2_1
XFILLER_139_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8566_ _8565_/Y _8559_/Y _8560_/X _8486_/A VGND VGND VPWR VPWR _8569_/C sky130_fd_sc_hd__a31o_1
X_5778_ _9282_/Q _5773_/A _6008_/B1 _5773_/Y VGND VGND VPWR VPWR _9282_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7517_ _6824_/Y _7515_/X _6939_/Y _7516_/X VGND VGND VPWR VPWR _7517_/X sky130_fd_sc_hd__o22a_1
X_8497_ _8497_/A _8497_/B VGND VGND VPWR VPWR _8501_/A sky130_fd_sc_hd__or2_1
X_4729_ _4764_/B VGND VGND VPWR VPWR _4801_/B sky130_fd_sc_hd__buf_2
XFILLER_135_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7448_ _7471_/A _7476_/B _9297_/Q VGND VGND VPWR VPWR _7497_/A sky130_fd_sc_hd__or3_2
XFILLER_174_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7379_ _6762_/Y _7171_/X _6749_/Y _7172_/X _7378_/X VGND VGND VPWR VPWR _7384_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9118_ _9514_/CLK _9118_/D _9571_/SET_B VGND VGND VPWR VPWR _9118_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9049_ _9642_/Q _8833_/A VGND VGND VPWR VPWR _9049_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_130_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6750_ _9450_/Q VGND VGND VPWR VPWR _6750_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5701_ _9310_/Q _5700_/A _6064_/B1 _5700_/Y VGND VGND VPWR VPWR _9310_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6681_ _9114_/Q VGND VGND VPWR VPWR _6681_/Y sky130_fd_sc_hd__clkinv_2
X_8420_ _8607_/A _8420_/B VGND VGND VPWR VPWR _8762_/C sky130_fd_sc_hd__nor2_1
X_5632_ _9347_/Q _5630_/A _6065_/B1 _5630_/Y VGND VGND VPWR VPWR _9347_/D sky130_fd_sc_hd__a22o_1
X_5563_ _9394_/Q _5561_/A hold510/X _5561_/Y VGND VGND VPWR VPWR _5563_/X sky130_fd_sc_hd__a22o_1
X_8351_ _7903_/X _8540_/A _8383_/B _8540_/B VGND VGND VPWR VPWR _8351_/X sky130_fd_sc_hd__o22a_1
XFILLER_129_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7302_ _6171_/Y _7144_/X _6151_/Y _7145_/X _7301_/X VGND VGND VPWR VPWR _7309_/A
+ sky130_fd_sc_hd__o221a_1
X_4514_ _9827_/Q _4513_/A hold516/X _4513_/Y VGND VGND VPWR VPWR _9827_/D sky130_fd_sc_hd__a22o_1
Xhold124 _5310_/X VGND VGND VPWR VPWR hold125/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 hold135/A VGND VGND VPWR VPWR hold136/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold113/A VGND VGND VPWR VPWR _9236_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold102 _5461_/X VGND VGND VPWR VPWR hold103/A sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ _5494_/A VGND VGND VPWR VPWR _5495_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_132_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8282_ _8358_/A _8306_/B VGND VGND VPWR VPWR _8772_/B sky130_fd_sc_hd__nor2_1
Xhold157 hold157/A VGND VGND VPWR VPWR _9646_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold146 _5644_/X VGND VGND VPWR VPWR hold147/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/A VGND VGND VPWR VPWR hold169/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7233_ _6402_/Y _7137_/X _6492_/Y _7138_/X _7232_/X VGND VGND VPWR VPWR _7233_/X
+ sky130_fd_sc_hd__o221a_1
X_7164_ _6910_/Y _7160_/X _6939_/Y _7071_/B _7163_/X VGND VGND VPWR VPWR _7165_/D
+ sky130_fd_sc_hd__o221a_1
Xhold179 _6068_/X VGND VGND VPWR VPWR hold180/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_86_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _9781_/Q VGND VGND VPWR VPWR _6115_/Y sky130_fd_sc_hd__inv_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7127_/A _7095_/B _7095_/C _7095_/D VGND VGND VPWR VPWR _7096_/A sky130_fd_sc_hd__and4_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6071_/A VGND VGND VPWR VPWR _6047_/A sky130_fd_sc_hd__clkbuf_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9805_ _9810_/CLK _9805_/D _9817_/SET_B VGND VGND VPWR VPWR _9805_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7997_ _8005_/A _8230_/A _8140_/B VGND VGND VPWR VPWR _8236_/B sky130_fd_sc_hd__or3_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9736_ _9736_/CLK _9736_/D _9731_/SET_B VGND VGND VPWR VPWR _9736_/Q sky130_fd_sc_hd__dfrtp_1
X_6948_ _6946_/Y _5532_/B _6947_/Y _5570_/B VGND VGND VPWR VPWR _6948_/X sky130_fd_sc_hd__o22a_1
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9667_ _9734_/CLK _9667_/D _9731_/SET_B VGND VGND VPWR VPWR _9667_/Q sky130_fd_sc_hd__dfrtp_1
X_6879_ _9553_/Q VGND VGND VPWR VPWR _6879_/Y sky130_fd_sc_hd__clkinv_2
X_8618_ _8618_/A _8684_/D _8772_/D _8618_/D VGND VGND VPWR VPWR _8622_/A sky130_fd_sc_hd__or4_1
XFILLER_10_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9598_ _9600_/CLK _9598_/D _9821_/SET_B VGND VGND VPWR VPWR _9598_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8549_ _7918_/A _7920_/A _7887_/A _8342_/B _7970_/A VGND VGND VPWR VPWR _8642_/B
+ sky130_fd_sc_hd__o221ai_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold680 _5475_/X VGND VGND VPWR VPWR _5476_/A sky130_fd_sc_hd__clkbuf_2
Xhold691 _8985_/X VGND VGND VPWR VPWR hold691/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput207 _8873_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_181_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput218 _8874_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_2
Xoutput229 _8786_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_181_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7920_ _7920_/A VGND VGND VPWR VPWR _8608_/A sky130_fd_sc_hd__inv_2
X_7851_ _7851_/A VGND VGND VPWR VPWR _8053_/A sky130_fd_sc_hd__buf_6
XFILLER_82_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6802_ _6797_/Y _4929_/X _6798_/Y _5482_/B _6801_/X VGND VGND VPWR VPWR _6814_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7782_ _9108_/Q _7782_/B VGND VGND VPWR VPWR _7782_/X sky130_fd_sc_hd__and2_1
X_4994_ _5017_/A VGND VGND VPWR VPWR _4995_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_90_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9521_ _9569_/CLK hold59/X _9563_/SET_B VGND VGND VPWR VPWR _9521_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6733_ _6731_/Y _5505_/B _6732_/Y _5589_/B VGND VGND VPWR VPWR _6733_/X sky130_fd_sc_hd__o22a_1
XFILLER_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6664_ _9313_/Q VGND VGND VPWR VPWR _6664_/Y sky130_fd_sc_hd__inv_2
X_9452_ _9579_/CLK _9452_/D _7042_/B VGND VGND VPWR VPWR _9452_/Q sky130_fd_sc_hd__dfrtp_1
X_5615_ _9358_/Q _5611_/A hold53/X _5611_/Y VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__a22o_1
X_8403_ _8403_/A _8403_/B VGND VGND VPWR VPWR _8772_/C sky130_fd_sc_hd__or2_1
XFILLER_176_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9383_ _9522_/CLK _9383_/D _9563_/SET_B VGND VGND VPWR VPWR _9383_/Q sky130_fd_sc_hd__dfrtp_1
X_6595_ _6595_/A VGND VGND VPWR VPWR _6595_/Y sky130_fd_sc_hd__inv_2
X_8334_ _8556_/A _8334_/B VGND VGND VPWR VPWR _8336_/A sky130_fd_sc_hd__nor2_1
XFILLER_117_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5546_ _9405_/Q _5545_/A _6064_/B1 _5545_/Y VGND VGND VPWR VPWR _9405_/D sky130_fd_sc_hd__a22o_1
XFILLER_155_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8265_ _8265_/A _8265_/B VGND VGND VPWR VPWR _8265_/X sky130_fd_sc_hd__and2_1
X_5477_ _9452_/Q _5476_/A _6064_/B1 _5476_/Y VGND VGND VPWR VPWR _9452_/D sky130_fd_sc_hd__a22o_1
X_7216_ _8817_/A _7149_/X _8797_/A _7150_/X _7215_/X VGND VGND VPWR VPWR _7221_/B
+ sky130_fd_sc_hd__o221a_1
X_8196_ _8243_/B _8594_/A VGND VGND VPWR VPWR _8620_/A sky130_fd_sc_hd__nor2_1
XFILLER_59_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7147_ _6941_/Y _7071_/C _6830_/Y _7146_/X VGND VGND VPWR VPWR _7147_/X sky130_fd_sc_hd__o22a_1
XFILLER_100_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7078_ _9290_/Q _7081_/B _7129_/A VGND VGND VPWR VPWR _7099_/B sky130_fd_sc_hd__or3_1
XFILLER_104_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6029_ _6029_/A VGND VGND VPWR VPWR _6029_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9719_ _9723_/CLK _9719_/D _6177_/A VGND VGND VPWR VPWR _9719_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6380_ _9566_/Q VGND VGND VPWR VPWR _6380_/Y sky130_fd_sc_hd__inv_4
X_5400_ _9504_/Q _5399_/A _6064_/B1 _5399_/Y VGND VGND VPWR VPWR _9504_/D sky130_fd_sc_hd__a22o_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5331_ _5331_/A VGND VGND VPWR VPWR _5331_/Y sky130_fd_sc_hd__inv_2
X_8050_ _7903_/A _8126_/A _8049_/X VGND VGND VPWR VPWR _8056_/B sky130_fd_sc_hd__o21ai_1
X_7001_ _6816_/Y _6995_/A _9064_/Q _6995_/Y VGND VGND VPWR VPWR _9064_/D sky130_fd_sc_hd__o22a_1
X_5262_ _9596_/Q _5257_/A _8975_/A1 _5257_/Y VGND VGND VPWR VPWR _9596_/D sky130_fd_sc_hd__a22o_1
X_5193_ _9643_/Q _5192_/A hold516/X _5192_/Y VGND VGND VPWR VPWR _5193_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8952_ _7747_/Y _9126_/Q _9093_/Q VGND VGND VPWR VPWR _8952_/X sky130_fd_sc_hd__mux2_1
X_8883_ hold133/X hold251/X _8883_/S VGND VGND VPWR VPWR _8883_/X sky130_fd_sc_hd__mux2_8
X_7903_ _7903_/A VGND VGND VPWR VPWR _7903_/X sky130_fd_sc_hd__buf_6
X_7834_ _8552_/A _8229_/B VGND VGND VPWR VPWR _8693_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7765_ _7765_/A _7766_/A _9108_/Q VGND VGND VPWR VPWR _7765_/X sky130_fd_sc_hd__and3_1
X_6716_ _9727_/Q VGND VGND VPWR VPWR _6716_/Y sky130_fd_sc_hd__inv_2
X_9504_ _9729_/CLK _9504_/D _9727_/SET_B VGND VGND VPWR VPWR _9504_/Q sky130_fd_sc_hd__dfrtp_1
X_4977_ _4971_/Y _4973_/Y _4974_/Y _4976_/X VGND VGND VPWR VPWR _9751_/D sky130_fd_sc_hd__o22ai_1
XFILLER_137_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7696_ _6586_/Y _7485_/X _6528_/Y _7486_/X _7695_/X VGND VGND VPWR VPWR _7712_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9435_ _9522_/CLK _9435_/D _9563_/SET_B VGND VGND VPWR VPWR _9435_/Q sky130_fd_sc_hd__dfrtp_1
X_6647_ _9487_/Q VGND VGND VPWR VPWR _8835_/A sky130_fd_sc_hd__clkinv_8
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9366_ _9421_/CLK _9366_/D _9537_/SET_B VGND VGND VPWR VPWR _9366_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6578_ _6576_/Y _4634_/B _6577_/Y _4598_/B VGND VGND VPWR VPWR _6578_/X sky130_fd_sc_hd__o22a_2
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5529_ _9416_/Q _5523_/A _8965_/A1 _5523_/Y VGND VGND VPWR VPWR _9416_/D sky130_fd_sc_hd__a22o_1
X_8317_ _8317_/A _8735_/B VGND VGND VPWR VPWR _8317_/X sky130_fd_sc_hd__or2_2
X_9297_ _9297_/CLK _9297_/D _9730_/SET_B VGND VGND VPWR VPWR _9297_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_59_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8248_ _8314_/A _8268_/C VGND VGND VPWR VPWR _8249_/A sky130_fd_sc_hd__or2_1
XFILLER_78_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8179_ _8179_/A _8180_/A VGND VGND VPWR VPWR _8403_/A sky130_fd_sc_hd__nor2_1
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4900_ _4900_/A _4953_/B VGND VGND VPWR VPWR _5521_/B sky130_fd_sc_hd__or2_4
XFILLER_73_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5880_ _5878_/X _8912_/X _8960_/X _9217_/Q VGND VGND VPWR VPWR _9217_/D sky130_fd_sc_hd__o22a_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4831_ _9583_/Q VGND VGND VPWR VPWR _4831_/Y sky130_fd_sc_hd__inv_4
XANTENNA_191 _6383_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_180 _9811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7550_ _7550_/A _7550_/B _7550_/C _7550_/D VGND VGND VPWR VPWR _7550_/Y sky130_fd_sc_hd__nand4_4
X_4762_ _4827_/A _4801_/B VGND VGND VPWR VPWR _5847_/B sky130_fd_sc_hd__or2_4
XFILLER_159_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4693_ _4688_/Y _5902_/B _4691_/Y _5551_/B VGND VGND VPWR VPWR _4693_/X sky130_fd_sc_hd__o22a_1
X_7481_ _4688_/Y _7525_/A _7125_/A _7526_/A _7480_/X VGND VGND VPWR VPWR _7482_/D
+ sky130_fd_sc_hd__o221a_1
X_6501_ _6501_/A VGND VGND VPWR VPWR _6501_/Y sky130_fd_sc_hd__inv_2
X_9220_ _9830_/CLK _9220_/D _9537_/SET_B VGND VGND VPWR VPWR _9220_/Q sky130_fd_sc_hd__dfstp_1
X_6432_ _6427_/Y _5367_/B _6428_/Y _5321_/B _6431_/X VGND VGND VPWR VPWR _6439_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9151_ _9736_/CLK _9151_/D _9731_/SET_B VGND VGND VPWR VPWR _9151_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8102_ _8102_/A _8105_/B _8102_/C VGND VGND VPWR VPWR _8103_/B sky130_fd_sc_hd__and3_1
X_6363_ _6361_/Y _5313_/B _6362_/Y _5946_/B VGND VGND VPWR VPWR _6363_/X sky130_fd_sc_hd__o22a_2
X_9082_ _9705_/CLK _9082_/D VGND VGND VPWR VPWR _9082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6294_ _9593_/Q VGND VGND VPWR VPWR _6294_/Y sky130_fd_sc_hd__inv_6
X_5314_ _5314_/A VGND VGND VPWR VPWR _5315_/A sky130_fd_sc_hd__clkbuf_2
X_5245_ _9607_/Q _5241_/Y _8963_/X _5241_/A VGND VGND VPWR VPWR _5245_/X sky130_fd_sc_hd__o22a_1
X_8033_ _8175_/A VGND VGND VPWR VPWR _8178_/B sky130_fd_sc_hd__buf_2
XFILLER_102_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold17 hold17/A VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold28 hold28/A VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5176_ _9654_/Q _5170_/A _8965_/A1 _5170_/Y VGND VGND VPWR VPWR _9654_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8935_ _7407_/Y _9672_/Q _9001_/S VGND VGND VPWR VPWR _8935_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _9718_/CLK sky130_fd_sc_hd__clkbuf_2
X_8866_ _9620_/Q input3/X input1/X VGND VGND VPWR VPWR _8866_/X sky130_fd_sc_hd__mux2_2
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7817_ _7869_/A _7874_/B _7816_/Y _7874_/C _5964_/X VGND VGND VPWR VPWR _8260_/A
+ sky130_fd_sc_hd__a32o_2
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8797_ _8797_/A VGND VGND VPWR VPWR _8798_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7748_ _9128_/Q _7748_/B VGND VGND VPWR VPWR _7750_/A sky130_fd_sc_hd__nand2_1
XFILLER_177_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7679_ _6763_/Y _7493_/X _6793_/Y _7494_/X VGND VGND VPWR VPWR _7679_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9418_ _9418_/CLK _9418_/D _9731_/SET_B VGND VGND VPWR VPWR _9418_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9349_ _9678_/CLK _9349_/D _9730_/SET_B VGND VGND VPWR VPWR _9349_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput390 _9054_/Q VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold509 hold509/A VGND VGND VPWR VPWR hold509/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_171_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _4971_/A _9739_/Q _5030_/S VGND VGND VPWR VPWR _5031_/A sky130_fd_sc_hd__mux2_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6981_ _7005_/B _6981_/B VGND VGND VPWR VPWR _6982_/A sky130_fd_sc_hd__or2_1
XFILLER_65_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8720_ _8720_/A _8720_/B _8720_/C VGND VGND VPWR VPWR _8765_/C sky130_fd_sc_hd__or3_1
X_5932_ _9177_/Q _5929_/A _8965_/A1 _5929_/Y VGND VGND VPWR VPWR _9177_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8651_ _8651_/A VGND VGND VPWR VPWR _8708_/C sky130_fd_sc_hd__inv_2
X_5863_ _9229_/Q _5860_/A _8965_/A1 _5860_/Y VGND VGND VPWR VPWR _9229_/D sky130_fd_sc_hd__a22o_1
X_5794_ _9275_/Q _5788_/A _8965_/A1 _5788_/Y VGND VGND VPWR VPWR _9275_/D sky130_fd_sc_hd__a22o_1
X_7602_ _6333_/Y _7525_/X _7270_/A _7526_/X _7601_/X VGND VGND VPWR VPWR _7603_/D
+ sky130_fd_sc_hd__o221a_1
X_8582_ _8582_/A _8746_/B VGND VGND VPWR VPWR _8661_/D sky130_fd_sc_hd__or2_1
X_4814_ _9588_/Q VGND VGND VPWR VPWR _4814_/Y sky130_fd_sc_hd__clkinv_4
X_7533_ _6767_/Y _7487_/X _6704_/Y _7488_/X VGND VGND VPWR VPWR _7533_/X sky130_fd_sc_hd__o22a_1
X_4745_ _4741_/Y _5706_/B _4743_/Y _5797_/B VGND VGND VPWR VPWR _4745_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4676_ _9754_/Q _4657_/A _8994_/X _4657_/Y VGND VGND VPWR VPWR _9754_/D sky130_fd_sc_hd__a22o_1
X_7464_ _7478_/C _7473_/A _9297_/Q VGND VGND VPWR VPWR _7513_/A sky130_fd_sc_hd__or3_2
XFILLER_162_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9203_ _9326_/CLK _9203_/D _9571_/SET_B VGND VGND VPWR VPWR _9203_/Q sky130_fd_sc_hd__dfstp_1
X_6415_ _9794_/Q VGND VGND VPWR VPWR _6415_/Y sky130_fd_sc_hd__inv_2
X_7395_ _6612_/Y _7161_/A _6628_/Y _7162_/A VGND VGND VPWR VPWR _7395_/X sky130_fd_sc_hd__o22a_1
XFILLER_162_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6346_ _9153_/Q VGND VGND VPWR VPWR _6346_/Y sky130_fd_sc_hd__clkinv_2
X_9134_ _8879_/A1 _9134_/D _6010_/X VGND VGND VPWR VPWR _9134_/Q sky130_fd_sc_hd__dfrtp_4
X_9065_ _9723_/CLK _9065_/D VGND VGND VPWR VPWR _9065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8016_ _8005_/A _8006_/B _8236_/B VGND VGND VPWR VPWR _8028_/A sky130_fd_sc_hd__a21bo_1
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6277_ _9489_/Q VGND VGND VPWR VPWR _6277_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput118 sram_ro_data[3] VGND VGND VPWR VPWR _6595_/A sky130_fd_sc_hd__clkbuf_1
Xinput107 sram_ro_data[22] VGND VGND VPWR VPWR _6250_/A sky130_fd_sc_hd__clkbuf_1
Xinput129 usr1_vdd_pwrgood VGND VGND VPWR VPWR _6878_/A sky130_fd_sc_hd__clkbuf_1
X_5228_ _9618_/Q _5226_/Y _8968_/X _5226_/A VGND VGND VPWR VPWR _5228_/X sky130_fd_sc_hd__o22a_1
X_5159_ _5159_/A VGND VGND VPWR VPWR _5159_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8918_ _8917_/X _9181_/Q _9096_/Q VGND VGND VPWR VPWR _8918_/X sky130_fd_sc_hd__mux2_1
X_8849_ _8849_/A _8849_/B VGND VGND VPWR VPWR _8849_/Y sky130_fd_sc_hd__nor2_2
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_80 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4530_ _9817_/Q _4527_/A hold217/X _4527_/Y VGND VGND VPWR VPWR _9817_/D sky130_fd_sc_hd__a22o_1
Xhold306 _5564_/X VGND VGND VPWR VPWR hold307/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold317 hold317/A VGND VGND VPWR VPWR _9575_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold339 _9801_/Q VGND VGND VPWR VPWR hold340/A sky130_fd_sc_hd__dlygate4sd3_1
X_6200_ _9550_/Q VGND VGND VPWR VPWR _6200_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold328 hold328/A VGND VGND VPWR VPWR hold329/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7180_ _7180_/A VGND VGND VPWR VPWR _7180_/X sky130_fd_sc_hd__buf_6
XFILLER_131_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _6131_/A VGND VGND VPWR VPWR _6131_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _9118_/Q _6060_/A hold510/A _6060_/Y VGND VGND VPWR VPWR _6062_/X sky130_fd_sc_hd__a22o_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5013_ _7039_/A _6023_/B _4989_/A _6053_/B _5012_/X VGND VGND VPWR VPWR _5014_/A
+ sky130_fd_sc_hd__o32a_1
X_9821_ _9827_/CLK _9821_/D _9821_/SET_B VGND VGND VPWR VPWR _9821_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_38_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6964_ _9233_/Q VGND VGND VPWR VPWR _6964_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9752_ net399_3/A _9752_/D _4961_/X VGND VGND VPWR VPWR _9752_/Q sky130_fd_sc_hd__dfrtn_1
X_8703_ _8702_/C _8383_/A _8702_/B _8702_/X _8598_/Y VGND VGND VPWR VPWR _8703_/X
+ sky130_fd_sc_hd__o311a_1
X_9683_ _9686_/CLK _9683_/D _9817_/SET_B VGND VGND VPWR VPWR _9683_/Q sky130_fd_sc_hd__dfrtp_1
X_5915_ _5889_/X _8934_/X _8960_/X _9190_/Q VGND VGND VPWR VPWR _9190_/D sky130_fd_sc_hd__o22a_1
X_6895_ _6890_/Y _5521_/B _6891_/Y _5263_/B _6894_/X VGND VGND VPWR VPWR _6908_/B
+ sky130_fd_sc_hd__o221a_1
X_8634_ _8634_/A VGND VGND VPWR VPWR _8683_/A sky130_fd_sc_hd__inv_2
X_5846_ _9240_/Q _5841_/A _6008_/B1 _5841_/Y VGND VGND VPWR VPWR _9240_/D sky130_fd_sc_hd__a22o_1
XFILLER_166_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8565_ _8565_/A VGND VGND VPWR VPWR _8565_/Y sky130_fd_sc_hd__inv_2
X_5777_ _9283_/Q _5773_/A _6067_/B1 _5773_/Y VGND VGND VPWR VPWR _9283_/D sky130_fd_sc_hd__a22o_1
X_4728_ _9260_/Q VGND VGND VPWR VPWR _4728_/Y sky130_fd_sc_hd__inv_2
X_8496_ _8496_/A _8496_/B VGND VGND VPWR VPWR _8497_/B sky130_fd_sc_hd__nand2_1
X_7516_ _7516_/A VGND VGND VPWR VPWR _7516_/X sky130_fd_sc_hd__buf_6
XFILLER_147_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4659_ _4969_/A VGND VGND VPWR VPWR _4660_/A sky130_fd_sc_hd__clkbuf_1
X_7447_ _4728_/Y _7491_/A _4721_/Y _7492_/A _7446_/X VGND VGND VPWR VPWR _7483_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7378_ _6810_/Y _7173_/X _6699_/Y _7174_/X VGND VGND VPWR VPWR _7378_/X sky130_fd_sc_hd__o22a_1
X_6329_ _9237_/Q VGND VGND VPWR VPWR _6329_/Y sky130_fd_sc_hd__clkinv_2
X_9117_ _9577_/CLK _9117_/D _9571_/SET_B VGND VGND VPWR VPWR _9117_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9048_ _9641_/Q _8831_/A VGND VGND VPWR VPWR _9048_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_76_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_32_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9678_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_47_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9810_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_180_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5700_ _5700_/A VGND VGND VPWR VPWR _5700_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6680_ _6680_/A _6680_/B _6680_/C VGND VGND VPWR VPWR _6816_/A sky130_fd_sc_hd__and3_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5631_ _9348_/Q _5630_/A _6064_/B1 _5630_/Y VGND VGND VPWR VPWR _9348_/D sky130_fd_sc_hd__a22o_1
X_5562_ _9395_/Q _5561_/A hold516/X _5561_/Y VGND VGND VPWR VPWR _5562_/X sky130_fd_sc_hd__a22o_1
X_8350_ _7873_/A _8341_/A _7873_/B _7918_/Y VGND VGND VPWR VPWR _8539_/A sky130_fd_sc_hd__a31o_1
XFILLER_129_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7301_ _6160_/Y _7071_/C _6154_/Y _7146_/X VGND VGND VPWR VPWR _7301_/X sky130_fd_sc_hd__o22a_1
X_8281_ _8288_/A _8281_/B VGND VGND VPWR VPWR _8403_/B sky130_fd_sc_hd__nor2_1
X_4513_ _4513_/A VGND VGND VPWR VPWR _4513_/Y sky130_fd_sc_hd__clkinv_2
Xhold125 hold125/A VGND VGND VPWR VPWR hold126/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 _5206_/X VGND VGND VPWR VPWR hold115/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 hold103/A VGND VGND VPWR VPWR hold104/A sky130_fd_sc_hd__dlygate4sd3_1
X_5493_ _5570_/A _6112_/B VGND VGND VPWR VPWR _5494_/A sky130_fd_sc_hd__or2_1
X_7232_ _6446_/Y _7139_/X _6388_/Y _7140_/X VGND VGND VPWR VPWR _7232_/X sky130_fd_sc_hd__o22a_1
Xhold158 _5207_/X VGND VGND VPWR VPWR hold159/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 hold136/A VGND VGND VPWR VPWR hold136/X sky130_fd_sc_hd__buf_12
Xhold147 hold147/A VGND VGND VPWR VPWR hold148/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 hold169/A VGND VGND VPWR VPWR _9538_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7163_ _6921_/Y _7161_/X _6891_/Y _7162_/X VGND VGND VPWR VPWR _7163_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6114_ _9595_/Q VGND VGND VPWR VPWR _6114_/Y sky130_fd_sc_hd__inv_6
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _7094_/A _7094_/B _7094_/C _7094_/D VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__and4_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _9125_/Q _6026_/A _8950_/X _6026_/Y VGND VGND VPWR VPWR _9125_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9804_ _9810_/CLK _9804_/D _7042_/B VGND VGND VPWR VPWR _9804_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7996_ _8421_/C _7996_/B _7996_/C VGND VGND VPWR VPWR _8140_/B sky130_fd_sc_hd__or3_1
X_9735_ _9830_/CLK _9735_/D _9537_/SET_B VGND VGND VPWR VPWR _9735_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6947_ _9381_/Q VGND VGND VPWR VPWR _6947_/Y sky130_fd_sc_hd__inv_2
X_6878_ _6878_/A VGND VGND VPWR VPWR _6878_/Y sky130_fd_sc_hd__inv_4
XFILLER_169_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9666_ _9734_/CLK _9666_/D _9731_/SET_B VGND VGND VPWR VPWR _9666_/Q sky130_fd_sc_hd__dfrtp_1
X_5829_ _9253_/Q _5828_/A hold516/X _5828_/Y VGND VGND VPWR VPWR _5829_/X sky130_fd_sc_hd__a22o_1
X_8617_ _8617_/A _8617_/B _8617_/C VGND VGND VPWR VPWR _8618_/D sky130_fd_sc_hd__or3_1
X_9597_ _9600_/CLK _9597_/D _9821_/SET_B VGND VGND VPWR VPWR _9597_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8548_ _8657_/A _8548_/B _8548_/C VGND VGND VPWR VPWR _8735_/A sky130_fd_sc_hd__or3_2
XFILLER_135_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8479_ _8674_/A _8479_/B VGND VGND VPWR VPWR _8746_/B sky130_fd_sc_hd__nor2_1
XFILLER_108_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold670 _5232_/X VGND VGND VPWR VPWR _9614_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold681 _5474_/X VGND VGND VPWR VPWR _5475_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold692 _8856_/X VGND VGND VPWR VPWR _9833_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_76_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput208 _8794_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_2
Xoutput219 _8814_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_153_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7850_ _8421_/C _7876_/A _8436_/A _8436_/B VGND VGND VPWR VPWR _7851_/A sky130_fd_sc_hd__or4_1
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6801_ _6799_/Y _4585_/B _6800_/Y _6117_/X VGND VGND VPWR VPWR _6801_/X sky130_fd_sc_hd__o22a_1
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7781_ _9110_/Q _7781_/A2 _9109_/Q _7781_/B2 _7780_/X VGND VGND VPWR VPWR _7781_/X
+ sky130_fd_sc_hd__a221o_1
X_4993_ _9748_/Q _4989_/A _9747_/Q _4989_/Y VGND VGND VPWR VPWR _9748_/D sky130_fd_sc_hd__a22o_1
XFILLER_90_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9520_ _9569_/CLK _9520_/D _9563_/SET_B VGND VGND VPWR VPWR _9520_/Q sky130_fd_sc_hd__dfrtp_1
X_6732_ _9372_/Q VGND VGND VPWR VPWR _6732_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6663_ _9351_/Q VGND VGND VPWR VPWR _6663_/Y sky130_fd_sc_hd__inv_2
X_9451_ _9579_/CLK _9451_/D _7042_/B VGND VGND VPWR VPWR _9451_/Q sky130_fd_sc_hd__dfrtp_1
X_5614_ _9359_/Q _5611_/A hold577/A _5611_/Y VGND VGND VPWR VPWR _5614_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8402_ _8402_/A _8615_/C _8684_/C _8616_/C VGND VGND VPWR VPWR _8406_/A sky130_fd_sc_hd__or4_1
XFILLER_164_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9382_ _9522_/CLK _9382_/D _9563_/SET_B VGND VGND VPWR VPWR _9382_/Q sky130_fd_sc_hd__dfrtp_1
X_6594_ _9115_/Q VGND VGND VPWR VPWR _8825_/A sky130_fd_sc_hd__clkinv_8
X_8333_ _8714_/C _8692_/B _8333_/C VGND VGND VPWR VPWR _8334_/B sky130_fd_sc_hd__or3_1
X_5545_ _5545_/A VGND VGND VPWR VPWR _5545_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8264_ _8288_/A _8540_/A _8264_/C VGND VGND VPWR VPWR _8265_/B sky130_fd_sc_hd__or3_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5476_ _5476_/A VGND VGND VPWR VPWR _5476_/Y sky130_fd_sc_hd__inv_2
X_7215_ _8819_/A _7151_/X _8829_/A _7152_/X VGND VGND VPWR VPWR _7215_/X sky130_fd_sc_hd__o22a_1
XFILLER_132_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8195_ _8195_/A _8409_/A VGND VGND VPWR VPWR _8197_/A sky130_fd_sc_hd__or2_1
X_7146_ _7146_/A VGND VGND VPWR VPWR _7146_/X sky130_fd_sc_hd__buf_4
XFILLER_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7077_ _7108_/C _7128_/A _7084_/C VGND VGND VPWR VPWR _7157_/A sky130_fd_sc_hd__or3_4
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6028_ _6071_/A VGND VGND VPWR VPWR _6029_/A sky130_fd_sc_hd__clkbuf_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7979_ _8243_/A _8383_/A _7978_/X VGND VGND VPWR VPWR _7980_/B sky130_fd_sc_hd__o21ai_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9718_ _9718_/CLK _9718_/D _6177_/A VGND VGND VPWR VPWR _9718_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9649_ _9651_/CLK _9649_/D _9689_/SET_B VGND VGND VPWR VPWR _9649_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5330_ _5330_/A VGND VGND VPWR VPWR _5331_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_141_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5261_ _9597_/Q _5257_/A _6067_/B1 _5257_/Y VGND VGND VPWR VPWR _9597_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7000_ _6660_/Y _6995_/A _9065_/Q _6995_/Y VGND VGND VPWR VPWR _9065_/D sky130_fd_sc_hd__o22a_1
X_5192_ _5192_/A VGND VGND VPWR VPWR _5192_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8951_ _7744_/X _9125_/Q _9093_/Q VGND VGND VPWR VPWR _8951_/X sky130_fd_sc_hd__mux2_1
X_7902_ _8268_/C _8347_/A VGND VGND VPWR VPWR _7903_/A sky130_fd_sc_hd__or2_1
XFILLER_83_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8882_ hold120/X hold592/X _9629_/Q VGND VGND VPWR VPWR _8882_/X sky130_fd_sc_hd__mux2_8
X_7833_ _7833_/A VGND VGND VPWR VPWR _8229_/B sky130_fd_sc_hd__buf_2
XFILLER_51_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7764_ _7764_/A VGND VGND VPWR VPWR _9002_/S sky130_fd_sc_hd__clkbuf_1
XFILLER_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6715_ _6710_/Y _4883_/X _6711_/Y _6353_/A _6714_/X VGND VGND VPWR VPWR _6721_/C
+ sky130_fd_sc_hd__o221a_1
X_4976_ _4975_/Y _7039_/A _9134_/Q _9090_/Q _9133_/Q VGND VGND VPWR VPWR _4976_/X
+ sky130_fd_sc_hd__o2111a_1
X_9503_ _9579_/CLK _9503_/D _9727_/SET_B VGND VGND VPWR VPWR _9503_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7695_ _6620_/Y _7487_/A _6560_/Y _7488_/A VGND VGND VPWR VPWR _7695_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9434_ _9522_/CLK _9434_/D _9563_/SET_B VGND VGND VPWR VPWR _9434_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6646_ _9529_/Q VGND VGND VPWR VPWR _6646_/Y sky130_fd_sc_hd__inv_2
X_9365_ _9643_/CLK _9365_/D _9563_/SET_B VGND VGND VPWR VPWR _9365_/Q sky130_fd_sc_hd__dfrtp_1
X_6577_ _9785_/Q VGND VGND VPWR VPWR _6577_/Y sky130_fd_sc_hd__inv_2
X_5528_ _9417_/Q _5523_/A _8964_/A1 _5523_/Y VGND VGND VPWR VPWR _9417_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8316_ _8552_/A _8702_/B _8538_/A VGND VGND VPWR VPWR _8735_/B sky130_fd_sc_hd__nor3_1
X_9296_ _9297_/CLK _9296_/D _9730_/SET_B VGND VGND VPWR VPWR _9296_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5459_ _9464_/Q _5456_/X hold510/X _5457_/Y VGND VGND VPWR VPWR _5459_/X sky130_fd_sc_hd__a22o_1
X_8247_ _8277_/A _8347_/B _8268_/C VGND VGND VPWR VPWR _8637_/B sky130_fd_sc_hd__nor3_1
XFILLER_105_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8178_ _8255_/A _8178_/B VGND VGND VPWR VPWR _8616_/A sky130_fd_sc_hd__nor2_1
XFILLER_59_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7129_ _7129_/A _7129_/B _7129_/C VGND VGND VPWR VPWR _7183_/A sky130_fd_sc_hd__or3_2
XFILLER_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_opt_2_0_wb_clk_i _9297_/CLK VGND VGND VPWR VPWR clkbuf_opt_2_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 _8827_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4830_ _4830_/A VGND VGND VPWR VPWR _4830_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_192 _6710_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_181 _8847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4761_ _9232_/Q VGND VGND VPWR VPWR _4761_/Y sky130_fd_sc_hd__inv_4
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4692_ _4866_/A _4808_/A VGND VGND VPWR VPWR _5551_/B sky130_fd_sc_hd__or2_4
X_7480_ _4836_/Y _7527_/A _4747_/Y _7528_/A VGND VGND VPWR VPWR _7480_/X sky130_fd_sc_hd__o22a_1
X_6500_ _9808_/Q VGND VGND VPWR VPWR _6500_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6431_ _6429_/Y _5559_/B _6430_/Y _5389_/B VGND VGND VPWR VPWR _6431_/X sky130_fd_sc_hd__o22a_1
XFILLER_146_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9150_ _9491_/CLK _9150_/D _9731_/SET_B VGND VGND VPWR VPWR _9150_/Q sky130_fd_sc_hd__dfrtp_1
X_6362_ _9166_/Q VGND VGND VPWR VPWR _6362_/Y sky130_fd_sc_hd__clkinv_2
X_8101_ _8101_/A VGND VGND VPWR VPWR _8102_/C sky130_fd_sc_hd__inv_2
X_5313_ _5474_/A _5313_/B VGND VGND VPWR VPWR _5314_/A sky130_fd_sc_hd__or2_1
X_9081_ _9705_/CLK _9081_/D VGND VGND VPWR VPWR _9081_/Q sky130_fd_sc_hd__dfxtp_1
X_6293_ _6293_/A VGND VGND VPWR VPWR _6293_/Y sky130_fd_sc_hd__clkinv_2
X_5244_ _9608_/Q _5241_/Y hold379/X _5241_/A VGND VGND VPWR VPWR _5244_/X sky130_fd_sc_hd__o22a_1
XFILLER_142_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8032_ _8157_/A _8032_/B VGND VGND VPWR VPWR _8175_/A sky130_fd_sc_hd__or2_1
XFILLER_152_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5175_ _9655_/Q _5170_/A _8964_/A1 _5170_/Y VGND VGND VPWR VPWR _9655_/D sky130_fd_sc_hd__a22o_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8934_ _8933_/X _9189_/Q _9096_/Q VGND VGND VPWR VPWR _8934_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8865_ _9192_/Q _9832_/Q _9829_/Q VGND VGND VPWR VPWR _8865_/X sky130_fd_sc_hd__mux2_2
X_7816_ _7816_/A _7816_/B VGND VGND VPWR VPWR _7816_/Y sky130_fd_sc_hd__nand2_1
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8796_ _8796_/A VGND VGND VPWR VPWR _8796_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4959_ _4657_/Y _8999_/S _4958_/Y hold708/X _4657_/A VGND VGND VPWR VPWR _9753_/D
+ sky130_fd_sc_hd__a32o_1
X_7747_ _7748_/B _7747_/B VGND VGND VPWR VPWR _7747_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7678_ _6749_/Y _7485_/X _6676_/Y _7486_/X _7677_/X VGND VGND VPWR VPWR _7694_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9417_ _9695_/CLK _9417_/D _9537_/SET_B VGND VGND VPWR VPWR _9417_/Q sky130_fd_sc_hd__dfrtp_1
X_6629_ _9591_/Q VGND VGND VPWR VPWR _8827_/A sky130_fd_sc_hd__clkinv_8
XFILLER_20_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9348_ _9483_/CLK _9348_/D _9727_/SET_B VGND VGND VPWR VPWR _9348_/Q sky130_fd_sc_hd__dfstp_1
X_9279_ _9392_/CLK _9279_/D _9537_/SET_B VGND VGND VPWR VPWR _9279_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput380 _9082_/Q VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_126_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput391 _9055_/Q VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6980_ _9105_/Q VGND VGND VPWR VPWR _6981_/B sky130_fd_sc_hd__inv_2
XFILLER_38_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5931_ _9178_/Q _5929_/A _8964_/A1 _5929_/Y VGND VGND VPWR VPWR _9178_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8650_ _8538_/A _8557_/B _8347_/B _8059_/C _8489_/X VGND VGND VPWR VPWR _8651_/A
+ sky130_fd_sc_hd__o311a_1
X_5862_ _9230_/Q _5860_/A _8964_/A1 _5860_/Y VGND VGND VPWR VPWR _9230_/D sky130_fd_sc_hd__a22o_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5793_ _9276_/Q _5788_/A _8964_/A1 _5788_/Y VGND VGND VPWR VPWR _9276_/D sky130_fd_sc_hd__a22o_1
X_8581_ _8581_/A _8763_/C _8580_/X VGND VGND VPWR VPWR _8747_/D sky130_fd_sc_hd__or3b_2
X_7601_ _6322_/Y _7527_/X _6347_/Y _7528_/X VGND VGND VPWR VPWR _7601_/X sky130_fd_sc_hd__o22a_1
XFILLER_61_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4813_ _9790_/Q VGND VGND VPWR VPWR _4813_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7532_ _7532_/A _7532_/B _7532_/C _7532_/D VGND VGND VPWR VPWR _7532_/Y sky130_fd_sc_hd__nand4_4
X_4744_ _6142_/B _4801_/B VGND VGND VPWR VPWR _5797_/B sky130_fd_sc_hd__or2_4
XFILLER_147_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9202_ _9318_/CLK _9202_/D _9571_/SET_B VGND VGND VPWR VPWR _9202_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4675_ _4675_/A VGND VGND VPWR VPWR _4675_/X sky130_fd_sc_hd__clkbuf_1
X_7463_ _4800_/Y _7507_/A _4872_/Y _7508_/A _7462_/X VGND VGND VPWR VPWR _7482_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6414_ _6398_/Y _5826_/B _6401_/X _6407_/X _6413_/X VGND VGND VPWR VPWR _6506_/C
+ sky130_fd_sc_hd__o2111a_1
X_7394_ _6553_/Y _7155_/A _6588_/Y _7156_/A _7393_/X VGND VGND VPWR VPWR _7397_/C
+ sky130_fd_sc_hd__o221a_1
X_6345_ _9693_/Q VGND VGND VPWR VPWR _6345_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_162_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9133_ _9751_/CLK _9133_/D _6014_/X VGND VGND VPWR VPWR _9133_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_103_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9064_ _9064_/CLK _9064_/D VGND VGND VPWR VPWR _9064_/Q sky130_fd_sc_hd__dfxtp_1
X_6276_ _6276_/A VGND VGND VPWR VPWR _6276_/Y sky130_fd_sc_hd__clkinv_4
X_5227_ _9619_/Q _5226_/Y _8971_/X hold666/X VGND VGND VPWR VPWR _9619_/D sky130_fd_sc_hd__o22a_1
X_8015_ _8431_/A VGND VGND VPWR VPWR _8429_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput108 sram_ro_data[23] VGND VGND VPWR VPWR _6131_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput119 sram_ro_data[4] VGND VGND VPWR VPWR _6482_/A sky130_fd_sc_hd__clkbuf_1
X_5158_ _5158_/A VGND VGND VPWR VPWR _5159_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5089_ _9009_/X _9707_/Q _5101_/S VGND VGND VPWR VPWR _5090_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8917_ _7209_/Y _9676_/Q _9001_/S VGND VGND VPWR VPWR _8917_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8848_ _8848_/A VGND VGND VPWR VPWR _8848_/X sky130_fd_sc_hd__clkbuf_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8779_ _8178_/B _8596_/B _8778_/X _8670_/X VGND VGND VPWR VPWR _8779_/Y sky130_fd_sc_hd__o211ai_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_81 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_70 _6536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold307 hold307/A VGND VGND VPWR VPWR hold308/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold318 _5117_/X VGND VGND VPWR VPWR hold319/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold329 hold329/A VGND VGND VPWR VPWR _9515_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6130_ _6130_/A VGND VGND VPWR VPWR _6130_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_112_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _9119_/Q _6060_/A hold516/X _6060_/Y VGND VGND VPWR VPWR _6061_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _9133_/Q _9132_/Q _9134_/Q VGND VGND VPWR VPWR _5012_/X sky130_fd_sc_hd__o21a_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9820_ _9832_/CLK _9820_/D _9821_/SET_B VGND VGND VPWR VPWR _9820_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9751_ _9751_/CLK _9751_/D _4970_/X VGND VGND VPWR VPWR _9751_/Q sky130_fd_sc_hd__dfrtp_1
X_6963_ _9255_/Q VGND VGND VPWR VPWR _6963_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9682_ _4471_/A1 _9682_/D _6177_/A VGND VGND VPWR VPWR _9682_/Q sky130_fd_sc_hd__dfrtp_1
X_8702_ _8702_/A _8702_/B _8702_/C VGND VGND VPWR VPWR _8702_/X sky130_fd_sc_hd__or3_1
XFILLER_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6894_ _6892_/Y _4598_/B _8850_/A _4848_/X VGND VGND VPWR VPWR _6894_/X sky130_fd_sc_hd__o22a_1
XFILLER_34_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5914_ _5889_/X _8936_/X _8960_/X _9191_/Q VGND VGND VPWR VPWR _9191_/D sky130_fd_sc_hd__o22a_1
X_8633_ _8552_/A _8540_/A _7918_/B _8439_/A VGND VGND VPWR VPWR _8633_/Y sky130_fd_sc_hd__o211ai_1
X_5845_ _9241_/Q _5841_/A _6067_/B1 _5841_/Y VGND VGND VPWR VPWR _9241_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8564_ _8105_/C _8105_/B _8563_/Y _8056_/B VGND VGND VPWR VPWR _8569_/B sky130_fd_sc_hd__a31o_1
X_5776_ _9284_/Q _5773_/A hold217/X _5773_/Y VGND VGND VPWR VPWR _9284_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8495_ _8707_/A _8495_/B _8495_/C _8649_/C VGND VGND VPWR VPWR _8497_/A sky130_fd_sc_hd__or4_1
X_4727_ _4947_/A _4764_/B VGND VGND VPWR VPWR _5698_/B sky130_fd_sc_hd__or2_4
X_7515_ _7515_/A VGND VGND VPWR VPWR _7515_/X sky130_fd_sc_hd__buf_6
XFILLER_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7446_ _4794_/Y _7493_/A _4879_/Y _7494_/A VGND VGND VPWR VPWR _7446_/X sky130_fd_sc_hd__o22a_1
X_4658_ _9760_/Q _4657_/A _8942_/X _4657_/Y VGND VGND VPWR VPWR _9760_/D sky130_fd_sc_hd__a22o_1
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__buf_2
XFILLER_174_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9116_ _9514_/CLK _9116_/D _9727_/SET_B VGND VGND VPWR VPWR _9116_/Q sky130_fd_sc_hd__dfrtp_1
X_7377_ _6705_/Y _7070_/A _6693_/Y _7166_/X _7376_/X VGND VGND VPWR VPWR _7384_/A
+ sky130_fd_sc_hd__o221a_1
X_4589_ _9796_/Q _4587_/A hold510/X _4587_/Y VGND VGND VPWR VPWR _9796_/D sky130_fd_sc_hd__a22o_1
X_6328_ _9735_/Q VGND VGND VPWR VPWR _6328_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9047_ _9640_/Q _8829_/A VGND VGND VPWR VPWR _9047_/Z sky130_fd_sc_hd__ebufn_1
X_6259_ _6257_/Y _4545_/B _6258_/Y _4854_/X VGND VGND VPWR VPWR _6259_/X sky130_fd_sc_hd__o22a_2
XFILLER_130_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5630_ _5630_/A VGND VGND VPWR VPWR _5630_/Y sky130_fd_sc_hd__inv_2
X_5561_ _5561_/A VGND VGND VPWR VPWR _5561_/Y sky130_fd_sc_hd__clkinv_2
X_7300_ _6104_/Y _7135_/X _6145_/Y _7136_/X _7299_/X VGND VGND VPWR VPWR _7319_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_129_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8280_ _8280_/A _8302_/B VGND VGND VPWR VPWR _8616_/B sky130_fd_sc_hd__nor2_1
X_4512_ _4512_/A VGND VGND VPWR VPWR _4513_/A sky130_fd_sc_hd__clkbuf_4
X_5492_ _9440_/Q _5484_/A _6008_/B1 _5484_/Y VGND VGND VPWR VPWR _9440_/D sky130_fd_sc_hd__a22o_1
Xhold126 hold126/A VGND VGND VPWR VPWR _9563_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold115 hold115/A VGND VGND VPWR VPWR hold116/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 hold104/A VGND VGND VPWR VPWR _9462_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7231_ _7231_/A _7231_/B _7231_/C VGND VGND VPWR VPWR _7231_/Y sky130_fd_sc_hd__nand3_4
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold159 hold159/A VGND VGND VPWR VPWR hold160/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _5309_/X VGND VGND VPWR VPWR hold138/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 hold148/A VGND VGND VPWR VPWR _9338_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7162_ _7162_/A VGND VGND VPWR VPWR _7162_/X sky130_fd_sc_hd__buf_6
X_6113_ _6109_/Y _5367_/B _6110_/Y _5301_/B _6112_/X VGND VGND VPWR VPWR _6127_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7145_/A _7168_/A _7137_/A _7138_/A VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__and4_1
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6044_/A VGND VGND VPWR VPWR _6044_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7995_ _8479_/B _8205_/A VGND VGND VPWR VPWR _8627_/B sky130_fd_sc_hd__nor2_2
X_9803_ _9810_/CLK _9803_/D _7042_/B VGND VGND VPWR VPWR _9803_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_39_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6946_ _9407_/Q VGND VGND VPWR VPWR _6946_/Y sky130_fd_sc_hd__inv_2
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9734_ _9734_/CLK _9734_/D _9731_/SET_B VGND VGND VPWR VPWR _9734_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9665_ _9730_/CLK _9665_/D _9730_/SET_B VGND VGND VPWR VPWR _9665_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6877_ _6875_/Y _4511_/B _6876_/Y _5282_/B VGND VGND VPWR VPWR _6877_/X sky130_fd_sc_hd__o22a_1
X_5828_ _5828_/A VGND VGND VPWR VPWR _5828_/Y sky130_fd_sc_hd__inv_2
X_8616_ _8616_/A _8616_/B _8616_/C VGND VGND VPWR VPWR _8772_/D sky130_fd_sc_hd__or3_1
X_9596_ _9600_/CLK _9596_/D _9821_/SET_B VGND VGND VPWR VPWR _9596_/Q sky130_fd_sc_hd__dfrtp_1
X_8547_ _8639_/D _8641_/D _8699_/C _8546_/X VGND VGND VPWR VPWR _8551_/A sky130_fd_sc_hd__or4b_4
X_5759_ _9097_/Q _7072_/A _5741_/Y VGND VGND VPWR VPWR _5759_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8478_ _8478_/A _8478_/B VGND VGND VPWR VPWR _8529_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7429_ _7429_/A _7429_/B _7429_/C VGND VGND VPWR VPWR _7429_/Y sky130_fd_sc_hd__nand3_1
Xhold671 _5234_/X VGND VGND VPWR VPWR _9612_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold660 _5473_/X VGND VGND VPWR VPWR _9453_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_150_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold682 _4823_/B VGND VGND VPWR VPWR _4508_/B sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold693 _9611_/Q VGND VGND VPWR VPWR hold710/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput209 _8796_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_95_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6800_ input5/X VGND VGND VPWR VPWR _6800_/Y sky130_fd_sc_hd__inv_2
X_7780_ _9108_/Q _7780_/B VGND VGND VPWR VPWR _7780_/X sky130_fd_sc_hd__and2_1
X_4992_ _4992_/A VGND VGND VPWR VPWR _4992_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6731_ _9429_/Q VGND VGND VPWR VPWR _6731_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6662_ _9338_/Q VGND VGND VPWR VPWR _7204_/A sky130_fd_sc_hd__clkinv_4
XFILLER_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9450_ _9582_/CLK _9450_/D _9727_/SET_B VGND VGND VPWR VPWR _9450_/Q sky130_fd_sc_hd__dfstp_1
X_5613_ _9360_/Q _5611_/A hold510/X _5611_/Y VGND VGND VPWR VPWR _5613_/X sky130_fd_sc_hd__a22o_1
X_9381_ _9522_/CLK _9381_/D _9537_/SET_B VGND VGND VPWR VPWR _9381_/Q sky130_fd_sc_hd__dfstp_1
X_8401_ _8401_/A _8401_/B VGND VGND VPWR VPWR _8616_/C sky130_fd_sc_hd__or2_1
XFILLER_176_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8332_ _8648_/B _8332_/B VGND VGND VPWR VPWR _8333_/C sky130_fd_sc_hd__or2_1
X_6593_ _9513_/Q VGND VGND VPWR VPWR _8833_/A sky130_fd_sc_hd__inv_8
XFILLER_129_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5544_ _5544_/A VGND VGND VPWR VPWR _5545_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8263_ _8277_/A _8540_/A _8264_/C VGND VGND VPWR VPWR _8265_/A sky130_fd_sc_hd__or3_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5475_ _5475_/A VGND VGND VPWR VPWR _5475_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7214_ _8791_/A _7144_/X _8787_/A _7145_/X _7213_/X VGND VGND VPWR VPWR _7221_/A
+ sky130_fd_sc_hd__o221a_2
X_8194_ _8594_/A _8420_/B VGND VGND VPWR VPWR _8409_/A sky130_fd_sc_hd__nor2_1
X_7145_ _7145_/A VGND VGND VPWR VPWR _7145_/X sky130_fd_sc_hd__buf_4
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7076_ _7424_/B _7144_/A _7174_/A _7160_/A VGND VGND VPWR VPWR _7094_/A sky130_fd_sc_hd__and4_1
XFILLER_104_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6027_ _9131_/Q _6026_/A _8948_/X _6026_/Y VGND VGND VPWR VPWR _9131_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7978_ _8243_/A _8552_/A _7977_/Y VGND VGND VPWR VPWR _7978_/X sky130_fd_sc_hd__o21ba_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9717_ _9723_/CLK _9717_/D _6177_/A VGND VGND VPWR VPWR _9717_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9679_/CLK sky130_fd_sc_hd__clkbuf_16
X_6929_ _9376_/Q VGND VGND VPWR VPWR _6929_/Y sky130_fd_sc_hd__clkinv_2
X_9648_ _9651_/CLK _9648_/D _9563_/SET_B VGND VGND VPWR VPWR _9648_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9579_ _9579_/CLK _9579_/D _7042_/B VGND VGND VPWR VPWR _9579_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_46_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9817_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold490 hold490/A VGND VGND VPWR VPWR hold491/A sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_89_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5260_ _9598_/Q _5257_/A hold217/A _5257_/Y VGND VGND VPWR VPWR _9598_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5191_ _5191_/A VGND VGND VPWR VPWR _5192_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8950_ _7742_/X _9124_/Q _9093_/Q VGND VGND VPWR VPWR _8950_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7901_ _8302_/A VGND VGND VPWR VPWR _7901_/Y sky130_fd_sc_hd__clkinv_2
X_8881_ _4971_/A hold176/X _8987_/S VGND VGND VPWR VPWR _8881_/X sky130_fd_sc_hd__mux2_8
XFILLER_36_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7832_ _8125_/A _8126_/A VGND VGND VPWR VPWR _7833_/A sky130_fd_sc_hd__or2_1
XFILLER_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7763_ _7763_/A _9017_/S VGND VGND VPWR VPWR _7764_/A sky130_fd_sc_hd__and2_1
X_4975_ _9750_/Q VGND VGND VPWR VPWR _4975_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6714_ _6712_/Y _5036_/B _6713_/Y _5858_/B VGND VGND VPWR VPWR _6714_/X sky130_fd_sc_hd__o22a_1
X_9502_ _9729_/CLK _9502_/D _9727_/SET_B VGND VGND VPWR VPWR _9502_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9433_ _9522_/CLK _9433_/D _9563_/SET_B VGND VGND VPWR VPWR _9433_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7694_ _7694_/A _7694_/B _7694_/C _7694_/D VGND VGND VPWR VPWR _7694_/Y sky130_fd_sc_hd__nand4_2
XFILLER_192_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6645_ _6640_/Y _5274_/B _8807_/A _5559_/B _6644_/X VGND VGND VPWR VPWR _6658_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9364_ _9643_/CLK _9364_/D _9563_/SET_B VGND VGND VPWR VPWR _9364_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6576_ _9766_/Q VGND VGND VPWR VPWR _6576_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5527_ _9418_/Q _5523_/A _8959_/A1 _5523_/Y VGND VGND VPWR VPWR _9418_/D sky130_fd_sc_hd__a22o_1
X_8315_ _8315_/A _8757_/B VGND VGND VPWR VPWR _8317_/A sky130_fd_sc_hd__or2_1
X_9295_ _9297_/CLK _9295_/D _9730_/SET_B VGND VGND VPWR VPWR _9295_/Q sky130_fd_sc_hd__dfrtp_2
X_8246_ _8246_/A _8682_/A VGND VGND VPWR VPWR _8720_/A sky130_fd_sc_hd__nor2_1
XFILLER_133_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5458_ _9465_/Q _5456_/X hold516/X _5457_/Y VGND VGND VPWR VPWR _5458_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8177_ _8177_/A _8400_/A _8684_/A _8401_/A VGND VGND VPWR VPWR _8181_/A sky130_fd_sc_hd__or4_1
X_5389_ _5474_/A _5389_/B VGND VGND VPWR VPWR _5390_/A sky130_fd_sc_hd__or2_1
XFILLER_99_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7128_ _7128_/A _7129_/B _7129_/C VGND VGND VPWR VPWR _7182_/A sky130_fd_sc_hd__or3_2
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7059_ _7113_/A _7118_/C VGND VGND VPWR VPWR _7127_/B sky130_fd_sc_hd__or2_1
XFILLER_59_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_160 _6534_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_182 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_171 _8829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_193 _6794_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4760_/A VGND VGND VPWR VPWR _6165_/A sky130_fd_sc_hd__buf_8
X_4691_ _9396_/Q VGND VGND VPWR VPWR _4691_/Y sky130_fd_sc_hd__clkinv_2
X_6430_ _9509_/Q VGND VGND VPWR VPWR _6430_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6361_ _9561_/Q VGND VGND VPWR VPWR _6361_/Y sky130_fd_sc_hd__inv_2
X_8100_ _8126_/A VGND VGND VPWR VPWR _8105_/B sky130_fd_sc_hd__inv_2
X_5312_ _6083_/A VGND VGND VPWR VPWR _5474_/A sky130_fd_sc_hd__clkbuf_4
X_9080_ _9705_/CLK _9080_/D VGND VGND VPWR VPWR _9080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6292_ _6287_/Y _5378_/B _6288_/Y _4892_/X _6291_/X VGND VGND VPWR VPWR _6311_/A
+ sky130_fd_sc_hd__o221a_1
X_5243_ _9609_/Q _5241_/Y hold569/X _5241_/A VGND VGND VPWR VPWR _5243_/X sky130_fd_sc_hd__o22a_1
XFILLER_130_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8031_ _8180_/A VGND VGND VPWR VPWR _8592_/A sky130_fd_sc_hd__buf_2
X_5174_ _9656_/Q _5170_/A _8959_/A1 _5170_/Y VGND VGND VPWR VPWR _9656_/D sky130_fd_sc_hd__a22o_1
Xhold19 hold19/A VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8933_ _7385_/Y _9671_/Q _9001_/S VGND VGND VPWR VPWR _8933_/X sky130_fd_sc_hd__mux2_1
X_8864_ _9218_/Q _9121_/Q _9829_/Q VGND VGND VPWR VPWR _8864_/X sky130_fd_sc_hd__mux2_4
X_7815_ _8260_/B VGND VGND VPWR VPWR _8009_/A sky130_fd_sc_hd__inv_2
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8795_ _8795_/A VGND VGND VPWR VPWR _8796_/A sky130_fd_sc_hd__clkbuf_1
X_4958_ _4958_/A _4958_/B _4958_/C VGND VGND VPWR VPWR _4958_/Y sky130_fd_sc_hd__nand3_4
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7746_ _9126_/Q _7745_/B _9127_/Q VGND VGND VPWR VPWR _7747_/B sky130_fd_sc_hd__a21oi_1
X_4889_ _4889_/A VGND VGND VPWR VPWR _4889_/Y sky130_fd_sc_hd__inv_4
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7677_ _6760_/Y _7487_/X _6716_/Y _7488_/X VGND VGND VPWR VPWR _7677_/X sky130_fd_sc_hd__o22a_1
XFILLER_124_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9416_ _9416_/CLK _9416_/D _9731_/SET_B VGND VGND VPWR VPWR _9416_/Q sky130_fd_sc_hd__dfrtp_1
X_6628_ _9599_/Q VGND VGND VPWR VPWR _6628_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9347_ _9483_/CLK _9347_/D _9727_/SET_B VGND VGND VPWR VPWR _9347_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6559_ _9178_/Q VGND VGND VPWR VPWR _6559_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_193_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9278_ _9392_/CLK _9278_/D _9563_/SET_B VGND VGND VPWR VPWR _9278_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput370 _9073_/Q VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_2
X_8229_ _8229_/A _8229_/B VGND VGND VPWR VPWR _8648_/B sky130_fd_sc_hd__nor2_1
XFILLER_105_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput381 _9083_/Q VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_126_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5930_ _9179_/Q _5929_/A _8959_/A1 _5929_/Y VGND VGND VPWR VPWR _9179_/D sky130_fd_sc_hd__a22o_1
XFILLER_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7600_ _6315_/Y _7519_/X _6302_/Y _7520_/X _7599_/X VGND VGND VPWR VPWR _7603_/C
+ sky130_fd_sc_hd__o221a_1
X_5861_ _9231_/Q _5860_/A _8959_/A1 _5860_/Y VGND VGND VPWR VPWR _9231_/D sky130_fd_sc_hd__a22o_1
X_8580_ _8625_/A _8580_/B _8580_/C _8580_/D VGND VGND VPWR VPWR _8580_/X sky130_fd_sc_hd__or4_1
X_5792_ _9277_/Q _5788_/A _8959_/A1 _5788_/Y VGND VGND VPWR VPWR _9277_/D sky130_fd_sc_hd__a22o_1
X_4812_ _4812_/A _4812_/B _4812_/C _4812_/D VGND VGND VPWR VPWR _4958_/B sky130_fd_sc_hd__and4_1
XFILLER_21_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7531_ _7531_/A _7531_/B _7531_/C _7531_/D VGND VGND VPWR VPWR _7532_/D sky130_fd_sc_hd__and4_1
X_4743_ _9268_/Q VGND VGND VPWR VPWR _4743_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7462_ _4936_/Y _7509_/A _4950_/Y _7510_/A VGND VGND VPWR VPWR _7462_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9201_ _9326_/CLK _9201_/D _9571_/SET_B VGND VGND VPWR VPWR _9201_/Q sky130_fd_sc_hd__dfrtp_1
X_6413_ _6408_/Y _5687_/B _7424_/A _5658_/B _6412_/X VGND VGND VPWR VPWR _6413_/X
+ sky130_fd_sc_hd__o221a_1
X_4674_ _4969_/A VGND VGND VPWR VPWR _4675_/A sky130_fd_sc_hd__clkbuf_1
X_7393_ _6608_/Y _7056_/A _6541_/Y _7157_/A VGND VGND VPWR VPWR _7393_/X sky130_fd_sc_hd__o22a_1
X_6344_ _6339_/Y _5786_/B _6340_/Y _5706_/B _6343_/X VGND VGND VPWR VPWR _6356_/A
+ sky130_fd_sc_hd__o221a_1
X_9132_ _8879_/A1 _9132_/D _6018_/X VGND VGND VPWR VPWR _9132_/Q sky130_fd_sc_hd__dfrtp_1
X_6275_ _9541_/Q VGND VGND VPWR VPWR _6275_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9063_ _9723_/CLK _9063_/D VGND VGND VPWR VPWR _9063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5226_ _5226_/A VGND VGND VPWR VPWR _5226_/Y sky130_fd_sc_hd__inv_2
X_8014_ _8421_/B _8134_/A VGND VGND VPWR VPWR _8431_/A sky130_fd_sc_hd__or2_4
XFILLER_142_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput109 sram_ro_data[24] VGND VGND VPWR VPWR _4853_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5157_ _6196_/A _5179_/B VGND VGND VPWR VPWR _5158_/A sky130_fd_sc_hd__or2_1
XFILLER_69_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5088_ _5088_/A VGND VGND VPWR VPWR _9708_/D sky130_fd_sc_hd__clkbuf_1
X_8916_ _8915_/X _9180_/Q _9096_/Q VGND VGND VPWR VPWR _8916_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8847_ _8847_/A input1/X VGND VGND VPWR VPWR _8848_/A sky130_fd_sc_hd__and2_1
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8778_ _8205_/A _8592_/A _8070_/X _8453_/Y VGND VGND VPWR VPWR _8778_/X sky130_fd_sc_hd__o211a_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7729_ _7729_/A _7729_/B _7729_/C _7729_/D VGND VGND VPWR VPWR _7730_/D sky130_fd_sc_hd__and4_1
XFILLER_184_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_93 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_60 _8807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold308 hold308/A VGND VGND VPWR VPWR _9393_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold319 hold319/A VGND VGND VPWR VPWR hold320/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6060_/A VGND VGND VPWR VPWR _6060_/Y sky130_fd_sc_hd__inv_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _9742_/Q _9741_/Q VGND VGND VPWR VPWR _6023_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6962_ _6957_/Y _5687_/B _6958_/Y _5771_/B _6961_/X VGND VGND VPWR VPWR _6975_/A
+ sky130_fd_sc_hd__o221a_1
X_9750_ _8879_/A1 _9750_/D _4980_/X VGND VGND VPWR VPWR _9750_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8701_ _8701_/A _8701_/B _8701_/C _7932_/X VGND VGND VPWR VPWR _8769_/C sky130_fd_sc_hd__or4b_2
X_9681_ _9833_/CLK _9681_/D _9730_/SET_B VGND VGND VPWR VPWR _9681_/Q sky130_fd_sc_hd__dfrtp_1
X_6893_ _9602_/Q VGND VGND VPWR VPWR _8850_/A sky130_fd_sc_hd__inv_2
X_5913_ _5889_/X _8938_/X _8960_/X _9192_/Q VGND VGND VPWR VPWR _9192_/D sky130_fd_sc_hd__o22a_1
XFILLER_179_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8632_ _8647_/B _8585_/Y _8606_/X _8631_/X VGND VGND VPWR VPWR _8632_/Y sky130_fd_sc_hd__o211ai_1
X_5844_ _9242_/Q _5841_/A hold217/A _5841_/Y VGND VGND VPWR VPWR _9242_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8563_ _8563_/A _8563_/B VGND VGND VPWR VPWR _8563_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5775_ _9285_/Q _5773_/A _6065_/B1 _5773_/Y VGND VGND VPWR VPWR _9285_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7514_ _7514_/A VGND VGND VPWR VPWR _7514_/X sky130_fd_sc_hd__buf_6
XFILLER_147_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8494_ _8280_/A _7903_/X _8053_/A _8171_/B VGND VGND VPWR VPWR _8649_/C sky130_fd_sc_hd__o22ai_1
X_4726_ _9306_/Q VGND VGND VPWR VPWR _4726_/Y sky130_fd_sc_hd__inv_2
X_4657_ _4657_/A VGND VGND VPWR VPWR _4657_/Y sky130_fd_sc_hd__inv_2
X_7445_ _7478_/C _7473_/A _7471_/C VGND VGND VPWR VPWR _7494_/A sky130_fd_sc_hd__or3_2
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__buf_6
X_7376_ _6663_/Y _7167_/X _6781_/Y _7168_/X VGND VGND VPWR VPWR _7376_/X sky130_fd_sc_hd__o22a_1
X_6327_ _9333_/Q VGND VGND VPWR VPWR _6327_/Y sky130_fd_sc_hd__clkinv_2
X_9115_ _9577_/CLK _9115_/D _9571_/SET_B VGND VGND VPWR VPWR _9115_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4588_ _9797_/Q _4587_/A hold516/X _4587_/Y VGND VGND VPWR VPWR _9797_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9046_ _9639_/Q _8827_/A VGND VGND VPWR VPWR _9046_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6258_ _6258_/A VGND VGND VPWR VPWR _6258_/Y sky130_fd_sc_hd__inv_2
X_5209_ _9630_/Q _5203_/A _8975_/A1 _5203_/Y VGND VGND VPWR VPWR _9630_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6189_ _6189_/A _6189_/B VGND VGND VPWR VPWR _6189_/X sky130_fd_sc_hd__or2_4
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5560_ _5560_/A VGND VGND VPWR VPWR _5561_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5491_ _9441_/Q _5484_/A _6067_/B1 _5484_/Y VGND VGND VPWR VPWR _9441_/D sky130_fd_sc_hd__a22o_1
X_4511_ _5201_/A _4511_/B VGND VGND VPWR VPWR _4511_/X sky130_fd_sc_hd__or2_1
Xhold105 _5186_/X VGND VGND VPWR VPWR hold106/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 hold116/A VGND VGND VPWR VPWR _9633_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7230_ _7230_/A _7230_/B _7230_/C _7230_/D VGND VGND VPWR VPWR _7231_/C sky130_fd_sc_hd__and4_1
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold127 _5415_/X VGND VGND VPWR VPWR hold128/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _5567_/X VGND VGND VPWR VPWR hold150/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 hold138/A VGND VGND VPWR VPWR hold139/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7161_ _7161_/A VGND VGND VPWR VPWR _7161_/X sky130_fd_sc_hd__buf_6
X_6112_ _6112_/A _6112_/B VGND VGND VPWR VPWR _6112_/X sky130_fd_sc_hd__or2_1
XFILLER_98_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7092_/A _7127_/B VGND VGND VPWR VPWR _7138_/A sky130_fd_sc_hd__or2_2
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6071_/A VGND VGND VPWR VPWR _6044_/A sky130_fd_sc_hd__clkbuf_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7994_ _8179_/A VGND VGND VPWR VPWR _8205_/A sky130_fd_sc_hd__buf_6
XFILLER_81_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9802_ _9810_/CLK _9802_/D _7042_/B VGND VGND VPWR VPWR _9802_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_54_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6945_ _9329_/Q VGND VGND VPWR VPWR _6945_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9733_ _9734_/CLK _9733_/D _9731_/SET_B VGND VGND VPWR VPWR _9733_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_9664_ _9730_/CLK _9664_/D _9730_/SET_B VGND VGND VPWR VPWR _9664_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6876_ _9579_/Q VGND VGND VPWR VPWR _6876_/Y sky130_fd_sc_hd__clkinv_2
X_5827_ _5827_/A VGND VGND VPWR VPWR _5828_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_139_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8615_ _8615_/A _8615_/B _8615_/C VGND VGND VPWR VPWR _8684_/D sky130_fd_sc_hd__or3_1
X_9595_ _9832_/CLK _9595_/D _9821_/SET_B VGND VGND VPWR VPWR _9595_/Q sky130_fd_sc_hd__dfrtp_2
X_8546_ _8543_/X _8546_/B _8546_/C VGND VGND VPWR VPWR _8546_/X sky130_fd_sc_hd__and3b_1
XFILLER_6_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5758_ _5758_/A VGND VGND VPWR VPWR _9292_/D sky130_fd_sc_hd__clkinv_2
XFILLER_163_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8477_ _8678_/B _8477_/B VGND VGND VPWR VPWR _8478_/B sky130_fd_sc_hd__or2_1
X_4709_ _4933_/B _4865_/B VGND VGND VPWR VPWR _5979_/B sky130_fd_sc_hd__or2_4
XFILLER_162_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5689_ _5689_/A VGND VGND VPWR VPWR _5689_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7428_ _7428_/A _7428_/B _7428_/C _7428_/D VGND VGND VPWR VPWR _7429_/C sky130_fd_sc_hd__and4_1
XFILLER_150_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold650 _8975_/X VGND VGND VPWR VPWR hold650/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7359_ _6887_/Y _5756_/X _6933_/Y _7071_/A _7358_/X VGND VGND VPWR VPWR _7362_/C
+ sky130_fd_sc_hd__o221a_1
Xhold661 _5130_/X VGND VGND VPWR VPWR _9683_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold672 _9125_/Q VGND VGND VPWR VPWR hold672/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold683 _4913_/B VGND VGND VPWR VPWR _4925_/A sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_1_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold694 _7016_/Y VGND VGND VPWR VPWR _8851_/A sky130_fd_sc_hd__buf_6
XFILLER_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9029_ _9029_/A _8793_/A VGND VGND VPWR VPWR _9029_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_89_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4991_ _5017_/A VGND VGND VPWR VPWR _4992_/A sky130_fd_sc_hd__clkbuf_1
X_6730_ _9784_/Q VGND VGND VPWR VPWR _6730_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6661_ _6180_/A _6660_/Y _9081_/Q _6180_/Y VGND VGND VPWR VPWR _9081_/D sky130_fd_sc_hd__o22a_1
X_5612_ _9361_/Q _5611_/A hold516/X _5611_/Y VGND VGND VPWR VPWR _5612_/X sky130_fd_sc_hd__a22o_1
X_9380_ _9522_/CLK _9380_/D _9537_/SET_B VGND VGND VPWR VPWR _9380_/Q sky130_fd_sc_hd__dfstp_1
X_8400_ _8400_/A _8400_/B VGND VGND VPWR VPWR _8684_/C sky130_fd_sc_hd__or2_1
X_6592_ _6592_/A VGND VGND VPWR VPWR _6592_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8331_ _8667_/A _8382_/B _8382_/C _8330_/X VGND VGND VPWR VPWR _8332_/B sky130_fd_sc_hd__a31o_1
XFILLER_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5543_ _5698_/A _5543_/B VGND VGND VPWR VPWR _5544_/A sky130_fd_sc_hd__or2_1
XFILLER_160_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8262_ _8608_/B _8256_/Y _8259_/Y _8151_/C _8261_/Y VGND VGND VPWR VPWR _8266_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_117_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5474_ _5474_/A _5474_/B VGND VGND VPWR VPWR _5474_/X sky130_fd_sc_hd__or2_1
XFILLER_172_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7213_ _8785_/A _7071_/C _7733_/A _7146_/X VGND VGND VPWR VPWR _7213_/X sky130_fd_sc_hd__o22a_1
X_8193_ _8193_/A _8716_/A VGND VGND VPWR VPWR _8195_/A sky130_fd_sc_hd__or2_1
XFILLER_132_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7144_ _7144_/A VGND VGND VPWR VPWR _7144_/X sky130_fd_sc_hd__buf_4
XFILLER_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7075_ _7128_/A _7129_/B _7091_/C VGND VGND VPWR VPWR _7160_/A sky130_fd_sc_hd__or3_4
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6026_ _6026_/A VGND VGND VPWR VPWR _6026_/Y sky130_fd_sc_hd__inv_2
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7977_ _8135_/A _7977_/B VGND VGND VPWR VPWR _7977_/Y sky130_fd_sc_hd__nand2_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9716_ _9731_/CLK _9716_/D _9731_/SET_B VGND VGND VPWR VPWR _9716_/Q sky130_fd_sc_hd__dfrtp_1
X_6928_ _9241_/Q VGND VGND VPWR VPWR _6928_/Y sky130_fd_sc_hd__inv_2
X_9647_ _9651_/CLK _9647_/D _9689_/SET_B VGND VGND VPWR VPWR _9647_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6859_ _6854_/Y _6058_/B _6855_/Y _5359_/B _6858_/X VGND VGND VPWR VPWR _6860_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9578_ _9819_/CLK _9578_/D _7042_/B VGND VGND VPWR VPWR _9578_/Q sky130_fd_sc_hd__dfrtp_1
X_8529_ _8529_/A _8528_/X VGND VGND VPWR VPWR _8530_/A sky130_fd_sc_hd__or2b_1
XFILLER_136_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold480 hold480/A VGND VGND VPWR VPWR _9602_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_145_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold491 hold491/A VGND VGND VPWR VPWR hold491/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_92_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _4467_/A1
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_126_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5190_ _5378_/A _6353_/A VGND VGND VPWR VPWR _5191_/A sky130_fd_sc_hd__or2_1
X_7900_ _8347_/A VGND VGND VPWR VPWR _8341_/B sky130_fd_sc_hd__inv_2
XFILLER_110_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8880_ input85/X _4971_/A _9668_/Q VGND VGND VPWR VPWR _8880_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7831_ _8580_/C _8558_/B VGND VGND VPWR VPWR _8126_/A sky130_fd_sc_hd__or2_2
XFILLER_63_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4974_ _9751_/Q VGND VGND VPWR VPWR _4974_/Y sky130_fd_sc_hd__inv_2
X_7762_ _7759_/Y _7758_/Y _9742_/Q _7761_/Y VGND VGND VPWR VPWR _7762_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6713_ _9229_/Q VGND VGND VPWR VPWR _6713_/Y sky130_fd_sc_hd__clkinv_2
X_7693_ _7693_/A _7693_/B _7693_/C _7693_/D VGND VGND VPWR VPWR _7694_/D sky130_fd_sc_hd__and4_1
X_9501_ _9729_/CLK _9501_/D _9727_/SET_B VGND VGND VPWR VPWR _9501_/Q sky130_fd_sc_hd__dfrtp_1
X_9432_ _9522_/CLK _9432_/D _9537_/SET_B VGND VGND VPWR VPWR _9432_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6644_ _8813_/A _4937_/X _6643_/Y _5466_/B VGND VGND VPWR VPWR _6644_/X sky130_fd_sc_hd__o22a_1
X_9363_ _9643_/CLK _9363_/D _9563_/SET_B VGND VGND VPWR VPWR _9363_/Q sky130_fd_sc_hd__dfstp_1
X_6575_ _9677_/Q VGND VGND VPWR VPWR _6575_/Y sky130_fd_sc_hd__inv_2
X_5526_ _9419_/Q _5523_/A hold577/A _5523_/Y VGND VGND VPWR VPWR _5526_/X sky130_fd_sc_hd__a22o_1
X_8314_ _8314_/A _8702_/B _8538_/A VGND VGND VPWR VPWR _8757_/B sky130_fd_sc_hd__nor3_2
X_9294_ _9297_/CLK _9294_/D _9730_/SET_B VGND VGND VPWR VPWR _9294_/Q sky130_fd_sc_hd__dfstp_1
X_8245_ _8264_/C VGND VGND VPWR VPWR _8682_/A sky130_fd_sc_hd__buf_2
X_5457_ _5457_/A VGND VGND VPWR VPWR _5457_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5388_ _9510_/Q _5380_/A hold601/A _5380_/Y VGND VGND VPWR VPWR _5388_/X sky130_fd_sc_hd__a22o_1
X_8176_ _8178_/B _8182_/B VGND VGND VPWR VPWR _8401_/A sky130_fd_sc_hd__nor2_1
X_7127_ _7127_/A _7127_/B VGND VGND VPWR VPWR _7180_/A sky130_fd_sc_hd__or2_1
XFILLER_59_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7058_ _7084_/C VGND VGND VPWR VPWR _7091_/C sky130_fd_sc_hd__buf_2
XFILLER_86_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6009_ _6017_/A VGND VGND VPWR VPWR _6010_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_161 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_150 _4919_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _8829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_183 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 _8815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4690_ _4949_/A _4865_/B VGND VGND VPWR VPWR _5902_/B sky130_fd_sc_hd__or2_4
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6360_ _9548_/Q VGND VGND VPWR VPWR _6360_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5311_ _9562_/Q _5303_/A hold601/A _5303_/Y VGND VGND VPWR VPWR _5311_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8030_ _8091_/B _8032_/B VGND VGND VPWR VPWR _8180_/A sky130_fd_sc_hd__or2_2
X_6291_ _6289_/Y _4611_/B _6290_/Y _6117_/X VGND VGND VPWR VPWR _6291_/X sky130_fd_sc_hd__o22a_1
X_5242_ _9610_/Q _5241_/Y hold563/X _5241_/A VGND VGND VPWR VPWR _5242_/X sky130_fd_sc_hd__o22a_1
XFILLER_130_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5173_ _9657_/Q _5170_/A hold696/A _5170_/Y VGND VGND VPWR VPWR _5173_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_30_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9418_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_4
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_45_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9819_/CLK sky130_fd_sc_hd__clkbuf_16
X_8932_ _8931_/X _9188_/Q _9096_/Q VGND VGND VPWR VPWR _8932_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8863_ _9099_/Q _9120_/Q _9829_/Q VGND VGND VPWR VPWR _8863_/X sky130_fd_sc_hd__mux2_1
X_7814_ _7869_/A _7874_/B _5964_/X VGND VGND VPWR VPWR _8260_/B sky130_fd_sc_hd__o21ai_2
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8794_ _8794_/A VGND VGND VPWR VPWR _8794_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7745_ _9126_/Q _7745_/B _9127_/Q VGND VGND VPWR VPWR _7748_/B sky130_fd_sc_hd__and3_1
X_4957_ _4957_/A _4957_/B _4957_/C _4957_/D VGND VGND VPWR VPWR _4958_/C sky130_fd_sc_hd__and4_2
X_7676_ _7676_/A _7676_/B _7676_/C _7676_/D VGND VGND VPWR VPWR _7676_/Y sky130_fd_sc_hd__nand4_2
X_4888_ _4933_/A _4947_/A VGND VGND VPWR VPWR _5359_/B sky130_fd_sc_hd__or2_4
XFILLER_192_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9415_ _9416_/CLK _9415_/D _9731_/SET_B VGND VGND VPWR VPWR _9415_/Q sky130_fd_sc_hd__dfstp_1
X_6627_ _6622_/Y _4585_/B _6623_/Y _6117_/X _6626_/X VGND VGND VPWR VPWR _6627_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6558_ _9409_/Q VGND VGND VPWR VPWR _8841_/A sky130_fd_sc_hd__inv_4
XFILLER_117_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9346_ _9483_/CLK _9346_/D _9727_/SET_B VGND VGND VPWR VPWR _9346_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9277_ _9392_/CLK _9277_/D _9537_/SET_B VGND VGND VPWR VPWR _9277_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5509_ _9430_/Q _5507_/A _6065_/B1 _5507_/Y VGND VGND VPWR VPWR _9430_/D sky130_fd_sc_hd__a22o_1
X_6489_ _9147_/Q VGND VGND VPWR VPWR _6489_/Y sky130_fd_sc_hd__clkinv_2
X_8228_ _8228_/A VGND VGND VPWR VPWR _8692_/B sky130_fd_sc_hd__inv_2
XFILLER_121_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput371 _9063_/Q VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput360 _9062_/Q VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8159_ _8436_/A _8421_/B _8158_/A VGND VGND VPWR VPWR _8159_/X sky130_fd_sc_hd__or3b_1
Xoutput382 _9064_/Q VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_99_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5860_ _5860_/A VGND VGND VPWR VPWR _5860_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4811_ _4811_/A _4811_/B _4811_/C _4811_/D VGND VGND VPWR VPWR _4812_/D sky130_fd_sc_hd__and4_1
XFILLER_73_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5791_ _9278_/Q _5788_/A hold577/A _5788_/Y VGND VGND VPWR VPWR _5791_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7530_ _6920_/Y _7525_/X _7178_/A _7526_/X _7529_/X VGND VGND VPWR VPWR _7531_/D
+ sky130_fd_sc_hd__o221a_1
X_4742_ _4939_/A _4764_/B VGND VGND VPWR VPWR _5706_/B sky130_fd_sc_hd__or2_4
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4673_ _9755_/Q _4657_/A _8993_/X _4657_/Y VGND VGND VPWR VPWR _9755_/D sky130_fd_sc_hd__a22o_1
X_7461_ _7467_/A _7477_/A _7478_/D VGND VGND VPWR VPWR _7510_/A sky130_fd_sc_hd__or3_2
X_9200_ _9225_/CLK _9200_/D _9731_/SET_B VGND VGND VPWR VPWR _9200_/Q sky130_fd_sc_hd__dfrtp_1
X_6412_ _6410_/Y _5698_/B _7248_/A _5636_/B VGND VGND VPWR VPWR _6412_/X sky130_fd_sc_hd__o22a_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7392_ _6620_/Y _7149_/A _6508_/Y _7150_/A _7391_/X VGND VGND VPWR VPWR _7397_/B
+ sky130_fd_sc_hd__o221a_1
X_6343_ _6341_/Y _6112_/B _6342_/Y _5609_/B VGND VGND VPWR VPWR _6343_/X sky130_fd_sc_hd__o22a_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9131_ net399_3/A _9131_/D _6022_/X VGND VGND VPWR VPWR _9131_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9062_ _9062_/CLK _9062_/D VGND VGND VPWR VPWR _9062_/Q sky130_fd_sc_hd__dfxtp_1
X_6274_ _9787_/Q VGND VGND VPWR VPWR _6274_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5225_ hold665/X _6353_/A _5250_/A _9019_/X VGND VGND VPWR VPWR _5226_/A sky130_fd_sc_hd__a211o_4
X_8013_ _8013_/A VGND VGND VPWR VPWR _8596_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_130_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5156_ _5770_/A _9019_/S VGND VGND VPWR VPWR _5179_/B sky130_fd_sc_hd__or2_1
XFILLER_96_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5087_ _9010_/X _9708_/Q _5101_/S VGND VGND VPWR VPWR _5088_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8915_ _7187_/Y _9675_/Q _9001_/S VGND VGND VPWR VPWR _8915_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8846_ _8846_/A VGND VGND VPWR VPWR _8846_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _9148_/Q _5981_/A _8975_/A1 _5981_/Y VGND VGND VPWR VPWR _9148_/D sky130_fd_sc_hd__a22o_1
X_8777_ _8777_/A _8777_/B _8777_/C _8777_/D VGND VGND VPWR VPWR _8777_/X sky130_fd_sc_hd__or4_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7728_ _6472_/Y _7525_/A _7424_/A _7526_/A _7727_/X VGND VGND VPWR VPWR _7729_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_50 _6793_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _4471_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_83 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7659_ _6897_/Y _7487_/X _6933_/Y _7488_/X VGND VGND VPWR VPWR _7659_/X sky130_fd_sc_hd__o22a_1
XANTENNA_94 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9329_ _9391_/CLK _9329_/D _9563_/SET_B VGND VGND VPWR VPWR _9329_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold309 _5791_/X VGND VGND VPWR VPWR hold310/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _9723_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_98_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5010_/A VGND VGND VPWR VPWR _5010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8700_ _8718_/B _8700_/B VGND VGND VPWR VPWR _8701_/B sky130_fd_sc_hd__or2_1
X_6961_ _6959_/Y _5698_/B _6960_/Y _5990_/B VGND VGND VPWR VPWR _6961_/X sky130_fd_sc_hd__o22a_1
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5912_ _9193_/Q _5904_/A _8975_/A1 _5904_/Y VGND VGND VPWR VPWR _9193_/D sky130_fd_sc_hd__a22o_1
X_9680_ _9730_/CLK _9680_/D _9797_/SET_B VGND VGND VPWR VPWR _9680_/Q sky130_fd_sc_hd__dfrtp_1
X_6892_ _9783_/Q VGND VGND VPWR VPWR _6892_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8631_ _8692_/B _8692_/C _8693_/B _8630_/X VGND VGND VPWR VPWR _8631_/X sky130_fd_sc_hd__or4b_2
X_5843_ _9243_/Q _5841_/A _6065_/B1 _5841_/Y VGND VGND VPWR VPWR _9243_/D sky130_fd_sc_hd__a22o_1
XFILLER_179_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8562_ _8514_/Y _8559_/Y _8560_/X _8486_/B VGND VGND VPWR VPWR _8654_/B sky130_fd_sc_hd__a31o_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5774_ _9286_/Q _5773_/A _6064_/B1 _5773_/Y VGND VGND VPWR VPWR _9286_/D sky130_fd_sc_hd__a22o_1
X_7513_ _7513_/A VGND VGND VPWR VPWR _7513_/X sky130_fd_sc_hd__buf_6
XFILLER_159_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8493_ _8493_/A _8725_/A VGND VGND VPWR VPWR _8495_/C sky130_fd_sc_hd__or2_1
X_4725_ _4725_/A _4725_/B _4725_/C _4725_/D VGND VGND VPWR VPWR _4958_/A sky130_fd_sc_hd__and4_1
XFILLER_190_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7444_ _7479_/A _9293_/Q _7467_/A _9297_/Q VGND VGND VPWR VPWR _7493_/A sky130_fd_sc_hd__or4_2
X_4656_ _4656_/A VGND VGND VPWR VPWR _4657_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_162_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_6
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _6091_/A sky130_fd_sc_hd__clkbuf_1
X_7375_ _7375_/A _7375_/B _7375_/C _7375_/D VGND VGND VPWR VPWR _7385_/B sky130_fd_sc_hd__and4_1
X_4587_ _4587_/A VGND VGND VPWR VPWR _4587_/Y sky130_fd_sc_hd__inv_2
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__clkbuf_2
X_6326_ _6318_/Y _5570_/B _6319_/Y _5826_/B _6325_/X VGND VGND VPWR VPWR _6338_/B
+ sky130_fd_sc_hd__o221a_1
X_9114_ _9514_/CLK _9114_/D _9727_/SET_B VGND VGND VPWR VPWR _9114_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9045_ _9638_/Q _8825_/A VGND VGND VPWR VPWR _9045_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6257_ _9810_/Q VGND VGND VPWR VPWR _6257_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6188_ _9694_/Q VGND VGND VPWR VPWR _6188_/Y sky130_fd_sc_hd__inv_2
X_5208_ _9631_/Q _5203_/A hold593/X _5203_/Y VGND VGND VPWR VPWR _9631_/D sky130_fd_sc_hd__a22o_1
X_5139_ _9678_/Q _5135_/A _8959_/A1 _5135_/Y VGND VGND VPWR VPWR _9678_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8829_ _8829_/A VGND VGND VPWR VPWR _8830_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4510_ _4913_/B _4827_/A VGND VGND VPWR VPWR _4511_/B sky130_fd_sc_hd__or2_4
X_5490_ _9442_/Q _5484_/A hold217/X _5484_/Y VGND VGND VPWR VPWR _9442_/D sky130_fd_sc_hd__a22o_1
Xhold117 _9743_/Q VGND VGND VPWR VPWR hold118/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 hold106/A VGND VGND VPWR VPWR hold107/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 hold128/A VGND VGND VPWR VPWR hold129/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 hold139/A VGND VGND VPWR VPWR _9564_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7160_ _7160_/A VGND VGND VPWR VPWR _7160_/X sky130_fd_sc_hd__buf_6
X_6111_ _9439_/Q VGND VGND VPWR VPWR _6112_/A sky130_fd_sc_hd__inv_2
XFILLER_98_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7108_/C _7129_/A _7091_/C VGND VGND VPWR VPWR _7137_/A sky130_fd_sc_hd__or3_4
XFILLER_98_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _9126_/Q _6026_/A _8951_/X _6026_/Y VGND VGND VPWR VPWR _9126_/D sky130_fd_sc_hd__a22o_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9801_ _4471_/A1 _9801_/D _6177_/A VGND VGND VPWR VPWR _9801_/Q sky130_fd_sc_hd__dfrtp_4
X_7993_ _8236_/A _8674_/A VGND VGND VPWR VPWR _8179_/A sky130_fd_sc_hd__or2_4
XFILLER_93_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6944_ _9136_/Q VGND VGND VPWR VPWR _6944_/Y sky130_fd_sc_hd__clkinv_2
X_9732_ _9734_/CLK _9732_/D _9731_/SET_B VGND VGND VPWR VPWR _9732_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9663_ _9734_/CLK _9663_/D _9731_/SET_B VGND VGND VPWR VPWR _9663_/Q sky130_fd_sc_hd__dfrtp_1
X_8614_ _8683_/B _8761_/A _8614_/C _8719_/C VGND VGND VPWR VPWR _8618_/A sky130_fd_sc_hd__or4_4
XFILLER_62_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6875_ _9821_/Q VGND VGND VPWR VPWR _6875_/Y sky130_fd_sc_hd__inv_6
XFILLER_167_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5826_ _5847_/A _5826_/B VGND VGND VPWR VPWR _5827_/A sky130_fd_sc_hd__or2_1
XFILLER_139_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9594_ _9827_/CLK _9594_/D _9797_/SET_B VGND VGND VPWR VPWR _9594_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8545_ _8383_/A _8281_/B _8280_/A _8540_/B _7949_/X VGND VGND VPWR VPWR _8546_/C
+ sky130_fd_sc_hd__o221a_1
X_5757_ _7025_/A _5719_/Y _5752_/Y _5723_/A _5756_/X VGND VGND VPWR VPWR _5758_/A
+ sky130_fd_sc_hd__o32a_1
X_8476_ _8476_/A _8678_/C VGND VGND VPWR VPWR _8477_/B sky130_fd_sc_hd__nor2_1
X_4708_ _4750_/A _4708_/B _4750_/C _4750_/D VGND VGND VPWR VPWR _6117_/B sky130_fd_sc_hd__or4_4
X_5688_ _5688_/A VGND VGND VPWR VPWR _5689_/A sky130_fd_sc_hd__clkbuf_4
X_7427_ _6435_/Y _7180_/A _6374_/Y _7181_/A _7426_/X VGND VGND VPWR VPWR _7428_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_135_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4639_ _9765_/Q hold673/X hold217/X _4636_/Y VGND VGND VPWR VPWR _9765_/D sky130_fd_sc_hd__a22o_1
Xhold651 _5249_/X VGND VGND VPWR VPWR _9603_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_118_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7358_ _7358_/A _7380_/B VGND VGND VPWR VPWR _7358_/X sky130_fd_sc_hd__or2_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold640 _4560_/X VGND VGND VPWR VPWR _9803_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold662 _5396_/X VGND VGND VPWR VPWR _9505_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold695 _8851_/Y VGND VGND VPWR VPWR _8855_/B sky130_fd_sc_hd__clkbuf_1
X_7289_ _6225_/Y _7071_/D _6185_/Y _7166_/X _7288_/X VGND VGND VPWR VPWR _7296_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6309_ _6307_/Y _5521_/B _6308_/Y _5559_/B VGND VGND VPWR VPWR _6309_/X sky130_fd_sc_hd__o22a_1
Xhold673 _4636_/A VGND VGND VPWR VPWR hold673/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold684 _5129_/X VGND VGND VPWR VPWR _9684_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_9028_ _9028_/A _8791_/A VGND VGND VPWR VPWR _9028_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4990_ _9749_/Q _4989_/A _9748_/Q _4989_/Y VGND VGND VPWR VPWR _9749_/D sky130_fd_sc_hd__a22o_1
X_6660_ _6660_/A _6660_/B _6660_/C _6660_/D VGND VGND VPWR VPWR _6660_/Y sky130_fd_sc_hd__nand4_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5611_ _5611_/A VGND VGND VPWR VPWR _5611_/Y sky130_fd_sc_hd__inv_2
X_6591_ _6586_/Y _5543_/B _6587_/Y _5428_/B _6590_/X VGND VGND VPWR VPWR _6598_/C
+ sky130_fd_sc_hd__o221a_1
X_5542_ _9406_/Q _5534_/A _8975_/A1 _5534_/Y VGND VGND VPWR VPWR _9406_/D sky130_fd_sc_hd__a22o_1
X_8330_ _8382_/C _8432_/B _8382_/B _8329_/X VGND VGND VPWR VPWR _8330_/X sky130_fd_sc_hd__a31o_1
XFILLER_129_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8261_ _8321_/C _8353_/B VGND VGND VPWR VPWR _8261_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5473_ _9453_/Q _5468_/A _6008_/B1 _5468_/Y VGND VGND VPWR VPWR _5473_/X sky130_fd_sc_hd__a22o_1
X_7212_ _8831_/A _7135_/X _8833_/A _7136_/X _7211_/X VGND VGND VPWR VPWR _7231_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8192_ _8594_/A _8682_/B VGND VGND VPWR VPWR _8716_/A sky130_fd_sc_hd__nor2_1
XFILLER_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7143_ _6856_/Y _7135_/X _6818_/Y _7136_/X _7142_/X VGND VGND VPWR VPWR _7187_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7074_ _7092_/A _7121_/B VGND VGND VPWR VPWR _7174_/A sky130_fd_sc_hd__or2_2
XFILLER_113_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6025_ _9093_/Q _6024_/X _6053_/B VGND VGND VPWR VPWR _6026_/A sky130_fd_sc_hd__o21ai_4
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7976_ _8324_/C _7873_/C _8324_/B _8745_/A _7975_/X VGND VGND VPWR VPWR _7977_/B
+ sky130_fd_sc_hd__a311oi_1
X_9715_ _9736_/CLK _9715_/D _9731_/SET_B VGND VGND VPWR VPWR _9715_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ _9176_/Q VGND VGND VPWR VPWR _6927_/Y sky130_fd_sc_hd__inv_2
X_9646_ _9651_/CLK _9646_/D _9563_/SET_B VGND VGND VPWR VPWR _9646_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6858_ _6856_/Y _5340_/B _6857_/Y _5436_/B VGND VGND VPWR VPWR _6858_/X sky130_fd_sc_hd__o22a_1
X_5809_ _9266_/Q _5807_/A hold510/X _5807_/Y VGND VGND VPWR VPWR _9266_/D sky130_fd_sc_hd__a22o_1
X_9577_ _9577_/CLK _9577_/D _9571_/SET_B VGND VGND VPWR VPWR _9577_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8528_ _8556_/B _8527_/X VGND VGND VPWR VPWR _8528_/X sky130_fd_sc_hd__or2b_1
X_6789_ _6784_/Y _6112_/B _6785_/Y _5935_/B _6788_/X VGND VGND VPWR VPWR _6790_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8459_ _8709_/B _8619_/A VGND VGND VPWR VPWR _8728_/A sky130_fd_sc_hd__or2_1
XFILLER_145_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold470 hold470/A VGND VGND VPWR VPWR hold470/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold481 _5251_/S VGND VGND VPWR VPWR hold482/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold492 _8981_/X VGND VGND VPWR VPWR hold493/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7830_ _7860_/A _7860_/B _8580_/B VGND VGND VPWR VPWR _8558_/B sky130_fd_sc_hd__o21ai_1
XFILLER_63_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4973_ _9090_/Q _4973_/B VGND VGND VPWR VPWR _4973_/Y sky130_fd_sc_hd__nand2_1
X_7761_ _7759_/Y _7758_/Y _9742_/Q VGND VGND VPWR VPWR _7761_/Y sky130_fd_sc_hd__a21oi_1
X_6712_ _9732_/Q VGND VGND VPWR VPWR _6712_/Y sky130_fd_sc_hd__inv_2
X_7692_ _6781_/Y _7525_/X _7380_/A _7526_/X _7691_/X VGND VGND VPWR VPWR _7693_/D
+ sky130_fd_sc_hd__o221a_1
X_9500_ _9579_/CLK _9500_/D _9727_/SET_B VGND VGND VPWR VPWR _9500_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9431_ _9431_/CLK _9431_/D _9797_/SET_B VGND VGND VPWR VPWR _9431_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6643_ _9456_/Q VGND VGND VPWR VPWR _6643_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9362_ _9421_/CLK _9362_/D _9537_/SET_B VGND VGND VPWR VPWR _9362_/Q sky130_fd_sc_hd__dfstp_1
X_6574_ _9503_/Q VGND VGND VPWR VPWR _6574_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_192_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5525_ _9420_/Q _5523_/A hold510/X _5523_/Y VGND VGND VPWR VPWR _5525_/X sky130_fd_sc_hd__a22o_1
X_8313_ _8313_/A _8548_/B VGND VGND VPWR VPWR _8315_/A sky130_fd_sc_hd__or2_1
X_9293_ _9297_/CLK _9293_/D _9730_/SET_B VGND VGND VPWR VPWR _9293_/Q sky130_fd_sc_hd__dfrtp_4
X_8244_ _8244_/A VGND VGND VPWR VPWR _8518_/B sky130_fd_sc_hd__inv_2
X_5456_ _5456_/A VGND VGND VPWR VPWR _5456_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_133_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5387_ _9511_/Q _5380_/A _6067_/B1 _5380_/Y VGND VGND VPWR VPWR _9511_/D sky130_fd_sc_hd__a22o_1
X_8175_ _8175_/A _8682_/B VGND VGND VPWR VPWR _8684_/A sky130_fd_sc_hd__nor2_1
XFILLER_113_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7126_ _4838_/Y _5756_/A _4864_/Y _7061_/A _7125_/X VGND VGND VPWR VPWR _7132_/C
+ sky130_fd_sc_hd__o221a_1
X_7057_ _9292_/Q _9291_/Q VGND VGND VPWR VPWR _7084_/C sky130_fd_sc_hd__or2_2
XFILLER_59_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6008_ _9135_/Q _6000_/A _6008_/B1 _6000_/Y VGND VGND VPWR VPWR _9135_/D sky130_fd_sc_hd__a22o_1
XFILLER_74_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ _7903_/X _8361_/A _7956_/Y _8534_/A _8362_/A VGND VGND VPWR VPWR _7959_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9629_ _4471_/A1 _9629_/D _6177_/A VGND VGND VPWR VPWR _9629_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_140 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_151 _4938_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 input89/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_173 _8833_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_162 _6902_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_195 _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5310_ _9563_/Q _5303_/A hold593/A _5303_/Y VGND VGND VPWR VPWR _5310_/X sky130_fd_sc_hd__a22o_1
X_6290_ input8/X VGND VGND VPWR VPWR _6290_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5241_ _5241_/A VGND VGND VPWR VPWR _5241_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5172_ _9658_/Q _5170_/A hold510/X _5170_/Y VGND VGND VPWR VPWR _5172_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8931_ _7363_/Y _9670_/Q _9001_/S VGND VGND VPWR VPWR _8931_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_opt_1_0_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR clkbuf_leaf_5_csclk/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8862_ _9259_/Q _9111_/Q _9829_/Q VGND VGND VPWR VPWR _8862_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7813_ _7789_/B _7812_/Y _7874_/B _7812_/A VGND VGND VPWR VPWR _7936_/A sky130_fd_sc_hd__o22a_1
X_8793_ _8793_/A VGND VGND VPWR VPWR _8794_/A sky130_fd_sc_hd__clkbuf_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7744_ _9126_/Q _7745_/B _9126_/Q _7745_/B VGND VGND VPWR VPWR _7744_/X sky130_fd_sc_hd__o2bb2a_1
X_4956_ _4956_/A _4956_/B _4956_/C _4956_/D VGND VGND VPWR VPWR _4957_/D sky130_fd_sc_hd__and4_1
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7675_ _7675_/A _7675_/B _7675_/C _7675_/D VGND VGND VPWR VPWR _7676_/D sky130_fd_sc_hd__and4_1
XFILLER_20_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4887_ _9526_/Q VGND VGND VPWR VPWR _4887_/Y sky130_fd_sc_hd__inv_2
X_6626_ _6624_/Y _4890_/X _8837_/A _5455_/B VGND VGND VPWR VPWR _6626_/X sky130_fd_sc_hd__o22a_4
X_9414_ _9418_/CLK _9414_/D _9731_/SET_B VGND VGND VPWR VPWR _9414_/Q sky130_fd_sc_hd__dfstp_1
X_6557_ _6557_/A _6557_/B _6557_/C _6557_/D VGND VGND VPWR VPWR _6660_/B sky130_fd_sc_hd__and4_1
X_9345_ _9729_/CLK _9345_/D _9727_/SET_B VGND VGND VPWR VPWR _9345_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5508_ _9431_/Q _5507_/A _6064_/B1 _5507_/Y VGND VGND VPWR VPWR _9431_/D sky130_fd_sc_hd__a22o_1
X_9276_ _9392_/CLK _9276_/D _9537_/SET_B VGND VGND VPWR VPWR _9276_/Q sky130_fd_sc_hd__dfrtp_1
X_6488_ _9223_/Q VGND VGND VPWR VPWR _6488_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8227_ _8227_/A VGND VGND VPWR VPWR _8714_/C sky130_fd_sc_hd__inv_2
Xoutput361 _9056_/Q VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput350 _9805_/Q VGND VGND VPWR VPWR sram_ro_addr[1] sky130_fd_sc_hd__buf_2
X_5439_ _9478_/Q _5438_/A _6064_/B1 _5438_/Y VGND VGND VPWR VPWR _9478_/D sky130_fd_sc_hd__a22o_1
Xoutput383 _9084_/Q VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_2
Xoutput372 _9074_/Q VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_126_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8158_ _8158_/A _8158_/B VGND VGND VPWR VPWR _8435_/A sky130_fd_sc_hd__nand2_2
XFILLER_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7109_ _4948_/Y _7151_/A _4932_/Y _7152_/A VGND VGND VPWR VPWR _7109_/X sky130_fd_sc_hd__o22a_1
XFILLER_59_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8089_ _8596_/A _8429_/A _8088_/X VGND VGND VPWR VPWR _8089_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4810_ _4800_/Y _5786_/B _4802_/Y _6353_/A _4809_/X VGND VGND VPWR VPWR _4811_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5790_ _9279_/Q _5788_/A hold510/X _5788_/Y VGND VGND VPWR VPWR _5790_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4741_ _9298_/Q VGND VGND VPWR VPWR _4741_/Y sky130_fd_sc_hd__inv_4
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4672_ _4672_/A VGND VGND VPWR VPWR _4672_/X sky130_fd_sc_hd__clkbuf_1
X_7460_ _7460_/A _7476_/B _7478_/D VGND VGND VPWR VPWR _7509_/A sky130_fd_sc_hd__or3_2
X_6411_ _9340_/Q VGND VGND VPWR VPWR _7248_/A sky130_fd_sc_hd__inv_2
X_7391_ _6635_/Y _7151_/A _6581_/Y _7152_/A VGND VGND VPWR VPWR _7391_/X sky130_fd_sc_hd__o22a_1
X_9130_ net399_3/A _9130_/D _6029_/X VGND VGND VPWR VPWR _9130_/Q sky130_fd_sc_hd__dfrtp_2
X_6342_ _9359_/Q VGND VGND VPWR VPWR _6342_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9061_ _9718_/CLK _9061_/D VGND VGND VPWR VPWR _9061_/Q sky130_fd_sc_hd__dfxtp_1
X_6273_ _6271_/Y _5329_/B _6272_/Y _4511_/B VGND VGND VPWR VPWR _6273_/X sky130_fd_sc_hd__o22a_1
XFILLER_115_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8012_ _8137_/B _8157_/A VGND VGND VPWR VPWR _8013_/A sky130_fd_sc_hd__or2_1
X_5224_ _9620_/Q _5216_/Y _8972_/X _5216_/A VGND VGND VPWR VPWR _9620_/D sky130_fd_sc_hd__o22a_1
XFILLER_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5155_ hold1/A VGND VGND VPWR VPWR _9019_/S sky130_fd_sc_hd__clkinv_8
X_5086_ _5086_/A VGND VGND VPWR VPWR _5101_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_84_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8914_ _8913_/X _9217_/Q _9096_/Q VGND VGND VPWR VPWR _8914_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8845_ _8845_/A _8875_/S VGND VGND VPWR VPWR _8846_/A sky130_fd_sc_hd__and2_1
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5988_ _9149_/Q _5981_/A _8969_/A1 _5981_/Y VGND VGND VPWR VPWR _9149_/D sky130_fd_sc_hd__a22o_1
X_8776_ _8776_/A _8776_/B _8776_/C _8776_/D VGND VGND VPWR VPWR _8777_/B sky130_fd_sc_hd__or4_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4939_ _4939_/A _4953_/B VGND VGND VPWR VPWR _5406_/B sky130_fd_sc_hd__or2_4
X_7727_ _6460_/Y _7527_/A _6410_/Y _7528_/A VGND VGND VPWR VPWR _7727_/X sky130_fd_sc_hd__o22a_1
XANTENNA_40 _6427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7658_ _7658_/A _7658_/B _7658_/C _7658_/D VGND VGND VPWR VPWR _7658_/Y sky130_fd_sc_hd__nand4_2
XANTENNA_84 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_62 _5290_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _6830_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _8821_/A _4869_/X _6608_/Y _5436_/B VGND VGND VPWR VPWR _6609_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_95 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7589_ _6313_/Y _7493_/X _6272_/Y _7494_/X VGND VGND VPWR VPWR _7589_/X sky130_fd_sc_hd__o22a_1
X_9328_ _9391_/CLK _9328_/D _9563_/SET_B VGND VGND VPWR VPWR _9328_/Q sky130_fd_sc_hd__dfstp_1
Xclkbuf_opt_1_0_wb_clk_i _9297_/CLK VGND VGND VPWR VPWR clkbuf_opt_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9259_ _9322_/CLK _9259_/D _9797_/SET_B VGND VGND VPWR VPWR _9259_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_44_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9686_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6960_ _9144_/Q VGND VGND VPWR VPWR _6960_/Y sky130_fd_sc_hd__clkinv_2
X_5911_ _9194_/Q _5904_/A _8969_/A1 _5904_/Y VGND VGND VPWR VPWR _9194_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6891_ _9589_/Q VGND VGND VPWR VPWR _6891_/Y sky130_fd_sc_hd__inv_6
X_8630_ _8762_/B _8630_/B _8747_/A _8723_/A VGND VGND VPWR VPWR _8630_/X sky130_fd_sc_hd__or4_1
XFILLER_61_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5842_ _9244_/Q _5841_/A _6064_/B1 _5841_/Y VGND VGND VPWR VPWR _9244_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8561_ _8558_/Y _8559_/Y _8560_/X _8495_/C VGND VGND VPWR VPWR _8649_/A sky130_fd_sc_hd__a31o_1
X_5773_ _5773_/A VGND VGND VPWR VPWR _5773_/Y sky130_fd_sc_hd__inv_2
X_7512_ _6970_/Y _7507_/X _6818_/Y _7508_/X _7511_/X VGND VGND VPWR VPWR _7531_/A
+ sky130_fd_sc_hd__o221a_1
X_4724_ _4714_/Y _4715_/X _4716_/Y _6196_/A _4723_/X VGND VGND VPWR VPWR _4725_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8492_ _8492_/A VGND VGND VPWR VPWR _8725_/A sky130_fd_sc_hd__inv_2
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4655_ _5237_/A _4987_/B VGND VGND VPWR VPWR _4656_/A sky130_fd_sc_hd__or2_1
X_7443_ _7473_/A _7476_/B _9297_/Q VGND VGND VPWR VPWR _7492_/A sky130_fd_sc_hd__or3_2
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR _6163_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_190_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__buf_4
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR _4758_/A sky130_fd_sc_hd__clkbuf_1
X_7374_ _6677_/Y _7160_/X _6776_/Y _7064_/A _7373_/X VGND VGND VPWR VPWR _7375_/D
+ sky130_fd_sc_hd__o221a_1
X_4586_ _4586_/A VGND VGND VPWR VPWR _4587_/A sky130_fd_sc_hd__buf_2
X_9113_ _9514_/CLK _9113_/D _9571_/SET_B VGND VGND VPWR VPWR _9113_/Q sky130_fd_sc_hd__dfstp_1
X_6325_ _6320_/Y _4585_/B _6321_/Y _5367_/B _6324_/X VGND VGND VPWR VPWR _6325_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_1_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput93 sram_ro_data[0] VGND VGND VPWR VPWR _4882_/A sky130_fd_sc_hd__clkbuf_1
X_9044_ _9637_/Q _8823_/A VGND VGND VPWR VPWR _9044_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_143_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6256_ _9472_/Q VGND VGND VPWR VPWR _6256_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_67_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5207_ _9632_/Q _5203_/A hold136/X _5203_/Y VGND VGND VPWR VPWR _5207_/X sky130_fd_sc_hd__a22o_1
X_6187_ _6182_/Y _5570_/B _6183_/Y _5521_/B _6186_/X VGND VGND VPWR VPWR _6205_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5138_ _9679_/Q _5135_/A hold696/A _5135_/Y VGND VGND VPWR VPWR _9679_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5069_ _5069_/A VGND VGND VPWR VPWR _5070_/A sky130_fd_sc_hd__clkbuf_4
X_8828_ _8828_/A VGND VGND VPWR VPWR _8828_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8759_ _8682_/A _8205_/A _8682_/A _8682_/B VGND VGND VPWR VPWR _8759_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold107 hold107/A VGND VGND VPWR VPWR _9647_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold118 hold118/A VGND VGND VPWR VPWR hold119/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 hold129/A VGND VGND VPWR VPWR _9493_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6110_ _9569_/Q VGND VGND VPWR VPWR _6110_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ _7107_/B _7091_/C VGND VGND VPWR VPWR _7168_/A sky130_fd_sc_hd__or2_4
XFILLER_140_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6041_/A VGND VGND VPWR VPWR _6041_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9800_ _9800_/CLK _9800_/D _9817_/SET_B VGND VGND VPWR VPWR _9800_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_39_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7992_ _7992_/A VGND VGND VPWR VPWR _8479_/B sky130_fd_sc_hd__clkbuf_4
X_9731_ _9731_/CLK _9731_/D _9731_/SET_B VGND VGND VPWR VPWR _9731_/Q sky130_fd_sc_hd__dfstp_1
X_6943_ _6939_/Y _5112_/B _6940_/Y _4715_/X _6942_/X VGND VGND VPWR VPWR _6956_/B
+ sky130_fd_sc_hd__o221a_1
X_9662_ _9734_/CLK _9662_/D _9730_/SET_B VGND VGND VPWR VPWR _9662_/Q sky130_fd_sc_hd__dfrtp_1
X_6874_ _9532_/Q VGND VGND VPWR VPWR _6874_/Y sky130_fd_sc_hd__inv_2
X_8613_ _8613_/A _8613_/B _8613_/C VGND VGND VPWR VPWR _8719_/C sky130_fd_sc_hd__or3_2
X_5825_ _9254_/Q _5820_/A _8975_/A1 _5820_/Y VGND VGND VPWR VPWR _9254_/D sky130_fd_sc_hd__a22o_1
X_9593_ _9673_/CLK _9593_/D _9797_/SET_B VGND VGND VPWR VPWR _9593_/Q sky130_fd_sc_hd__dfrtp_2
X_8544_ _8272_/A _8540_/B _7916_/X _8275_/A VGND VGND VPWR VPWR _8546_/B sky130_fd_sc_hd__o211a_1
XFILLER_22_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5756_ _5756_/A VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__buf_6
X_8475_ _8556_/A _8475_/B VGND VGND VPWR VPWR _8678_/C sky130_fd_sc_hd__or2_1
X_5687_ _5847_/A _5687_/B VGND VGND VPWR VPWR _5688_/A sky130_fd_sc_hd__or2_1
X_4707_ _9148_/Q VGND VGND VPWR VPWR _4707_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_175_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4638_ _9766_/Q hold673/X _6065_/B1 _4636_/Y VGND VGND VPWR VPWR _9766_/D sky130_fd_sc_hd__a22o_1
X_7426_ _6460_/Y _7182_/A _6372_/Y _7183_/A VGND VGND VPWR VPWR _7426_/X sky130_fd_sc_hd__o22a_1
XFILLER_135_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold630 _5342_/A VGND VGND VPWR VPWR hold630/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4569_ _4569_/A VGND VGND VPWR VPWR _9017_/S sky130_fd_sc_hd__clkbuf_16
X_7357_ _6960_/Y _7171_/X _6832_/Y _7172_/X _7356_/X VGND VGND VPWR VPWR _7362_/B
+ sky130_fd_sc_hd__o221a_1
Xhold641 _4559_/S VGND VGND VPWR VPWR _4561_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xhold663 _4555_/X VGND VGND VPWR VPWR _9804_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold652 _4541_/X VGND VGND VPWR VPWR _4542_/A sky130_fd_sc_hd__clkdlybuf4s25_1
X_6308_ _9393_/Q VGND VGND VPWR VPWR _6308_/Y sky130_fd_sc_hd__inv_2
Xhold696 hold696/A VGND VGND VPWR VPWR hold696/X sky130_fd_sc_hd__buf_12
X_7288_ _6207_/Y _7167_/X _6243_/Y _7168_/X VGND VGND VPWR VPWR _7288_/X sky130_fd_sc_hd__o22a_1
XFILLER_103_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold674 _4634_/X VGND VGND VPWR VPWR _4635_/A sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_1_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold685 _5125_/A VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__dlymetal6s2s_1
X_9027_ _9027_/A _8789_/A VGND VGND VPWR VPWR _9027_/Z sky130_fd_sc_hd__ebufn_1
X_6239_ _6239_/A VGND VGND VPWR VPWR _6239_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5610_ _5610_/A VGND VGND VPWR VPWR _5611_/A sky130_fd_sc_hd__clkbuf_4
X_6590_ _6588_/Y _5474_/B _6589_/Y _4863_/X VGND VGND VPWR VPWR _6590_/X sky130_fd_sc_hd__o22a_1
X_5541_ _9407_/Q _5534_/A hold593/X _5534_/Y VGND VGND VPWR VPWR _9407_/D sky130_fd_sc_hd__a22o_1
XFILLER_157_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8260_ _8260_/A _8260_/B _8260_/C VGND VGND VPWR VPWR _8321_/C sky130_fd_sc_hd__or3_2
XFILLER_8_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7211_ _8799_/A _7137_/X _6522_/Y _7138_/X _7210_/X VGND VGND VPWR VPWR _7211_/X
+ sky130_fd_sc_hd__o221a_1
X_5472_ _9454_/Q _5468_/A _6067_/B1 _5468_/Y VGND VGND VPWR VPWR _9454_/D sky130_fd_sc_hd__a22o_1
X_8191_ _8191_/A _8727_/B VGND VGND VPWR VPWR _8193_/A sky130_fd_sc_hd__or2_1
X_7142_ _6922_/Y _7137_/X _6947_/Y _7138_/X _7141_/X VGND VGND VPWR VPWR _7142_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7073_ _7129_/A _7129_/B _7091_/C VGND VGND VPWR VPWR _7144_/A sky130_fd_sc_hd__or3_4
X_6024_ _9092_/Q _6024_/B _7039_/B VGND VGND VPWR VPWR _6024_/X sky130_fd_sc_hd__and3_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7975_ _8518_/A _7975_/B VGND VGND VPWR VPWR _7975_/X sky130_fd_sc_hd__or2_1
X_6926_ _9363_/Q VGND VGND VPWR VPWR _6926_/Y sky130_fd_sc_hd__clkinv_4
X_9714_ _9731_/CLK _9714_/D _9731_/SET_B VGND VGND VPWR VPWR _9714_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9645_ _9651_/CLK _9645_/D _9563_/SET_B VGND VGND VPWR VPWR _9645_/Q sky130_fd_sc_hd__dfrtp_1
X_6857_ _9475_/Q VGND VGND VPWR VPWR _6857_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5808_ _9267_/Q _5807_/A hold516/X _5807_/Y VGND VGND VPWR VPWR _9267_/D sky130_fd_sc_hd__a22o_1
X_9576_ _9576_/CLK _9576_/D _9571_/SET_B VGND VGND VPWR VPWR _9576_/Q sky130_fd_sc_hd__dfrtp_1
X_6788_ _6786_/Y _5902_/B _6787_/Y _5551_/B VGND VGND VPWR VPWR _6788_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8527_ _8527_/A _8556_/C VGND VGND VPWR VPWR _8527_/X sky130_fd_sc_hd__or2_1
XFILLER_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5739_ _9095_/Q _9097_/Q VGND VGND VPWR VPWR _5741_/A sky130_fd_sc_hd__or2_2
XFILLER_135_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8458_ _8458_/A VGND VGND VPWR VPWR _8709_/B sky130_fd_sc_hd__inv_2
X_8389_ _8419_/B _8392_/C VGND VGND VPWR VPWR _8389_/X sky130_fd_sc_hd__or2_1
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7409_ _6393_/Y _7137_/A _6471_/Y _7138_/A _7408_/X VGND VGND VPWR VPWR _7409_/X
+ sky130_fd_sc_hd__o221a_1
Xhold460 hold460/A VGND VGND VPWR VPWR _9327_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold471 _4477_/X VGND VGND VPWR VPWR hold472/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold493 hold493/A VGND VGND VPWR VPWR _4823_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold482 hold482/A VGND VGND VPWR VPWR _5253_/S sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_145_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4972_ _9134_/Q _9133_/Q _6053_/C VGND VGND VPWR VPWR _4973_/B sky130_fd_sc_hd__and3_1
X_7760_ _7759_/Y _7758_/Y _9741_/Q _9740_/Q VGND VGND VPWR VPWR _7760_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6711_ _6711_/A VGND VGND VPWR VPWR _6711_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_149_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7691_ _6683_/Y _7527_/X _6665_/Y _7528_/X VGND VGND VPWR VPWR _7691_/X sky130_fd_sc_hd__o22a_1
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6642_ _9469_/Q VGND VGND VPWR VPWR _8813_/A sky130_fd_sc_hd__inv_6
X_9430_ _9431_/CLK _9430_/D _9797_/SET_B VGND VGND VPWR VPWR _9430_/Q sky130_fd_sc_hd__dfrtp_1
X_9361_ _9391_/CLK _9361_/D _9689_/SET_B VGND VGND VPWR VPWR _9361_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6573_ _8841_/A _5532_/B _6561_/X _6567_/X _6572_/X VGND VGND VPWR VPWR _6660_/C
+ sky130_fd_sc_hd__o2111a_1
X_8312_ _8383_/A _8312_/B VGND VGND VPWR VPWR _8548_/B sky130_fd_sc_hd__nor2_1
X_5524_ _9421_/Q _5523_/A hold516/X _5523_/Y VGND VGND VPWR VPWR _5524_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_1_1_1_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_2
X_9292_ _9322_/CLK _9292_/D _9730_/SET_B VGND VGND VPWR VPWR _9292_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8243_ _8243_/A _8243_/B VGND VGND VPWR VPWR _8763_/A sky130_fd_sc_hd__nor2_4
X_5455_ _5570_/A _5455_/B VGND VGND VPWR VPWR _5456_/A sky130_fd_sc_hd__or2_1
XFILLER_172_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8174_ _8174_/A VGND VGND VPWR VPWR _8400_/A sky130_fd_sc_hd__inv_2
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5386_ _9512_/Q _5380_/A hold217/X _5380_/Y VGND VGND VPWR VPWR _5386_/X sky130_fd_sc_hd__a22o_1
X_7125_ _7125_/A _7424_/B VGND VGND VPWR VPWR _7125_/X sky130_fd_sc_hd__or2_1
XFILLER_113_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7056_ _7056_/A VGND VGND VPWR VPWR _7095_/B sky130_fd_sc_hd__buf_6
X_6007_ _9136_/Q _6000_/A _6067_/B1 _6000_/Y VGND VGND VPWR VPWR _9136_/D sky130_fd_sc_hd__a22o_1
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7958_ _8563_/B _8296_/B VGND VGND VPWR VPWR _8362_/A sky130_fd_sc_hd__or2_1
XFILLER_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7889_ _7953_/A VGND VGND VPWR VPWR _8563_/B sky130_fd_sc_hd__buf_6
X_6909_ _6909_/A _6909_/B _6909_/C _6909_/D VGND VGND VPWR VPWR _6977_/B sky130_fd_sc_hd__and4_2
X_9628_ _9751_/CLK _9628_/D _5213_/X VGND VGND VPWR VPWR _9628_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9559_ _9561_/CLK _9559_/D _7042_/B VGND VGND VPWR VPWR _9559_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_148_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold290 hold290/A VGND VGND VPWR VPWR _9303_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _9111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_130 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_152 _5570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 _7918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _9297_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_185 _5250_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_196 _6794_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5240_ _6166_/A _6353_/A _5250_/A _9018_/X VGND VGND VPWR VPWR _5241_/A sky130_fd_sc_hd__a211o_4
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5171_ _9659_/Q _5170_/A hold516/X _5170_/Y VGND VGND VPWR VPWR _5171_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8930_ _8929_/X hold709/X _9096_/Q VGND VGND VPWR VPWR _8930_/X sky130_fd_sc_hd__mux2_1
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8861_ _9281_/Q _9814_/Q _9829_/Q VGND VGND VPWR VPWR _8861_/X sky130_fd_sc_hd__mux2_4
X_7812_ _7812_/A VGND VGND VPWR VPWR _7812_/Y sky130_fd_sc_hd__inv_2
X_8792_ _8792_/A VGND VGND VPWR VPWR _8792_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7743_ _7743_/A VGND VGND VPWR VPWR _7745_/B sky130_fd_sc_hd__inv_2
X_4955_ _4946_/Y _5389_/B _4948_/Y _5329_/B _4954_/X VGND VGND VPWR VPWR _4956_/D
+ sky130_fd_sc_hd__o221a_1
X_7674_ _6927_/Y _7525_/X _7358_/A _7526_/X _7673_/X VGND VGND VPWR VPWR _7675_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4886_ _4886_/A _4886_/B _4886_/C _4886_/D VGND VGND VPWR VPWR _4957_/B sky130_fd_sc_hd__and4_1
X_9413_ _9695_/CLK _9413_/D _9689_/SET_B VGND VGND VPWR VPWR _9413_/Q sky130_fd_sc_hd__dfrtp_1
X_6625_ _9461_/Q VGND VGND VPWR VPWR _8837_/A sky130_fd_sc_hd__inv_4
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6556_ _8789_/A _5866_/B _6552_/Y _6166_/A _6555_/X VGND VGND VPWR VPWR _6557_/D
+ sky130_fd_sc_hd__o221a_1
X_9344_ _9831_/CLK _9344_/D _9727_/SET_B VGND VGND VPWR VPWR _9344_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9275_ _9392_/CLK _9275_/D _9537_/SET_B VGND VGND VPWR VPWR _9275_/Q sky130_fd_sc_hd__dfrtp_1
X_5507_ _5507_/A VGND VGND VPWR VPWR _5507_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8226_ _8226_/A VGND VGND VPWR VPWR _8556_/A sky130_fd_sc_hd__inv_2
X_6487_ _9152_/Q VGND VGND VPWR VPWR _6487_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput362 _9057_/Q VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_105_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5438_ _5438_/A VGND VGND VPWR VPWR _5438_/Y sky130_fd_sc_hd__inv_2
Xoutput340 _8864_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_2
Xoutput351 _9806_/Q VGND VGND VPWR VPWR sram_ro_addr[2] sky130_fd_sc_hd__buf_2
X_5369_ _5369_/A VGND VGND VPWR VPWR _5369_/Y sky130_fd_sc_hd__inv_2
Xoutput384 _9085_/Q VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput373 _9075_/Q VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_2
X_8157_ _8157_/A _8157_/B VGND VGND VPWR VPWR _8158_/B sky130_fd_sc_hd__or2_2
XFILLER_99_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8088_ _8088_/A _8509_/A VGND VGND VPWR VPWR _8088_/X sky130_fd_sc_hd__and2_1
X_7108_ _9288_/Q _9287_/Q _7108_/C _7129_/C VGND VGND VPWR VPWR _7152_/A sky130_fd_sc_hd__or4_4
X_7039_ _7039_/A _7039_/B VGND VGND VPWR VPWR _7039_/X sky130_fd_sc_hd__or2_1
XFILLER_47_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4925_/B _4801_/B VGND VGND VPWR VPWR _5620_/B sky130_fd_sc_hd__or2_4
XFILLER_159_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4671_ _4969_/A VGND VGND VPWR VPWR _4672_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6410_ _9310_/Q VGND VGND VPWR VPWR _6410_/Y sky130_fd_sc_hd__inv_2
X_7390_ _6535_/Y _7144_/A _6570_/Y _7145_/A _7389_/X VGND VGND VPWR VPWR _7397_/A
+ sky130_fd_sc_hd__o221a_1
X_6341_ _9437_/Q VGND VGND VPWR VPWR _6341_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9060_ _9718_/CLK _9060_/D VGND VGND VPWR VPWR _9060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6272_ _9825_/Q VGND VGND VPWR VPWR _6272_/Y sky130_fd_sc_hd__inv_6
X_8011_ _8011_/A _8139_/A VGND VGND VPWR VPWR _8157_/A sky130_fd_sc_hd__or2_1
XFILLER_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5223_ _9621_/Q _5216_/Y _8969_/X _5216_/A VGND VGND VPWR VPWR _9621_/D sky130_fd_sc_hd__o22a_1
X_5154_ _9090_/Q _4973_/B _9750_/Q _9668_/Q _4973_/Y VGND VGND VPWR VPWR _9668_/D
+ sky130_fd_sc_hd__a32o_1
X_5085_ _5085_/A _5085_/B _5085_/C _5085_/D VGND VGND VPWR VPWR _5086_/A sky130_fd_sc_hd__or4_1
XFILLER_84_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8913_ _7730_/Y _9673_/Q _9020_/S VGND VGND VPWR VPWR _8913_/X sky130_fd_sc_hd__mux2_1
X_8844_ _8844_/A VGND VGND VPWR VPWR _8844_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ _9150_/Q _5981_/A _8965_/A1 _5981_/Y VGND VGND VPWR VPWR _9150_/D sky130_fd_sc_hd__a22o_1
X_8775_ _8775_/A VGND VGND VPWR VPWR _8775_/Y sky130_fd_sc_hd__inv_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4938_ _9492_/Q VGND VGND VPWR VPWR _4938_/Y sky130_fd_sc_hd__inv_6
X_7726_ _6465_/Y _7519_/A _6371_/Y _7520_/A _7725_/X VGND VGND VPWR VPWR _7729_/C
+ sky130_fd_sc_hd__o221a_1
XANTENNA_30 _6287_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _4869_/A _4951_/B VGND VGND VPWR VPWR _4869_/X sky130_fd_sc_hd__or2_4
XANTENNA_41 _6429_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7657_ _7657_/A _7657_/B _7657_/C _7657_/D VGND VGND VPWR VPWR _7658_/D sky130_fd_sc_hd__and4_1
XANTENNA_74 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 _6875_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_63 _8864_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6608_ _9477_/Q VGND VGND VPWR VPWR _6608_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_192_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_85 input82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7588_ _6307_/Y _7485_/X _6340_/Y _7486_/X _7587_/X VGND VGND VPWR VPWR _7604_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_96 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9327_ _9574_/CLK _9327_/D _9571_/SET_B VGND VGND VPWR VPWR _9327_/Q sky130_fd_sc_hd__dfrtp_1
X_6539_ _9378_/Q VGND VGND VPWR VPWR _6539_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9258_ _9673_/CLK _9258_/D _9730_/SET_B VGND VGND VPWR VPWR _9258_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8209_ _8209_/A _8420_/B VGND VGND VPWR VPWR _8210_/A sky130_fd_sc_hd__or2_1
X_9189_ _9322_/CLK _9189_/D _9797_/SET_B VGND VGND VPWR VPWR _9189_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5910_ _9195_/Q _5904_/A _8965_/A1 _5904_/Y VGND VGND VPWR VPWR _9195_/D sky130_fd_sc_hd__a22o_1
X_6890_ _9415_/Q VGND VGND VPWR VPWR _6890_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5841_ _5841_/A VGND VGND VPWR VPWR _5841_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8560_ _8560_/A _8560_/B VGND VGND VPWR VPWR _8560_/X sky130_fd_sc_hd__or2_4
X_5772_ _5772_/A VGND VGND VPWR VPWR _5773_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7511_ _6886_/Y _7509_/X _6902_/Y _7510_/X VGND VGND VPWR VPWR _7511_/X sky130_fd_sc_hd__o22a_1
X_8491_ _8491_/A _8491_/B VGND VGND VPWR VPWR _8495_/B sky130_fd_sc_hd__or2_1
X_4723_ _4719_/Y _5927_/B _4721_/Y _5036_/B VGND VGND VPWR VPWR _4723_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7442_ _7478_/C _7477_/A _9297_/Q VGND VGND VPWR VPWR _7491_/A sky130_fd_sc_hd__or3_2
XFILLER_174_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4654_ _9092_/Q VGND VGND VPWR VPWR _4987_/B sky130_fd_sc_hd__inv_2
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_4
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR _6972_/A sky130_fd_sc_hd__clkbuf_1
X_7373_ _6671_/Y _7161_/X _6756_/Y _7162_/X VGND VGND VPWR VPWR _7373_/X sky130_fd_sc_hd__o22a_1
X_4585_ _5201_/A _4585_/B VGND VGND VPWR VPWR _4586_/A sky130_fd_sc_hd__or2_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__clkbuf_8
XFILLER_143_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9112_ _9514_/CLK _9112_/D _9727_/SET_B VGND VGND VPWR VPWR _9112_/Q sky130_fd_sc_hd__dfstp_1
X_6324_ _6322_/Y _6058_/B _6323_/Y _4915_/X VGND VGND VPWR VPWR _6324_/X sky130_fd_sc_hd__o22a_1
Xinput94 sram_ro_data[10] VGND VGND VPWR VPWR _6809_/A sky130_fd_sc_hd__clkbuf_1
X_9043_ _9636_/Q _8821_/A VGND VGND VPWR VPWR _9043_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_143_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6255_ _9173_/Q VGND VGND VPWR VPWR _6255_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_130_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5206_ _9633_/Q _5203_/A hold42/X _5203_/Y VGND VGND VPWR VPWR _5206_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6186_ _6184_/Y _4892_/X _6185_/Y _5559_/B VGND VGND VPWR VPWR _6186_/X sky130_fd_sc_hd__o22a_1
XFILLER_123_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5137_ _9680_/Q _5135_/A hold510/X _5135_/Y VGND VGND VPWR VPWR _9680_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5068_ _5201_/A _5068_/B VGND VGND VPWR VPWR _5069_/A sky130_fd_sc_hd__or2_1
XFILLER_57_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8827_ _8827_/A VGND VGND VPWR VPWR _8828_/A sky130_fd_sc_hd__clkbuf_1
X_8758_ _8758_/A _8758_/B _8758_/C _8758_/D VGND VGND VPWR VPWR _8771_/A sky130_fd_sc_hd__or4_2
XFILLER_185_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7709_ _6580_/Y _7527_/A _6541_/Y _7528_/A VGND VGND VPWR VPWR _7709_/X sky130_fd_sc_hd__o22a_1
X_8689_ _8689_/A _8758_/C _8720_/C _8763_/C VGND VGND VPWR VPWR _8689_/Y sky130_fd_sc_hd__nor4_1
XFILLER_193_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold108 _5185_/X VGND VGND VPWR VPWR hold109/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold119 hold119/A VGND VGND VPWR VPWR hold120/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6071_/A VGND VGND VPWR VPWR _6041_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_100_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7991_ _8567_/A _8580_/B _8580_/C _8125_/A VGND VGND VPWR VPWR _7992_/A sky130_fd_sc_hd__or4_1
XFILLER_26_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6942_ input62/X _4700_/Y _6941_/Y _5068_/B VGND VGND VPWR VPWR _6942_/X sky130_fd_sc_hd__o2bb2a_1
X_9730_ _9730_/CLK _9730_/D _9730_/SET_B VGND VGND VPWR VPWR _9730_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_19_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9661_ _9730_/CLK _9661_/D _9730_/SET_B VGND VGND VPWR VPWR _9661_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6873_ _6868_/Y _5144_/B _6869_/Y _5133_/B _6872_/X VGND VGND VPWR VPWR _6909_/B
+ sky130_fd_sc_hd__o221a_1
X_8612_ _8243_/B _8158_/A _8383_/B _8302_/B _8394_/B VGND VGND VPWR VPWR _8614_/C
+ sky130_fd_sc_hd__o221ai_4
X_5824_ _9255_/Q _5820_/A _8969_/A1 _5820_/Y VGND VGND VPWR VPWR _9255_/D sky130_fd_sc_hd__a22o_1
XFILLER_167_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9592_ _9832_/CLK _9592_/D _9821_/SET_B VGND VGND VPWR VPWR _9592_/Q sky130_fd_sc_hd__dfrtp_1
X_8543_ _8636_/A _8737_/C _8543_/C _8543_/D VGND VGND VPWR VPWR _8543_/X sky130_fd_sc_hd__or4_2
X_5755_ _7072_/A _7127_/A VGND VGND VPWR VPWR _5756_/A sky130_fd_sc_hd__or2_4
X_8474_ _8604_/A _8714_/C _8474_/C VGND VGND VPWR VPWR _8476_/A sky130_fd_sc_hd__or3_1
X_4706_ _4808_/B _4764_/B VGND VGND VPWR VPWR _5839_/B sky130_fd_sc_hd__or2_4
X_5686_ _5673_/A _5685_/A _9319_/Q _5685_/Y _5677_/X VGND VGND VPWR VPWR _9319_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7425_ _6422_/Y _5756_/A _6449_/Y _7061_/A _7424_/X VGND VGND VPWR VPWR _7428_/C
+ sky130_fd_sc_hd__o221a_1
X_4637_ _9767_/Q hold673/X _6064_/B1 _4636_/Y VGND VGND VPWR VPWR _9767_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold620 _5291_/X VGND VGND VPWR VPWR _5292_/A sky130_fd_sc_hd__buf_2
X_4568_ _8852_/A _8854_/A _8855_/A VGND VGND VPWR VPWR _4569_/A sky130_fd_sc_hd__and3_1
Xhold642 _5576_/X VGND VGND VPWR VPWR _9384_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold631 _5872_/X VGND VGND VPWR VPWR _9223_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_118_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold653 _4953_/A VGND VGND VPWR VPWR _4776_/B sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7356_ _6905_/Y _7173_/X _6923_/Y _7174_/X VGND VGND VPWR VPWR _7356_/X sky130_fd_sc_hd__o22a_1
Xhold697 _9629_/Q VGND VGND VPWR VPWR _8883_/S sky130_fd_sc_hd__clkbuf_2
X_6307_ _9419_/Q VGND VGND VPWR VPWR _6307_/Y sky130_fd_sc_hd__clkinv_2
Xhold664 _5228_/X VGND VGND VPWR VPWR _9618_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7287_ _7287_/A _7287_/B _7287_/C _7287_/D VGND VGND VPWR VPWR _7297_/B sky130_fd_sc_hd__and4_1
XFILLER_116_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold675 _5978_/X VGND VGND VPWR VPWR _9156_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_4499_ _4883_/A VGND VGND VPWR VPWR _6142_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold686 _5123_/X VGND VGND VPWR VPWR _5124_/A sky130_fd_sc_hd__clkdlybuf4s25_1
X_9026_ _9627_/Q _7731_/A VGND VGND VPWR VPWR _9026_/Z sky130_fd_sc_hd__ebufn_2
X_6238_ _6238_/A VGND VGND VPWR VPWR _6238_/Y sky130_fd_sc_hd__inv_2
X_6169_ _9343_/Q VGND VGND VPWR VPWR _7314_/A sky130_fd_sc_hd__clkinv_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9791_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5540_ _9408_/Q _5534_/A hold136/X _5534_/Y VGND VGND VPWR VPWR _5540_/X sky130_fd_sc_hd__a22o_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5471_ _9455_/Q _5468_/A hold217/X _5468_/Y VGND VGND VPWR VPWR _9455_/D sky130_fd_sc_hd__a22o_1
X_7210_ _8815_/A _7139_/X _8813_/A _7140_/X VGND VGND VPWR VPWR _7210_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8190_ _8205_/A _8190_/B VGND VGND VPWR VPWR _8727_/B sky130_fd_sc_hd__nor2_1
XFILLER_125_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7141_ _6884_/Y _7139_/X _6886_/Y _7140_/X VGND VGND VPWR VPWR _7141_/X sky130_fd_sc_hd__o22a_1
X_7072_ _7072_/A _7084_/C VGND VGND VPWR VPWR _7424_/B sky130_fd_sc_hd__or2_2
XFILLER_113_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6023_ _9740_/Q _6023_/B VGND VGND VPWR VPWR _7039_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7974_ _8418_/A _7974_/B VGND VGND VPWR VPWR _7975_/B sky130_fd_sc_hd__or2_1
XFILLER_94_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6925_ _6920_/Y _5902_/B _6921_/Y _5805_/B _6924_/X VGND VGND VPWR VPWR _6932_/C
+ sky130_fd_sc_hd__o221a_1
X_9713_ _9730_/CLK _9713_/D _9730_/SET_B VGND VGND VPWR VPWR _9713_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9644_ _9651_/CLK _9644_/D _9563_/SET_B VGND VGND VPWR VPWR _9644_/Q sky130_fd_sc_hd__dfrtp_1
X_6856_ _9537_/Q VGND VGND VPWR VPWR _6856_/Y sky130_fd_sc_hd__inv_4
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5807_ _5807_/A VGND VGND VPWR VPWR _5807_/Y sky130_fd_sc_hd__inv_2
X_9575_ _9576_/CLK _9575_/D _9571_/SET_B VGND VGND VPWR VPWR _9575_/Q sky130_fd_sc_hd__dfrtp_1
X_6787_ _9398_/Q VGND VGND VPWR VPWR _6787_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8526_ _8229_/B _8429_/A _8127_/B VGND VGND VPWR VPWR _8556_/C sky130_fd_sc_hd__o21ai_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5738_ _7477_/A VGND VGND VPWR VPWR _5738_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8457_ _8593_/A _8443_/B _8454_/X _8456_/Y VGND VGND VPWR VPWR _8457_/X sky130_fd_sc_hd__o211a_1
X_5669_ _9098_/Q VGND VGND VPWR VPWR _5669_/Y sky130_fd_sc_hd__inv_2
X_8388_ _8388_/A _8388_/B _8237_/X VGND VGND VPWR VPWR _8392_/C sky130_fd_sc_hd__or3b_1
XFILLER_163_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7408_ _6379_/Y _7139_/A _6440_/Y _7140_/A VGND VGND VPWR VPWR _7408_/X sky130_fd_sc_hd__o22a_1
Xhold450 hold450/A VGND VGND VPWR VPWR hold451/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold461 _9723_/Q VGND VGND VPWR VPWR hold462/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 hold472/A VGND VGND VPWR VPWR hold473/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7339_ _4940_/Y _7180_/X _4784_/Y _7181_/X _7338_/X VGND VGND VPWR VPWR _7340_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold494 _4937_/B VGND VGND VPWR VPWR hold495/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _4848_/X VGND VGND VPWR VPWR _5250_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_9009_ _7781_/X _9009_/A1 _9017_/S VGND VGND VPWR VPWR _9009_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4971_ _4971_/A VGND VGND VPWR VPWR _4971_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_189_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7690_ _6705_/Y _7519_/X _6742_/Y _7520_/X _7689_/X VGND VGND VPWR VPWR _7693_/C
+ sky130_fd_sc_hd__o221a_1
X_6710_ _6710_/A VGND VGND VPWR VPWR _6710_/Y sky130_fd_sc_hd__inv_4
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6641_ _9391_/Q VGND VGND VPWR VPWR _8807_/A sky130_fd_sc_hd__clkinv_8
XFILLER_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9360_ _9391_/CLK _9360_/D _9689_/SET_B VGND VGND VPWR VPWR _9360_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6572_ _7735_/A _5979_/B _6569_/Y _5201_/B _6571_/X VGND VGND VPWR VPWR _6572_/X
+ sky130_fd_sc_hd__o221a_1
X_8311_ _8311_/A _8621_/B VGND VGND VPWR VPWR _8313_/A sky130_fd_sc_hd__or2_1
XFILLER_185_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5523_ _5523_/A VGND VGND VPWR VPWR _5523_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9291_ _9297_/CLK _9291_/D _9797_/SET_B VGND VGND VPWR VPWR _9291_/Q sky130_fd_sc_hd__dfstp_1
X_8242_ _8419_/C VGND VGND VPWR VPWR _8382_/C sky130_fd_sc_hd__inv_2
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5454_ _9466_/Q _5446_/A hold601/A _5446_/Y VGND VGND VPWR VPWR _5454_/X sky130_fd_sc_hd__a22o_1
XFILLER_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5385_ _9513_/Q _5380_/A _6065_/B1 _5380_/Y VGND VGND VPWR VPWR _9513_/D sky130_fd_sc_hd__a22o_1
X_8173_ _8179_/A _8175_/A VGND VGND VPWR VPWR _8174_/A sky130_fd_sc_hd__or2_1
X_7124_ _4707_/Y _7171_/A _4899_/Y _7172_/A _7123_/X VGND VGND VPWR VPWR _7132_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7055_ _9288_/Q _9287_/Q _7118_/C _7092_/A VGND VGND VPWR VPWR _7056_/A sky130_fd_sc_hd__or4_4
X_6006_ _9137_/Q _6000_/A hold217/X _6000_/Y VGND VGND VPWR VPWR _9137_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7957_ _7957_/A _8296_/B VGND VGND VPWR VPWR _8534_/A sky130_fd_sc_hd__or2_1
X_7888_ _8421_/D _8421_/B _8436_/C _8236_/A VGND VGND VPWR VPWR _7953_/A sky130_fd_sc_hd__or4_4
XFILLER_23_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6908_ _6908_/A _6908_/B _6908_/C _6908_/D VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__and4_1
X_9627_ _9734_/CLK _9627_/D _9731_/SET_B VGND VGND VPWR VPWR _9627_/Q sky130_fd_sc_hd__dfrtp_1
X_6839_ _6839_/A VGND VGND VPWR VPWR _6839_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9558_ _9561_/CLK _9558_/D _9817_/SET_B VGND VGND VPWR VPWR _9558_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9489_ _9491_/CLK _9489_/D _9731_/SET_B VGND VGND VPWR VPWR _9489_/Q sky130_fd_sc_hd__dfrtp_1
X_8509_ _8509_/A VGND VGND VPWR VPWR _8672_/A sky130_fd_sc_hd__inv_2
XFILLER_40_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold280 hold280/A VGND VGND VPWR VPWR hold281/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 _6063_/X VGND VGND VPWR VPWR hold292/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_142 _8971_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _4923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_153 _5570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_164 _7907_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 _9814_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_197 _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5170_ _5170_/A VGND VGND VPWR VPWR _5170_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
X_8860_ _8860_/A VGND VGND VPWR VPWR _8860_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7811_ _7904_/D _7827_/B _8006_/A _8006_/C VGND VGND VPWR VPWR _7812_/A sky130_fd_sc_hd__or4_1
X_8791_ _8791_/A VGND VGND VPWR VPWR _8792_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7742_ _9125_/Q _9124_/Q _7743_/A VGND VGND VPWR VPWR _7742_/X sky130_fd_sc_hd__o21a_1
X_4954_ _4950_/Y _5482_/B _4952_/Y _5351_/B VGND VGND VPWR VPWR _4954_/X sky130_fd_sc_hd__o22a_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9412_ _9695_/CLK _9412_/D _9563_/SET_B VGND VGND VPWR VPWR _9412_/Q sky130_fd_sc_hd__dfrtp_1
X_7673_ _6843_/Y _7527_/X _6959_/Y _7528_/X VGND VGND VPWR VPWR _7673_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4885_ _4877_/Y _5340_/B _4879_/Y _4511_/B _4884_/X VGND VGND VPWR VPWR _4886_/D
+ sky130_fd_sc_hd__o221a_1
X_6624_ _6624_/A VGND VGND VPWR VPWR _6624_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_177_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9343_ _9421_/CLK _9343_/D _9537_/SET_B VGND VGND VPWR VPWR _9343_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6555_ _6553_/Y _5628_/B _8785_/A _5068_/B VGND VGND VPWR VPWR _6555_/X sky130_fd_sc_hd__o22a_1
X_9274_ _9392_/CLK _9274_/D _9537_/SET_B VGND VGND VPWR VPWR _9274_/Q sky130_fd_sc_hd__dfstp_1
X_5506_ _5506_/A VGND VGND VPWR VPWR _5507_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8225_ _8225_/A _8678_/B VGND VGND VPWR VPWR _8337_/A sky130_fd_sc_hd__or2_1
XFILLER_133_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6486_ _6486_/A VGND VGND VPWR VPWR _8850_/B sky130_fd_sc_hd__clkinv_4
XFILLER_105_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput341 _8865_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_2
Xoutput352 _9807_/Q VGND VGND VPWR VPWR sram_ro_addr[3] sky130_fd_sc_hd__buf_2
Xoutput330 _9781_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_2
X_5437_ _5437_/A VGND VGND VPWR VPWR _5437_/X sky130_fd_sc_hd__clkbuf_2
Xoutput374 _9076_/Q VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_2
X_5368_ _5368_/A VGND VGND VPWR VPWR _5369_/A sky130_fd_sc_hd__clkbuf_4
Xoutput363 _9058_/Q VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput385 _9065_/Q VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_2
X_8156_ _8443_/A VGND VGND VPWR VPWR _8156_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_59_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5299_ _9571_/Q _5292_/A _6067_/B1 _5292_/Y VGND VGND VPWR VPWR _9571_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8087_ _8666_/B _8596_/A VGND VGND VPWR VPWR _8509_/A sky130_fd_sc_hd__or2_1
X_7107_ _7129_/C _7107_/B VGND VGND VPWR VPWR _7151_/A sky130_fd_sc_hd__or2_2
XFILLER_101_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7038_ _4974_/Y _4975_/Y _6054_/Y _9093_/Q _7039_/A VGND VGND VPWR VPWR _9093_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_47_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8989_ _8988_/X hold415/X _9629_/Q VGND VGND VPWR VPWR _8989_/X sky130_fd_sc_hd__mux2_4
XFILLER_82_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4670_ _9756_/Q _4657_/A _8995_/X _4657_/Y VGND VGND VPWR VPWR _9756_/D sky130_fd_sc_hd__a22o_1
X_6340_ _9303_/Q VGND VGND VPWR VPWR _6340_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6271_ _9549_/Q VGND VGND VPWR VPWR _6271_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_115_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8010_ _8010_/A VGND VGND VPWR VPWR _8139_/A sky130_fd_sc_hd__buf_4
XFILLER_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5222_ _9622_/Q _5216_/Y _8961_/X _5216_/A VGND VGND VPWR VPWR _9622_/D sky130_fd_sc_hd__o22a_1
X_5153_ _5153_/A VGND VGND VPWR VPWR _5153_/X sky130_fd_sc_hd__clkbuf_1
X_5084_ _8854_/A _5081_/X _8853_/A _5083_/X VGND VGND VPWR VPWR _5085_/C sky130_fd_sc_hd__o22ai_1
XFILLER_110_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8912_ _8911_/X hold707/X _9096_/Q VGND VGND VPWR VPWR _8912_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8843_ _8843_/A _8843_/B VGND VGND VPWR VPWR _8844_/A sky130_fd_sc_hd__and2_1
XFILLER_52_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5986_ _9151_/Q _5981_/A _8964_/A1 _5981_/Y VGND VGND VPWR VPWR _9151_/D sky130_fd_sc_hd__a22o_1
X_8774_ _8774_/A VGND VGND VPWR VPWR _8774_/Y sky130_fd_sc_hd__inv_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4937_ _6117_/B _4937_/B VGND VGND VPWR VPWR _4937_/X sky130_fd_sc_hd__or2_4
X_7725_ _6400_/Y _7521_/A _6428_/Y _7522_/A VGND VGND VPWR VPWR _7725_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_20 _6127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _9570_/Q VGND VGND VPWR VPWR _4868_/Y sky130_fd_sc_hd__clkinv_4
X_7656_ _4719_/Y _7525_/X _7336_/A _7526_/X _7655_/X VGND VGND VPWR VPWR _7657_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA_31 _6287_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6607_ _9573_/Q VGND VGND VPWR VPWR _8821_/A sky130_fd_sc_hd__clkinv_8
XANTENNA_53 _6875_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 _6434_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _7050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7587_ _6321_/Y _7487_/X _6334_/Y _7488_/X VGND VGND VPWR VPWR _7587_/X sky130_fd_sc_hd__o22a_1
X_9326_ _9326_/CLK _9326_/D _9571_/SET_B VGND VGND VPWR VPWR _9326_/Q sky130_fd_sc_hd__dfrtp_1
X_4799_ _4790_/Y _5112_/B _4792_/Y _5609_/B _4798_/X VGND VGND VPWR VPWR _4811_/C
+ sky130_fd_sc_hd__o221a_1
XANTENNA_86 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6538_ _8797_/A _5786_/B _6534_/Y _5513_/B _6537_/X VGND VGND VPWR VPWR _6557_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9257_ _9673_/CLK _9257_/D _9730_/SET_B VGND VGND VPWR VPWR _9257_/Q sky130_fd_sc_hd__dfrtp_1
X_6469_ _6469_/A VGND VGND VPWR VPWR _6469_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8208_ _8208_/A _8757_/A VGND VGND VPWR VPWR _8213_/A sky130_fd_sc_hd__or2_1
XFILLER_79_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9188_ _9322_/CLK _9188_/D _9797_/SET_B VGND VGND VPWR VPWR _9188_/Q sky130_fd_sc_hd__dfrtp_1
X_8139_ _8139_/A _8139_/B VGND VGND VPWR VPWR _8730_/A sky130_fd_sc_hd__nor2_1
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5840_ _5840_/A VGND VGND VPWR VPWR _5841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5771_ _5990_/A _5771_/B VGND VGND VPWR VPWR _5772_/A sky130_fd_sc_hd__or2_1
X_8490_ _8654_/A _8490_/B _8490_/C _8489_/X VGND VGND VPWR VPWR _8491_/B sky130_fd_sc_hd__or4b_1
X_4722_ _4915_/B _4806_/B VGND VGND VPWR VPWR _5036_/B sky130_fd_sc_hd__or2_4
X_7510_ _7510_/A VGND VGND VPWR VPWR _7510_/X sky130_fd_sc_hd__buf_4
XFILLER_187_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7441_ _7441_/A _9295_/Q VGND VGND VPWR VPWR _7478_/C sky130_fd_sc_hd__or2_2
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR _6348_/A sky130_fd_sc_hd__clkbuf_1
X_4653_ _9739_/Q VGND VGND VPWR VPWR _5237_/A sky130_fd_sc_hd__inv_2
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__buf_2
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4584_ _4913_/A _4643_/A VGND VGND VPWR VPWR _4585_/B sky130_fd_sc_hd__or2_4
X_7372_ _6738_/Y _7155_/X _6750_/Y _7156_/X _7371_/X VGND VGND VPWR VPWR _7375_/C
+ sky130_fd_sc_hd__o221a_1
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _7049_/B sky130_fd_sc_hd__clkbuf_1
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_4
XFILLER_115_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9111_ _9832_/CLK _9111_/D _9821_/SET_B VGND VGND VPWR VPWR _9111_/Q sky130_fd_sc_hd__dfrtp_4
Xinput95 sram_ro_data[11] VGND VGND VPWR VPWR _6583_/A sky130_fd_sc_hd__clkbuf_1
X_6323_ _6323_/A VGND VGND VPWR VPWR _6323_/Y sky130_fd_sc_hd__inv_2
X_9042_ _9610_/Q _8819_/A VGND VGND VPWR VPWR _9042_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_170_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6254_ _6249_/Y _5979_/B _6250_/Y _4863_/X _6253_/X VGND VGND VPWR VPWR _6267_/B
+ sky130_fd_sc_hd__o221a_1
X_5205_ _9634_/Q _5203_/A hold53/X _5203_/Y VGND VGND VPWR VPWR _9634_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6185_ _9394_/Q VGND VGND VPWR VPWR _6185_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5136_ _9681_/Q _5135_/A hold516/X _5135_/Y VGND VGND VPWR VPWR _9681_/D sky130_fd_sc_hd__a22o_1
X_5067_ _9011_/X _4572_/B _9717_/Q _5085_/D VGND VGND VPWR VPWR _9717_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8826_ _8826_/A VGND VGND VPWR VPWR _8826_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5969_ _5969_/A _5969_/B VGND VGND VPWR VPWR _5969_/X sky130_fd_sc_hd__or2_1
X_8757_ _8757_/A _8757_/B _8757_/C VGND VGND VPWR VPWR _8758_/B sky130_fd_sc_hd__or3_1
X_7708_ _6517_/Y _7519_/A _6581_/Y _7520_/A _7707_/X VGND VGND VPWR VPWR _7711_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8688_ _8688_/A _8688_/B VGND VGND VPWR VPWR _8720_/C sky130_fd_sc_hd__or2_1
XFILLER_32_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7639_ _7639_/A _7639_/B _7639_/C _7639_/D VGND VGND VPWR VPWR _7640_/D sky130_fd_sc_hd__and4_1
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9309_ _9831_/CLK _9309_/D _9727_/SET_B VGND VGND VPWR VPWR _9309_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold109 hold109/A VGND VGND VPWR VPWR hold110/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7990_ _8436_/D _8557_/B _8702_/C VGND VGND VPWR VPWR _8228_/A sky130_fd_sc_hd__or3_1
X_6941_ _9710_/Q VGND VGND VPWR VPWR _6941_/Y sky130_fd_sc_hd__inv_2
X_9660_ _9734_/CLK _9660_/D _9731_/SET_B VGND VGND VPWR VPWR _9660_/Q sky130_fd_sc_hd__dfrtp_1
X_6872_ _6870_/Y _4579_/B _6871_/Y _5474_/B VGND VGND VPWR VPWR _6872_/X sky130_fd_sc_hd__o22a_1
X_8611_ _8682_/A _8610_/X _8265_/A _8394_/C VGND VGND VPWR VPWR _8761_/A sky130_fd_sc_hd__o211ai_2
X_9591_ _9832_/CLK _9591_/D _9797_/SET_B VGND VGND VPWR VPWR _9591_/Q sky130_fd_sc_hd__dfrtp_4
X_5823_ _9256_/Q _5820_/A _8965_/A1 _5820_/Y VGND VGND VPWR VPWR _9256_/D sky130_fd_sc_hd__a22o_1
X_8542_ _8737_/A _8701_/A _8636_/B _7931_/X VGND VGND VPWR VPWR _8543_/D sky130_fd_sc_hd__or4b_1
XFILLER_34_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5754_ _7129_/C VGND VGND VPWR VPWR _7127_/A sky130_fd_sc_hd__buf_2
XFILLER_175_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8473_ _8473_/A _8473_/B VGND VGND VPWR VPWR _8474_/C sky130_fd_sc_hd__or2_1
XFILLER_147_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4705_ _9240_/Q VGND VGND VPWR VPWR _4705_/Y sky130_fd_sc_hd__inv_2
X_5685_ _5685_/A VGND VGND VPWR VPWR _5685_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7424_ _7424_/A _7424_/B VGND VGND VPWR VPWR _7424_/X sky130_fd_sc_hd__or2_1
X_4636_ _4636_/A VGND VGND VPWR VPWR _4636_/Y sky130_fd_sc_hd__inv_2
Xhold610 _5200_/X VGND VGND VPWR VPWR _9636_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_190_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold621 _5290_/X VGND VGND VPWR VPWR _5291_/A sky130_fd_sc_hd__clkdlybuf4s25_1
X_7355_ _6940_/Y _7071_/D _6929_/Y _7166_/X _7354_/X VGND VGND VPWR VPWR _7362_/A
+ sky130_fd_sc_hd__o221a_1
X_4567_ _9110_/Q VGND VGND VPWR VPWR _8855_/A sky130_fd_sc_hd__inv_2
Xhold632 _5495_/A VGND VGND VPWR VPWR hold632/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6306_ _9575_/Q VGND VGND VPWR VPWR _6306_/Y sky130_fd_sc_hd__clkinv_2
Xhold654 _5054_/X VGND VGND VPWR VPWR _9725_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold643 _4603_/X VGND VGND VPWR VPWR _9787_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7286_ _6215_/Y _7160_/X _6188_/Y _7071_/B _7285_/X VGND VGND VPWR VPWR _7287_/D
+ sky130_fd_sc_hd__o221a_1
Xhold676 _5907_/X VGND VGND VPWR VPWR _9198_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_4498_ _4498_/A VGND VGND VPWR VPWR _4498_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold665 _6165_/A VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__buf_2
Xhold687 _4883_/A VGND VGND VPWR VPWR _4482_/A sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_170_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9025_ _9025_/A _7733_/A VGND VGND VPWR VPWR _9025_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6237_ input9/X VGND VGND VPWR VPWR _6237_/Y sky130_fd_sc_hd__inv_2
Xhold698 _9752_/Q VGND VGND VPWR VPWR hold698/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6168_ _6163_/Y _6353_/A _6164_/Y _5570_/B _6167_/Y VGND VGND VPWR VPWR _6175_/C
+ sky130_fd_sc_hd__o221a_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _9691_/Q _5114_/A hold42/X _5114_/Y VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__a22o_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6099_ _9413_/Q VGND VGND VPWR VPWR _6099_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _9297_/CLK sky130_fd_sc_hd__clkbuf_2
X_8809_ _8809_/A VGND VGND VPWR VPWR _8810_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_43_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9789_ _9791_/CLK _9789_/D _9821_/SET_B VGND VGND VPWR VPWR _9789_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_159_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5470_ _9456_/Q _5468_/A _6065_/B1 _5468_/Y VGND VGND VPWR VPWR _9456_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7140_ _7140_/A VGND VGND VPWR VPWR _7140_/X sky130_fd_sc_hd__buf_4
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7071_ _7071_/A _7071_/B _7071_/C _7071_/D VGND VGND VPWR VPWR _7095_/C sky130_fd_sc_hd__and4_1
XFILLER_98_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6022_ _6022_/A VGND VGND VPWR VPWR _6022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7973_ _8324_/C _7873_/C _7868_/Y _7972_/X VGND VGND VPWR VPWR _7974_/B sky130_fd_sc_hd__a31o_1
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9712_ _9731_/CLK _9712_/D _9731_/SET_B VGND VGND VPWR VPWR _9712_/Q sky130_fd_sc_hd__dfrtp_2
X_6924_ _6922_/Y _5706_/B _6923_/Y _5513_/B VGND VGND VPWR VPWR _6924_/X sky130_fd_sc_hd__o22a_1
X_9643_ _9643_/CLK _9643_/D _9689_/SET_B VGND VGND VPWR VPWR _9643_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6855_ _9527_/Q VGND VGND VPWR VPWR _6855_/Y sky130_fd_sc_hd__clkinv_2
X_5806_ _5806_/A VGND VGND VPWR VPWR _5807_/A sky130_fd_sc_hd__clkbuf_4
X_6786_ _9195_/Q VGND VGND VPWR VPWR _6786_/Y sky130_fd_sc_hd__clkinv_2
X_9574_ _9574_/CLK _9574_/D _9571_/SET_B VGND VGND VPWR VPWR _9574_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8525_ _8525_/A _8647_/A VGND VGND VPWR VPWR _8527_/A sky130_fd_sc_hd__or2_1
X_5737_ _7479_/A _7432_/B VGND VGND VPWR VPWR _7477_/A sky130_fd_sc_hd__or2_4
XFILLER_148_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8456_ _8669_/C VGND VGND VPWR VPWR _8456_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5668_ _9096_/Q VGND VGND VPWR VPWR _7028_/A sky130_fd_sc_hd__clkinv_2
X_7407_ _7407_/A _7407_/B _7407_/C VGND VGND VPWR VPWR _7407_/Y sky130_fd_sc_hd__nand3_1
X_8387_ _8387_/A _8387_/B VGND VGND VPWR VPWR _8419_/B sky130_fd_sc_hd__or2_1
X_5599_ _5599_/A VGND VGND VPWR VPWR _5600_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4619_ _9776_/Q _4613_/A hold217/X _4613_/Y VGND VGND VPWR VPWR _9776_/D sky130_fd_sc_hd__a22o_1
XFILLER_150_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold451 hold451/A VGND VGND VPWR VPWR _5446_/A sky130_fd_sc_hd__clkbuf_4
Xhold440 hold440/A VGND VGND VPWR VPWR _9116_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold462 hold462/A VGND VGND VPWR VPWR hold463/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7338_ _4904_/Y _7182_/X _4831_/Y _7183_/X VGND VGND VPWR VPWR _7338_/X sky130_fd_sc_hd__o22a_1
X_7269_ _6346_/Y _7171_/X _6307_/Y _7172_/X _7268_/X VGND VGND VPWR VPWR _7274_/B
+ sky130_fd_sc_hd__o221a_1
Xhold484 _4848_/B VGND VGND VPWR VPWR _4949_/A sky130_fd_sc_hd__clkbuf_2
Xhold473 hold473/A VGND VGND VPWR VPWR _4685_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xhold495 hold495/A VGND VGND VPWR VPWR hold496/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9008_ _7779_/X _9008_/A1 _9017_/S VGND VGND VPWR VPWR _9008_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4970_ _4970_/A VGND VGND VPWR VPWR _4970_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6640_ _9586_/Q VGND VGND VPWR VPWR _6640_/Y sky130_fd_sc_hd__clkinv_4
X_6571_ hold23/A _8973_/S _6570_/Y _5971_/B VGND VGND VPWR VPWR _6571_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_192_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5522_ _5522_/A VGND VGND VPWR VPWR _5523_/A sky130_fd_sc_hd__buf_4
X_8310_ _8702_/A _8312_/B VGND VGND VPWR VPWR _8621_/B sky130_fd_sc_hd__nor2_1
XFILLER_157_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9290_ _9297_/CLK _9290_/D _9797_/SET_B VGND VGND VPWR VPWR _9290_/Q sky130_fd_sc_hd__dfrtp_2
X_8241_ _8260_/A _8241_/B _8241_/C VGND VGND VPWR VPWR _8419_/C sky130_fd_sc_hd__or3_2
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5453_ _9467_/Q _5446_/A _6067_/B1 _5446_/Y VGND VGND VPWR VPWR _5453_/X sky130_fd_sc_hd__a22o_1
X_5384_ _9514_/Q _5380_/A _6064_/B1 _5380_/Y VGND VGND VPWR VPWR _9514_/D sky130_fd_sc_hd__a22o_1
X_8172_ _8172_/A _8718_/A _8399_/A _8615_/A VGND VGND VPWR VPWR _8177_/A sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_42_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9798_/CLK sky130_fd_sc_hd__clkbuf_16
X_7123_ _4868_/Y _7173_/A _4695_/Y _7174_/A VGND VGND VPWR VPWR _7123_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7054_ _9290_/Q _9289_/Q VGND VGND VPWR VPWR _7118_/C sky130_fd_sc_hd__or2_2
X_6005_ _9138_/Q _5999_/X _6065_/B1 _6000_/Y VGND VGND VPWR VPWR _6005_/X sky130_fd_sc_hd__a22o_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7956_ _8776_/A _7956_/B _8359_/A _8639_/A VGND VGND VPWR VPWR _7956_/Y sky130_fd_sc_hd__nor4_1
X_7887_ _7887_/A _8118_/A VGND VGND VPWR VPWR _7968_/A sky130_fd_sc_hd__or2_1
X_6907_ _6902_/Y _5482_/B _6903_/Y _5505_/B _6906_/X VGND VGND VPWR VPWR _6908_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_168_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6838_ _9828_/Q VGND VGND VPWR VPWR _6838_/Y sky130_fd_sc_hd__inv_4
X_9626_ _9734_/CLK _9626_/D _9731_/SET_B VGND VGND VPWR VPWR _9626_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9557_ _9686_/CLK _9557_/D _9817_/SET_B VGND VGND VPWR VPWR _9557_/Q sky130_fd_sc_hd__dfrtp_1
X_6769_ _9356_/Q VGND VGND VPWR VPWR _6769_/Y sky130_fd_sc_hd__inv_2
X_8508_ _8508_/A _8657_/C VGND VGND VPWR VPWR _8512_/A sky130_fd_sc_hd__or2_1
XFILLER_176_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9488_ _9491_/CLK _9488_/D _9731_/SET_B VGND VGND VPWR VPWR _9488_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8439_ _8439_/A _8439_/B VGND VGND VPWR VPWR _8439_/Y sky130_fd_sc_hd__nor2_1
XFILLER_191_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold270 _5652_/X VGND VGND VPWR VPWR hold271/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 hold281/A VGND VGND VPWR VPWR _9649_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold292 hold292/A VGND VGND VPWR VPWR hold293/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _7604_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_110 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 _8858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_154 _8849_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _7912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_176 _8843_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_187 _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7810_ _8234_/A _7810_/B _7810_/C _7810_/D VGND VGND VPWR VPWR _8006_/C sky130_fd_sc_hd__or4_1
X_8790_ _8790_/A VGND VGND VPWR VPWR _8790_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7741_ _9125_/Q _9124_/Q VGND VGND VPWR VPWR _7743_/A sky130_fd_sc_hd__nand2_1
X_4953_ _4953_/A _4953_/B VGND VGND VPWR VPWR _5351_/B sky130_fd_sc_hd__or2_4
X_7672_ _6940_/Y _7519_/X _6876_/Y _7520_/X _7671_/X VGND VGND VPWR VPWR _7675_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9411_ _9695_/CLK _9411_/D _9563_/SET_B VGND VGND VPWR VPWR _9411_/Q sky130_fd_sc_hd__dfrtp_1
X_6623_ input6/X VGND VGND VPWR VPWR _6623_/Y sky130_fd_sc_hd__inv_2
X_4884_ _4880_/Y _5397_/B _4882_/Y _4883_/X VGND VGND VPWR VPWR _4884_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9342_ _9421_/CLK _9342_/D _9563_/SET_B VGND VGND VPWR VPWR _9342_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_158_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6554_ _9712_/Q VGND VGND VPWR VPWR _8785_/A sky130_fd_sc_hd__inv_6
XFILLER_20_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9273_ _9392_/CLK _9273_/D _9563_/SET_B VGND VGND VPWR VPWR _9273_/Q sky130_fd_sc_hd__dfstp_1
X_6485_ _6480_/Y _4611_/B _6481_/Y _6166_/A _6484_/X VGND VGND VPWR VPWR _6504_/A
+ sky130_fd_sc_hd__o221a_1
X_5505_ _5698_/A _5505_/B VGND VGND VPWR VPWR _5506_/A sky130_fd_sc_hd__or2_1
X_8224_ _8137_/A _8428_/A _8138_/B _9108_/Q VGND VGND VPWR VPWR _8678_/B sky130_fd_sc_hd__o31ai_4
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5436_ _5474_/A _5436_/B VGND VGND VPWR VPWR _5437_/A sky130_fd_sc_hd__or2_1
XFILLER_145_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput353 _9808_/Q VGND VGND VPWR VPWR sram_ro_addr[4] sky130_fd_sc_hd__buf_2
Xoutput342 _8862_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_2
Xoutput331 _9782_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_2
Xoutput320 _9795_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_2
Xoutput375 _9077_/Q VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_2
X_5367_ _5378_/A _5367_/B VGND VGND VPWR VPWR _5368_/A sky130_fd_sc_hd__or2_1
Xoutput364 _9059_/Q VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_2
XFILLER_120_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput386 _9066_/Q VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_2
X_8155_ _8179_/A VGND VGND VPWR VPWR _8155_/Y sky130_fd_sc_hd__inv_2
X_5298_ _9572_/Q _5292_/A hold217/X _5292_/Y VGND VGND VPWR VPWR _5298_/X sky130_fd_sc_hd__a22o_1
X_8086_ _8086_/A _8657_/B VGND VGND VPWR VPWR _8088_/A sky130_fd_sc_hd__nor2_1
X_7106_ _7127_/A _7106_/B VGND VGND VPWR VPWR _7149_/A sky130_fd_sc_hd__or2_2
XFILLER_101_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7037_ _9750_/Q _6024_/B _9090_/Q _9094_/Q VGND VGND VPWR VPWR _9094_/D sky130_fd_sc_hd__a31o_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8988_ hold672/X hold619/X _9093_/Q VGND VGND VPWR VPWR _8988_/X sky130_fd_sc_hd__mux2_2
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ _7939_/A _8570_/B VGND VGND VPWR VPWR _8559_/A sky130_fd_sc_hd__or2b_2
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9609_ _9651_/CLK _9609_/D _9689_/SET_B VGND VGND VPWR VPWR _9609_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6270_ _9471_/Q VGND VGND VPWR VPWR _6270_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5221_ _9623_/Q _5216_/Y _8943_/X _5216_/A VGND VGND VPWR VPWR _9623_/D sky130_fd_sc_hd__o22a_1
XFILLER_102_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5152_ _6017_/A VGND VGND VPWR VPWR _5153_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5083_ _5083_/A VGND VGND VPWR VPWR _5083_/X sky130_fd_sc_hd__clkbuf_1
X_8911_ _7712_/Y _9672_/Q _9020_/S VGND VGND VPWR VPWR _8911_/X sky130_fd_sc_hd__mux2_1
X_8842_ _8842_/A VGND VGND VPWR VPWR _8842_/X sky130_fd_sc_hd__clkbuf_1
X_8773_ _8773_/A _8773_/B _8773_/C _8773_/D VGND VGND VPWR VPWR _8773_/X sky130_fd_sc_hd__or4_1
X_5985_ _9152_/Q _5981_/A _8959_/A1 _5981_/Y VGND VGND VPWR VPWR _9152_/D sky130_fd_sc_hd__a22o_1
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7724_ _6498_/Y _7513_/A _6379_/Y _7514_/A _7723_/X VGND VGND VPWR VPWR _7729_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4936_ _9466_/Q VGND VGND VPWR VPWR _4936_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_21 _6125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7655_ _4904_/Y _7527_/X _4726_/Y _7528_/X VGND VGND VPWR VPWR _7655_/X sky130_fd_sc_hd__o22a_1
X_4867_ _4862_/Y _4863_/X _4864_/Y _4865_/X _4866_/X VGND VGND VPWR VPWR _4886_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA_32 _6302_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 _4889_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6606_ _9417_/Q VGND VGND VPWR VPWR _8809_/A sky130_fd_sc_hd__inv_6
X_7586_ _7586_/A _7586_/B _7586_/C _7586_/D VGND VGND VPWR VPWR _7586_/Y sky130_fd_sc_hd__nand4_2
XANTENNA_43 _6534_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 _7050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _6878_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9325_ _9326_/CLK _9325_/D _9571_/SET_B VGND VGND VPWR VPWR _9325_/Q sky130_fd_sc_hd__dfstp_1
X_4798_ _4794_/Y _5068_/B _4796_/Y _5946_/B VGND VGND VPWR VPWR _4798_/X sky130_fd_sc_hd__o22a_1
X_6537_ _6535_/Y _5858_/B _6536_/Y _6165_/A VGND VGND VPWR VPWR _6537_/X sky130_fd_sc_hd__o22a_1
XANTENNA_87 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6468_ _6466_/Y _5133_/B _6467_/Y _5532_/B VGND VGND VPWR VPWR _6468_/X sky130_fd_sc_hd__o22a_1
X_9256_ _9833_/CLK _9256_/D _9730_/SET_B VGND VGND VPWR VPWR _9256_/Q sky130_fd_sc_hd__dfstp_1
X_6399_ _9277_/Q VGND VGND VPWR VPWR _6399_/Y sky130_fd_sc_hd__inv_2
X_5419_ _5419_/A VGND VGND VPWR VPWR _5419_/Y sky130_fd_sc_hd__inv_2
X_8207_ _8209_/A _8682_/B VGND VGND VPWR VPWR _8757_/A sky130_fd_sc_hd__nor2_1
X_9187_ _9319_/CLK _9187_/D _9797_/SET_B VGND VGND VPWR VPWR _9187_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8138_ _8211_/A _8138_/B VGND VGND VPWR VPWR _8139_/B sky130_fd_sc_hd__or2_1
XFILLER_102_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8069_ _8563_/A _8592_/A VGND VGND VPWR VPWR _8452_/A sky130_fd_sc_hd__or2_1
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _5770_/A VGND VGND VPWR VPWR _5990_/A sky130_fd_sc_hd__buf_6
XFILLER_175_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4721_ _9730_/Q VGND VGND VPWR VPWR _4721_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7440_ _4899_/Y _7485_/A _4741_/Y _7486_/A _7439_/X VGND VGND VPWR VPWR _7483_/A
+ sky130_fd_sc_hd__o221a_1
X_4652_ _6081_/A VGND VGND VPWR VPWR _4969_/A sky130_fd_sc_hd__clkbuf_4
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR _6501_/A sky130_fd_sc_hd__clkbuf_1
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _8845_/A sky130_fd_sc_hd__buf_6
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR _4802_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_190_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9110_ _4471_/A1 _9110_/D _6177_/A VGND VGND VPWR VPWR _9110_/Q sky130_fd_sc_hd__dfrtp_4
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_2
X_7371_ _6688_/Y _7056_/A _6665_/Y _7157_/X VGND VGND VPWR VPWR _7371_/X sky130_fd_sc_hd__o22a_1
X_4583_ _4583_/A VGND VGND VPWR VPWR _9798_/D sky130_fd_sc_hd__clkbuf_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_4
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6322_ _9117_/Q VGND VGND VPWR VPWR _6322_/Y sky130_fd_sc_hd__inv_2
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _7051_/B sky130_fd_sc_hd__clkbuf_2
Xinput96 sram_ro_data[12] VGND VGND VPWR VPWR _6367_/A sky130_fd_sc_hd__clkbuf_1
X_9041_ _9609_/Q _8817_/A VGND VGND VPWR VPWR _9041_/Z sky130_fd_sc_hd__ebufn_1
X_6253_ _6251_/Y _4585_/B _6252_/Y _4915_/X VGND VGND VPWR VPWR _6253_/X sky130_fd_sc_hd__o22a_1
X_5204_ _9635_/Q _5203_/A hold577/A _5203_/Y VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6184_ _6184_/A VGND VGND VPWR VPWR _6184_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5135_ _5135_/A VGND VGND VPWR VPWR _5135_/Y sky130_fd_sc_hd__inv_2
X_5066_ _9012_/X _4572_/B _9718_/Q _5085_/D VGND VGND VPWR VPWR _9718_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8825_ _8825_/A VGND VGND VPWR VPWR _8826_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5968_ _6178_/B _7032_/B VGND VGND VPWR VPWR _5968_/Y sky130_fd_sc_hd__nor2_1
X_8756_ _8756_/A _8756_/B _8756_/C _8756_/D VGND VGND VPWR VPWR _8781_/A sky130_fd_sc_hd__or4_1
XFILLER_80_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4919_ _9518_/Q VGND VGND VPWR VPWR _4919_/Y sky130_fd_sc_hd__inv_6
X_7707_ _6529_/Y _7521_/A _6605_/Y _7522_/A VGND VGND VPWR VPWR _7707_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5899_ _9203_/Q _5896_/A hold217/X _5896_/Y VGND VGND VPWR VPWR _9203_/D sky130_fd_sc_hd__a22o_1
X_8687_ _8687_/A _8687_/B _8687_/C _8687_/D VGND VGND VPWR VPWR _8758_/C sky130_fd_sc_hd__or4_4
X_7638_ _6159_/Y _7525_/X _7314_/A _7526_/X _7637_/X VGND VGND VPWR VPWR _7639_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7569_ _6427_/Y _7487_/X _6365_/Y _7488_/X VGND VGND VPWR VPWR _7569_/X sky130_fd_sc_hd__o22a_1
X_9308_ _9831_/CLK _9308_/D _9727_/SET_B VGND VGND VPWR VPWR _9308_/Q sky130_fd_sc_hd__dfstp_1
X_9239_ _9421_/CLK _9239_/D _9537_/SET_B VGND VGND VPWR VPWR _9239_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6940_ _9202_/Q VGND VGND VPWR VPWR _6940_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6871_ _9449_/Q VGND VGND VPWR VPWR _6871_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8610_ _8243_/B _8682_/C _8257_/X VGND VGND VPWR VPWR _8610_/X sky130_fd_sc_hd__o21a_1
X_9590_ _9832_/CLK _9590_/D _9797_/SET_B VGND VGND VPWR VPWR _9590_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5822_ _9257_/Q _5820_/A _8964_/A1 _5820_/Y VGND VGND VPWR VPWR _9257_/D sky130_fd_sc_hd__a22o_1
X_8541_ _8613_/B _8541_/B VGND VGND VPWR VPWR _8701_/A sky130_fd_sc_hd__or2_1
X_5753_ _9292_/Q _5753_/B VGND VGND VPWR VPWR _7129_/C sky130_fd_sc_hd__or2_2
XFILLER_147_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4704_ _4695_/Y _5532_/B _4697_/Y _5103_/B _4703_/X VGND VGND VPWR VPWR _4725_/B
+ sky130_fd_sc_hd__o221a_1
X_8472_ _8472_/A _8602_/B VGND VGND VPWR VPWR _8473_/B sky130_fd_sc_hd__or2_1
X_5684_ _9096_/Q _9098_/Q _5723_/A _5673_/X _5683_/Y VGND VGND VPWR VPWR _9320_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4635_ _4635_/A VGND VGND VPWR VPWR _4636_/A sky130_fd_sc_hd__clkbuf_2
X_7423_ _6489_/Y _7171_/A _6455_/Y _7172_/A _7422_/X VGND VGND VPWR VPWR _7428_/B
+ sky130_fd_sc_hd__o221a_1
Xhold611 _9704_/Q VGND VGND VPWR VPWR hold611/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_4566_ _9109_/Q VGND VGND VPWR VPWR _8854_/A sky130_fd_sc_hd__inv_2
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold600 _5420_/X VGND VGND VPWR VPWR _9491_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7354_ _6969_/Y _7167_/X _6927_/Y _7168_/X VGND VGND VPWR VPWR _7354_/X sky130_fd_sc_hd__o22a_1
XFILLER_190_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6305_ _9497_/Q VGND VGND VPWR VPWR _6305_/Y sky130_fd_sc_hd__clkinv_4
Xhold633 _5499_/X VGND VGND VPWR VPWR _9436_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold644 _5832_/X VGND VGND VPWR VPWR _9250_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold622 _4869_/A VGND VGND VPWR VPWR _4898_/B sky130_fd_sc_hd__buf_2
Xhold688 _5245_/X VGND VGND VPWR VPWR _9607_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7285_ _6213_/Y _7161_/X _6230_/Y _7162_/X VGND VGND VPWR VPWR _7285_/X sky130_fd_sc_hd__o22a_1
Xhold666 _5226_/A VGND VGND VPWR VPWR hold666/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4497_ _6008_/B1 _9831_/Q _4497_/S VGND VGND VPWR VPWR _4497_/X sky130_fd_sc_hd__mux2_1
X_9024_ _9625_/Q _8787_/A VGND VGND VPWR VPWR _9024_/Z sky130_fd_sc_hd__ebufn_1
Xhold655 _5443_/X VGND VGND VPWR VPWR _9474_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold677 _5151_/X VGND VGND VPWR VPWR _9669_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold699 _7020_/Y VGND VGND VPWR VPWR _9110_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6236_ _9412_/Q VGND VGND VPWR VPWR _6236_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6167_ input42/X _8971_/S input51/X _8975_/S VGND VGND VPWR VPWR _6167_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_134_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _9692_/Q _5114_/A hold53/X _5114_/Y VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__a22o_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ _9335_/Q VGND VGND VPWR VPWR _6098_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5049_ _5049_/A VGND VGND VPWR VPWR _5049_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8808_ _8808_/A VGND VGND VPWR VPWR _8808_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9788_ _9791_/CLK _9788_/D _9817_/SET_B VGND VGND VPWR VPWR _9788_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_185_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8739_ _8739_/A VGND VGND VPWR VPWR _8739_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7070_ _7070_/A VGND VGND VPWR VPWR _7071_/D sky130_fd_sc_hd__buf_4
X_6021_ _6071_/A VGND VGND VPWR VPWR _6022_/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7972_ _8704_/A _7972_/B VGND VGND VPWR VPWR _7972_/X sky130_fd_sc_hd__or2_1
XFILLER_66_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6923_ _9423_/Q VGND VGND VPWR VPWR _6923_/Y sky130_fd_sc_hd__clkinv_2
X_9711_ _9734_/CLK _9711_/D _9731_/SET_B VGND VGND VPWR VPWR _9711_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9642_ _9643_/CLK _9642_/D _9689_/SET_B VGND VGND VPWR VPWR _9642_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6854_ _9113_/Q VGND VGND VPWR VPWR _6854_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5805_ _5847_/A _5805_/B VGND VGND VPWR VPWR _5806_/A sky130_fd_sc_hd__or2_1
X_9573_ _9574_/CLK _9573_/D _9571_/SET_B VGND VGND VPWR VPWR _9573_/Q sky130_fd_sc_hd__dfrtp_4
X_6785_ _9169_/Q VGND VGND VPWR VPWR _6785_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8524_ _8604_/A _8692_/B VGND VGND VPWR VPWR _8647_/A sky130_fd_sc_hd__or2_1
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5736_ _9293_/Q VGND VGND VPWR VPWR _7432_/B sky130_fd_sc_hd__inv_2
X_8455_ _8656_/B _8617_/A VGND VGND VPWR VPWR _8669_/C sky130_fd_sc_hd__or2_1
X_5667_ _9319_/Q VGND VGND VPWR VPWR _5673_/A sky130_fd_sc_hd__inv_2
XFILLER_163_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4618_ _9777_/Q _4613_/A _6065_/B1 _4613_/Y VGND VGND VPWR VPWR _9777_/D sky130_fd_sc_hd__a22o_1
X_7406_ _7406_/A _7406_/B _7406_/C _7406_/D VGND VGND VPWR VPWR _7407_/C sky130_fd_sc_hd__and4_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8386_ _8321_/A _8420_/B _8682_/A _8321_/C _8353_/B VGND VGND VPWR VPWR _8394_/A
+ sky130_fd_sc_hd__o32a_1
X_5598_ _5847_/A _5598_/B VGND VGND VPWR VPWR _5599_/A sky130_fd_sc_hd__or2_1
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold441 _6059_/X VGND VGND VPWR VPWR hold442/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 _5444_/X VGND VGND VPWR VPWR _5445_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold430 _6005_/X VGND VGND VPWR VPWR hold431/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 hold463/A VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_7337_ _4880_/Y _5756_/X _4712_/A _7071_/A _7336_/X VGND VGND VPWR VPWR _7340_/C
+ sky130_fd_sc_hd__o221a_1
X_4549_ _9810_/Q _4547_/A hold510/X _4547_/Y VGND VGND VPWR VPWR _9810_/D sky130_fd_sc_hd__a22o_1
X_7268_ _6306_/Y _7173_/X _6352_/Y _7174_/X VGND VGND VPWR VPWR _7268_/X sky130_fd_sc_hd__o22a_1
Xhold485 _5900_/X VGND VGND VPWR VPWR _9202_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold474 _4732_/B VGND VGND VPWR VPWR hold475/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 hold496/A VGND VGND VPWR VPWR _4951_/B sky130_fd_sc_hd__clkbuf_2
X_9007_ _7777_/X _9007_/A1 _9017_/S VGND VGND VPWR VPWR _9007_/X sky130_fd_sc_hd__mux2_1
X_6219_ _9118_/Q VGND VGND VPWR VPWR _6219_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7199_ _7199_/A _7199_/B _7199_/C _7199_/D VGND VGND VPWR VPWR _7209_/B sky130_fd_sc_hd__and4_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6570_ _9159_/Q VGND VGND VPWR VPWR _6570_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5521_ _5570_/A _5521_/B VGND VGND VPWR VPWR _5522_/A sky130_fd_sc_hd__or2_1
X_8240_ _8255_/B VGND VGND VPWR VPWR _8382_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_117_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5452_ _9468_/Q _5446_/A hold217/X _5446_/Y VGND VGND VPWR VPWR _5452_/X sky130_fd_sc_hd__a22o_1
X_5383_ _9515_/Q _5380_/A hold577/A _5380_/Y VGND VGND VPWR VPWR _5383_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8171_ _8255_/A _8171_/B VGND VGND VPWR VPWR _8615_/A sky130_fd_sc_hd__nor2_1
X_7122_ _9288_/Q _9287_/Q _7129_/B _7129_/C VGND VGND VPWR VPWR _7173_/A sky130_fd_sc_hd__or4_4
X_7053_ _7053_/A hold22/X VGND VGND VPWR VPWR _7053_/Y sky130_fd_sc_hd__nor2_2
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6004_ _9139_/Q _6000_/A _6064_/B1 _6000_/Y VGND VGND VPWR VPWR _9139_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7955_ _8118_/A _8296_/B VGND VGND VPWR VPWR _8639_/A sky130_fd_sc_hd__nor2_1
X_7886_ _8042_/B VGND VGND VPWR VPWR _8118_/A sky130_fd_sc_hd__buf_8
X_6906_ _6904_/Y _5428_/B _6905_/Y _5313_/B VGND VGND VPWR VPWR _6906_/X sky130_fd_sc_hd__o22a_1
X_9625_ _9730_/CLK _9625_/D _9797_/SET_B VGND VGND VPWR VPWR _9625_/Q sky130_fd_sc_hd__dfrtp_1
X_6837_ _6837_/A VGND VGND VPWR VPWR _6837_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9556_ _9686_/CLK _9556_/D _7042_/B VGND VGND VPWR VPWR _9556_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6768_ _9390_/Q VGND VGND VPWR VPWR _6768_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8507_ _8229_/A _8312_/B _8138_/B _8594_/A VGND VGND VPWR VPWR _8657_/C sky130_fd_sc_hd__o22ai_1
XFILLER_148_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6699_ _9424_/Q VGND VGND VPWR VPWR _6699_/Y sky130_fd_sc_hd__clkinv_2
X_9487_ _9491_/CLK _9487_/D _9731_/SET_B VGND VGND VPWR VPWR _9487_/Q sky130_fd_sc_hd__dfrtp_4
X_5719_ _5719_/A VGND VGND VPWR VPWR _5719_/Y sky130_fd_sc_hd__inv_2
X_8438_ _8438_/A VGND VGND VPWR VPWR _8438_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8369_ _8369_/A _8641_/C _8548_/C _8735_/C VGND VGND VPWR VPWR _8369_/Y sky130_fd_sc_hd__nor4_2
XFILLER_2_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold260 hold260/A VGND VGND VPWR VPWR hold261/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 hold271/A VGND VGND VPWR VPWR hold272/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _5460_/X VGND VGND VPWR VPWR hold283/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold293/A VGND VGND VPWR VPWR _9117_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_172_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 _8858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _8101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _6106_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_144 _7604_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _4790_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_177 _7052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7740_ _9124_/Q VGND VGND VPWR VPWR _7740_/Y sky130_fd_sc_hd__clkinv_2
X_4952_ _9531_/Q VGND VGND VPWR VPWR _4952_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4883_ _4883_/A _4947_/A VGND VGND VPWR VPWR _4883_/X sky130_fd_sc_hd__or2_4
X_7671_ _6928_/Y _7521_/X _6879_/Y _7522_/X VGND VGND VPWR VPWR _7671_/X sky130_fd_sc_hd__o22a_1
XFILLER_32_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9410_ _9695_/CLK hold83/X _9689_/SET_B VGND VGND VPWR VPWR _9410_/Q sky130_fd_sc_hd__dfrtp_1
X_6622_ _9793_/Q VGND VGND VPWR VPWR _6622_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9341_ _9643_/CLK _9341_/D _9563_/SET_B VGND VGND VPWR VPWR _9341_/Q sky130_fd_sc_hd__dfrtp_1
X_6553_ _9347_/Q VGND VGND VPWR VPWR _6553_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5504_ _5770_/A VGND VGND VPWR VPWR _5698_/A sky130_fd_sc_hd__buf_6
X_9272_ _9431_/CLK _9272_/D _9817_/SET_B VGND VGND VPWR VPWR _9272_/Q sky130_fd_sc_hd__dfrtp_1
X_6484_ _6482_/Y _4883_/X _6483_/Y _4623_/B VGND VGND VPWR VPWR _6484_/X sky130_fd_sc_hd__o22a_4
X_8223_ _8475_/B _8223_/B VGND VGND VPWR VPWR _8225_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput310 _9786_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_2
X_5435_ _9479_/Q _5430_/A _6008_/B1 _5430_/Y VGND VGND VPWR VPWR _9479_/D sky130_fd_sc_hd__a22o_1
XFILLER_133_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 _8863_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_2
Xoutput332 _9783_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_2
Xoutput321 _9796_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_2
Xoutput376 _9078_/Q VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_2
Xoutput365 _9060_/Q VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_2
Xoutput387 _9067_/Q VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_2
X_8154_ _8443_/A _8182_/B VGND VGND VPWR VPWR _8396_/A sky130_fd_sc_hd__nor2_1
Xoutput354 _9809_/Q VGND VGND VPWR VPWR sram_ro_addr[5] sky130_fd_sc_hd__buf_2
X_5366_ _9526_/Q _5361_/A _6008_/B1 _5361_/Y VGND VGND VPWR VPWR _9526_/D sky130_fd_sc_hd__a22o_1
X_5297_ _9573_/Q _5292_/A _6065_/B1 _5292_/Y VGND VGND VPWR VPWR _9573_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8085_ _8563_/A _8596_/A VGND VGND VPWR VPWR _8657_/B sky130_fd_sc_hd__nor2_1
X_7105_ _4761_/Y _7144_/A _4721_/Y _7145_/A _7104_/X VGND VGND VPWR VPWR _7116_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7036_ _7036_/A VGND VGND VPWR VPWR _9090_/D sky130_fd_sc_hd__inv_2
XFILLER_59_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8987_ _8986_/X hold350/X _8987_/S VGND VGND VPWR VPWR _8987_/X sky130_fd_sc_hd__mux2_4
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7938_ _7938_/A _8567_/C VGND VGND VPWR VPWR _8514_/A sky130_fd_sc_hd__or2_2
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9608_ _9651_/CLK _9608_/D _9689_/SET_B VGND VGND VPWR VPWR _9608_/Q sky130_fd_sc_hd__dfrtp_1
X_7869_ _7869_/A _7874_/B _7874_/C VGND VGND VPWR VPWR _7870_/A sky130_fd_sc_hd__or3_1
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9539_ _9576_/CLK _9539_/D _9537_/SET_B VGND VGND VPWR VPWR _9539_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_41_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9800_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5220_ _9624_/Q _5216_/Y _8959_/X _5216_/A VGND VGND VPWR VPWR _9624_/D sky130_fd_sc_hd__o22a_1
XFILLER_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5151_ _9669_/Q _5146_/A _8975_/A1 _5146_/Y VGND VGND VPWR VPWR _5151_/X sky130_fd_sc_hd__a22o_1
X_5082_ _7766_/A _5082_/B VGND VGND VPWR VPWR _5083_/A sky130_fd_sc_hd__and2_1
XFILLER_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8910_ _8909_/X _9215_/Q _9096_/Q VGND VGND VPWR VPWR _8910_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8841_ _8841_/A VGND VGND VPWR VPWR _8842_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8772_ _8772_/A _8772_/B _8772_/C _8772_/D VGND VGND VPWR VPWR _8773_/B sky130_fd_sc_hd__or4_2
X_5984_ _9153_/Q _5981_/A hold696/X _5981_/Y VGND VGND VPWR VPWR _9153_/D sky130_fd_sc_hd__a22o_1
X_7723_ _6394_/Y _7515_/A _6476_/Y _7516_/A VGND VGND VPWR VPWR _7723_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4935_ _4928_/Y _4929_/X _4930_/Y _4598_/B _4934_/X VGND VGND VPWR VPWR _4956_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_193_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_22 _6138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 _4904_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _4866_/A _6189_/A VGND VGND VPWR VPWR _4866_/X sky130_fd_sc_hd__or2_1
X_7654_ _4714_/Y _7519_/X _4905_/Y _7520_/X _7653_/X VGND VGND VPWR VPWR _7657_/C
+ sky130_fd_sc_hd__o221a_1
XANTENNA_66 _7050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7585_ _7585_/A _7585_/B _7585_/C _7585_/D VGND VGND VPWR VPWR _7586_/D sky130_fd_sc_hd__and4_1
XANTENNA_33 _6383_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4797_ _4947_/A _4865_/B VGND VGND VPWR VPWR _5946_/B sky130_fd_sc_hd__or2_4
XANTENNA_44 _6626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6605_ _9555_/Q VGND VGND VPWR VPWR _6605_/Y sky130_fd_sc_hd__inv_2
XANTENNA_55 _6908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _8859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9324_ _9326_/CLK _9324_/D _9571_/SET_B VGND VGND VPWR VPWR _9324_/Q sky130_fd_sc_hd__dfrtp_1
X_6536_ _6536_/A VGND VGND VPWR VPWR _6536_/Y sky130_fd_sc_hd__inv_2
XANTENNA_88 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6467_ _9410_/Q VGND VGND VPWR VPWR _6467_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9255_ _9833_/CLK _9255_/D _9730_/SET_B VGND VGND VPWR VPWR _9255_/Q sky130_fd_sc_hd__dfrtp_1
X_6398_ _9250_/Q VGND VGND VPWR VPWR _6398_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5418_ _5418_/A VGND VGND VPWR VPWR _5419_/A sky130_fd_sc_hd__clkbuf_4
X_8206_ _8206_/A _8750_/D VGND VGND VPWR VPWR _8208_/A sky130_fd_sc_hd__or2_1
X_9186_ _9319_/CLK _9186_/D _9797_/SET_B VGND VGND VPWR VPWR _9186_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5349_ _9537_/Q hold630/X hold593/X _5342_/Y VGND VGND VPWR VPWR _9537_/D sky130_fd_sc_hd__a22o_1
X_8137_ _8137_/A _8137_/B VGND VGND VPWR VPWR _8211_/A sky130_fd_sc_hd__or2_1
XFILLER_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8068_ _8068_/A VGND VGND VPWR VPWR _8563_/A sky130_fd_sc_hd__clkbuf_8
X_7019_ _8854_/A _8851_/A _6993_/B VGND VGND VPWR VPWR _7019_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_75_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4953_/A _4806_/B VGND VGND VPWR VPWR _5927_/B sky130_fd_sc_hd__or2_4
X_4651_ _6083_/B hold1/A VGND VGND VPWR VPWR _6081_/A sky130_fd_sc_hd__nor2_4
XFILLER_174_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR _6288_/A sky130_fd_sc_hd__clkbuf_1
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR _4843_/A sky130_fd_sc_hd__clkbuf_1
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_4
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR _6569_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7370_ _6760_/Y _7149_/X _6669_/Y _7150_/X _7369_/X VGND VGND VPWR VPWR _7375_/B
+ sky130_fd_sc_hd__o221a_1
X_4582_ _6008_/B1 _9798_/Q _4582_/S VGND VGND VPWR VPWR _4583_/A sky130_fd_sc_hd__mux2_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__buf_6
X_6321_ _9523_/Q VGND VGND VPWR VPWR _6321_/Y sky130_fd_sc_hd__clkinv_4
Xinput75 porb VGND VGND VPWR VPWR _7042_/B sky130_fd_sc_hd__buf_12
Xinput97 sram_ro_data[13] VGND VGND VPWR VPWR _6323_/A sky130_fd_sc_hd__clkbuf_1
X_9040_ _9608_/Q _8815_/A VGND VGND VPWR VPWR _9040_/Z sky130_fd_sc_hd__ebufn_1
X_6252_ _6252_/A VGND VGND VPWR VPWR _6252_/Y sky130_fd_sc_hd__clkinv_2
X_5203_ _5203_/A VGND VGND VPWR VPWR _5203_/Y sky130_fd_sc_hd__clkinv_2
X_6183_ _9420_/Q VGND VGND VPWR VPWR _6183_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_130_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5134_ _5134_/A VGND VGND VPWR VPWR _5135_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_111_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5065_ _9013_/X _4572_/B _9719_/Q _5085_/D VGND VGND VPWR VPWR _9719_/D sky130_fd_sc_hd__a22o_1
X_8824_ _8824_/A VGND VGND VPWR VPWR _8824_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5967_ _9101_/Q _5969_/B VGND VGND VPWR VPWR _7032_/B sky130_fd_sc_hd__and2_1
X_8755_ _8755_/A _8755_/B _8755_/C _8755_/D VGND VGND VPWR VPWR _8756_/B sky130_fd_sc_hd__or4_1
XFILLER_25_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8686_ _8719_/D _8761_/C _8773_/A _8717_/D VGND VGND VPWR VPWR _8689_/A sky130_fd_sc_hd__or4_4
XFILLER_80_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7706_ _6535_/Y _7513_/A _6587_/Y _7514_/A _7705_/X VGND VGND VPWR VPWR _7711_/B
+ sky130_fd_sc_hd__o221a_1
X_4918_ _4918_/A _4918_/B _4918_/C _4918_/D VGND VGND VPWR VPWR _4957_/C sky130_fd_sc_hd__and4_1
XFILLER_52_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7637_ _6135_/Y _7527_/X _6097_/Y _7528_/X VGND VGND VPWR VPWR _7637_/X sky130_fd_sc_hd__o22a_1
X_5898_ _9204_/Q _5896_/A _6065_/B1 _5896_/Y VGND VGND VPWR VPWR _5898_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4849_ _9245_/Q VGND VGND VPWR VPWR _4849_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7568_ _7568_/A _7568_/B _7568_/C _7568_/D VGND VGND VPWR VPWR _7568_/Y sky130_fd_sc_hd__nand4_2
X_7499_ _6849_/Y _7498_/X _6926_/Y _5727_/X VGND VGND VPWR VPWR _7499_/X sky130_fd_sc_hd__o22a_1
X_6519_ _8803_/A _5636_/B _6515_/Y _5620_/B _6518_/X VGND VGND VPWR VPWR _6532_/B
+ sky130_fd_sc_hd__o221a_1
X_9307_ _9831_/CLK _9307_/D _9727_/SET_B VGND VGND VPWR VPWR _9307_/Q sky130_fd_sc_hd__dfrtp_1
X_9238_ _9830_/CLK _9238_/D _9537_/SET_B VGND VGND VPWR VPWR _9238_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9169_ _9491_/CLK _9169_/D _9731_/SET_B VGND VGND VPWR VPWR _9169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6870_ _9799_/Q VGND VGND VPWR VPWR _6870_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5821_ _9258_/Q _5820_/A _8959_/A1 _5820_/Y VGND VGND VPWR VPWR _9258_/D sky130_fd_sc_hd__a22o_1
X_8540_ _8540_/A _8540_/B VGND VGND VPWR VPWR _8737_/A sky130_fd_sc_hd__nor2_1
X_5752_ _5753_/B _5752_/B _7072_/A VGND VGND VPWR VPWR _5752_/Y sky130_fd_sc_hd__nor3_1
X_4703_ input61/X _4700_/Y _4701_/Y _6083_/C VGND VGND VPWR VPWR _4703_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8471_ _8745_/A _8627_/B VGND VGND VPWR VPWR _8602_/B sky130_fd_sc_hd__or2_1
X_5683_ _5673_/A _5685_/A _5780_/C VGND VGND VPWR VPWR _5683_/Y sky130_fd_sc_hd__o21ai_1
X_4634_ _5282_/A _4634_/B VGND VGND VPWR VPWR _4634_/X sky130_fd_sc_hd__or2_1
X_7422_ _6361_/Y _7173_/A _6366_/Y _7174_/A VGND VGND VPWR VPWR _7422_/X sky130_fd_sc_hd__o22a_1
Xhold612 hold42/X VGND VGND VPWR VPWR hold612/X sky130_fd_sc_hd__buf_4
X_4565_ _9108_/Q VGND VGND VPWR VPWR _8852_/A sky130_fd_sc_hd__inv_2
Xhold601 hold601/A VGND VGND VPWR VPWR hold601/X sky130_fd_sc_hd__buf_8
X_7353_ _7353_/A _7353_/B _7353_/C _7353_/D VGND VGND VPWR VPWR _7363_/B sky130_fd_sc_hd__and4_1
Xhold634 _5462_/X VGND VGND VPWR VPWR _9461_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold645 _5604_/X VGND VGND VPWR VPWR _9366_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_162_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold623 _4869_/X VGND VGND VPWR VPWR _5290_/B sky130_fd_sc_hd__clkbuf_2
X_6304_ _6299_/Y _4545_/B _6300_/Y _5482_/B _6303_/X VGND VGND VPWR VPWR _6311_/C
+ sky130_fd_sc_hd__o221a_1
Xhold656 _9705_/Q VGND VGND VPWR VPWR hold656/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_143_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7284_ _6201_/Y _7155_/X _6232_/Y _7156_/X _7283_/X VGND VGND VPWR VPWR _7287_/C
+ sky130_fd_sc_hd__o221a_1
X_4496_ _4808_/A _4832_/A _5250_/A VGND VGND VPWR VPWR _4497_/S sky130_fd_sc_hd__or3_1
Xhold667 _5481_/X VGND VGND VPWR VPWR _9448_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_9023_ _9624_/Q _7735_/A VGND VGND VPWR VPWR _9023_/Z sky130_fd_sc_hd__ebufn_1
Xhold678 _5437_/X VGND VGND VPWR VPWR _5438_/A sky130_fd_sc_hd__clkbuf_2
Xhold689 _5241_/A VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__clkbuf_2
X_6235_ _6230_/Y _5263_/B _6231_/Y _5417_/B _6234_/X VGND VGND VPWR VPWR _6242_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_103_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6166_ _6166_/A VGND VGND VPWR VPWR _8975_/S sky130_fd_sc_hd__inv_8
XFILLER_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _9693_/Q _5114_/A hold577/A _5114_/Y VGND VGND VPWR VPWR _5117_/X sky130_fd_sc_hd__a22o_1
X_6097_ _9318_/Q VGND VGND VPWR VPWR _6097_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5048_ _5048_/A VGND VGND VPWR VPWR _5049_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8807_ _8807_/A VGND VGND VPWR VPWR _8808_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9787_ _9791_/CLK _9787_/D _9797_/SET_B VGND VGND VPWR VPWR _9787_/Q sky130_fd_sc_hd__dfstp_1
X_8738_ _8738_/A _8738_/B _8738_/C _8769_/D VGND VGND VPWR VPWR _8739_/A sky130_fd_sc_hd__or4_1
X_6999_ _6506_/Y _6995_/A _9066_/Q _6995_/Y VGND VGND VPWR VPWR _9066_/D sky130_fd_sc_hd__o22a_2
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8669_ _8669_/A _8669_/B _8669_/C _8669_/D VGND VGND VPWR VPWR _8728_/D sky130_fd_sc_hd__or4_2
XFILLER_193_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6020_ _6081_/A VGND VGND VPWR VPWR _6071_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7971_ _8436_/B _8340_/A _7970_/X VGND VGND VPWR VPWR _7972_/B sky130_fd_sc_hd__o21ai_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6922_ _9299_/Q VGND VGND VPWR VPWR _6922_/Y sky130_fd_sc_hd__inv_2
X_9710_ _9731_/CLK _9710_/D _9731_/SET_B VGND VGND VPWR VPWR _9710_/Q sky130_fd_sc_hd__dfstp_1
X_9641_ _9643_/CLK _9641_/D _9689_/SET_B VGND VGND VPWR VPWR _9641_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6853_ _6848_/Y _4854_/X _6849_/Y _5417_/B _6852_/X VGND VGND VPWR VPWR _6860_/C
+ sky130_fd_sc_hd__o221a_1
X_5804_ _9268_/Q _5799_/A _6008_/B1 _5799_/Y VGND VGND VPWR VPWR _9268_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6784_ _9434_/Q VGND VGND VPWR VPWR _6784_/Y sky130_fd_sc_hd__inv_2
X_9572_ _9574_/CLK _9572_/D _9571_/SET_B VGND VGND VPWR VPWR _9572_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8523_ _8523_/A _8748_/A VGND VGND VPWR VPWR _8525_/A sky130_fd_sc_hd__or2_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5735_ _9294_/Q VGND VGND VPWR VPWR _7479_/A sky130_fd_sc_hd__clkinv_2
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8454_ _8592_/A _8443_/B _8451_/X _8453_/Y VGND VGND VPWR VPWR _8454_/X sky130_fd_sc_hd__o211a_1
X_5666_ _9321_/Q VGND VGND VPWR VPWR _5675_/B sky130_fd_sc_hd__inv_2
XFILLER_190_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4617_ _9778_/Q _4613_/A _6064_/B1 _4613_/Y VGND VGND VPWR VPWR _9778_/D sky130_fd_sc_hd__a22o_1
X_7405_ _6618_/Y _7180_/A _6511_/Y _7181_/A _7404_/X VGND VGND VPWR VPWR _7406_/D
+ sky130_fd_sc_hd__o221a_1
X_8385_ _7925_/B _8043_/Y _8151_/C VGND VGND VPWR VPWR _8385_/Y sky130_fd_sc_hd__o21ai_2
X_5597_ _5770_/A VGND VGND VPWR VPWR _5847_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold420 _5897_/X VGND VGND VPWR VPWR hold421/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 hold442/A VGND VGND VPWR VPWR hold443/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 hold431/A VGND VGND VPWR VPWR hold432/A sky130_fd_sc_hd__dlygate4sd3_1
X_7336_ _7336_/A _7380_/B VGND VGND VPWR VPWR _7336_/X sky130_fd_sc_hd__or2_1
Xhold453 _4937_/X VGND VGND VPWR VPWR _5444_/B sky130_fd_sc_hd__clkbuf_2
X_4548_ _9811_/Q _4547_/A hold516/X _4547_/Y VGND VGND VPWR VPWR _4548_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7267_ _6315_/Y _7071_/D _6308_/Y _7166_/X _7266_/X VGND VGND VPWR VPWR _7274_/A
+ sky130_fd_sc_hd__o221a_1
Xhold486 _5662_/X VGND VGND VPWR VPWR _9326_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold464 _5659_/X VGND VGND VPWR VPWR hold465/A sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ _4689_/C VGND VGND VPWR VPWR _4750_/A sky130_fd_sc_hd__clkinv_2
Xhold475 hold475/A VGND VGND VPWR VPWR _4764_/B sky130_fd_sc_hd__clkbuf_2
X_9006_ _7775_/X _9006_/A1 _9017_/S VGND VGND VPWR VPWR _9006_/X sky130_fd_sc_hd__mux2_1
X_6218_ _6218_/A _6218_/B _6218_/C VGND VGND VPWR VPWR _6268_/B sky130_fd_sc_hd__and3_1
Xhold497 _4498_/X VGND VGND VPWR VPWR hold498/A sky130_fd_sc_hd__dlygate4sd3_1
X_7198_ _6668_/Y _7160_/X _6804_/Y _7071_/B _7197_/X VGND VGND VPWR VPWR _7199_/D
+ sky130_fd_sc_hd__o221a_1
X_6149_ _6144_/Y _5406_/B _6145_/Y _5378_/B _6148_/X VGND VGND VPWR VPWR _6150_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5520_ _9422_/Q _5515_/A _6008_/B1 _5515_/Y VGND VGND VPWR VPWR _5520_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5451_ _9469_/Q _5446_/A _6065_/B1 _5446_/Y VGND VGND VPWR VPWR _9469_/D sky130_fd_sc_hd__a22o_1
XFILLER_117_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5382_ _9516_/Q _5380_/A hold510/X _5380_/Y VGND VGND VPWR VPWR _5382_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8170_ _8171_/B _8182_/B VGND VGND VPWR VPWR _8399_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7121_ _7127_/A _7121_/B VGND VGND VPWR VPWR _7172_/A sky130_fd_sc_hd__or2_2
X_7052_ _7052_/A VGND VGND VPWR VPWR _7052_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_140_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6003_ _9140_/Q _5999_/X hold577/A _6000_/Y VGND VGND VPWR VPWR _6003_/X sky130_fd_sc_hd__a22o_1
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7954_ _8268_/C _8361_/A VGND VGND VPWR VPWR _8296_/B sky130_fd_sc_hd__or2_1
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6905_ _9558_/Q VGND VGND VPWR VPWR _6905_/Y sky130_fd_sc_hd__clkinv_2
X_7885_ _8436_/A _8436_/B _8436_/C _8236_/A VGND VGND VPWR VPWR _8042_/B sky130_fd_sc_hd__or4_4
X_9624_ _9730_/CLK _9624_/D _9797_/SET_B VGND VGND VPWR VPWR _9624_/Q sky130_fd_sc_hd__dfrtp_2
X_6836_ _9597_/Q VGND VGND VPWR VPWR _6836_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6767_ _9520_/Q VGND VGND VPWR VPWR _6767_/Y sky130_fd_sc_hd__inv_2
X_9555_ _9686_/CLK _9555_/D _7042_/B VGND VGND VPWR VPWR _9555_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8506_ _8506_/A _8506_/B _8710_/A _8506_/D VGND VGND VPWR VPWR _8508_/A sky130_fd_sc_hd__or4_1
X_5718_ _5718_/A _9097_/Q VGND VGND VPWR VPWR _5719_/A sky130_fd_sc_hd__or2_2
X_6698_ _9711_/Q VGND VGND VPWR VPWR _6698_/Y sky130_fd_sc_hd__clkinv_2
X_9486_ _9491_/CLK _9486_/D _9731_/SET_B VGND VGND VPWR VPWR _9486_/Q sky130_fd_sc_hd__dfrtp_1
X_5649_ _5649_/A VGND VGND VPWR VPWR _5649_/Y sky130_fd_sc_hd__inv_2
X_8437_ _8489_/A _8437_/B VGND VGND VPWR VPWR _8437_/X sky130_fd_sc_hd__or2_1
XFILLER_40_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8368_ _8510_/A _8757_/B VGND VGND VPWR VPWR _8735_/C sky130_fd_sc_hd__or2_1
Xhold261 hold261/A VGND VGND VPWR VPWR hold261/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold250 hold250/A VGND VGND VPWR VPWR _9569_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7319_ _7319_/A _7319_/B _7319_/C VGND VGND VPWR VPWR _7319_/Y sky130_fd_sc_hd__nand3_4
Xhold272 hold272/A VGND VGND VPWR VPWR _9333_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold294 _5334_/X VGND VGND VPWR VPWR hold295/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/A VGND VGND VPWR VPWR hold284/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8299_ _8299_/A _8716_/B VGND VGND VPWR VPWR _8301_/A sky130_fd_sc_hd__or2_1
XFILLER_2_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_123 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _8628_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _6230_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_145 _6083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_178 _7052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _5263_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_1_1_csclk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4951_ _4951_/A _4951_/B VGND VGND VPWR VPWR _5482_/B sky130_fd_sc_hd__or2_4
X_7670_ _6914_/Y _7513_/X _6904_/Y _7514_/X _7669_/X VGND VGND VPWR VPWR _7675_/B
+ sky130_fd_sc_hd__o221a_1
X_4882_ _4882_/A VGND VGND VPWR VPWR _4882_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6621_ _8819_/A _5329_/B _6620_/Y _5389_/B VGND VGND VPWR VPWR _6621_/X sky130_fd_sc_hd__o22a_1
X_9340_ _9421_/CLK _9340_/D _9537_/SET_B VGND VGND VPWR VPWR _9340_/Q sky130_fd_sc_hd__dfrtp_1
X_6552_ _6552_/A VGND VGND VPWR VPWR _6552_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_185_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5503_ _9432_/Q _5495_/A hold601/A _5495_/Y VGND VGND VPWR VPWR _5503_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6483_ _9772_/Q VGND VGND VPWR VPWR _6483_/Y sky130_fd_sc_hd__inv_2
X_9271_ _9431_/CLK _9271_/D _9817_/SET_B VGND VGND VPWR VPWR _9271_/Q sky130_fd_sc_hd__dfrtp_1
X_8222_ _8693_/A _8604_/A _8678_/A _8221_/Y VGND VGND VPWR VPWR _8223_/B sky130_fd_sc_hd__or4b_1
Xoutput300 _9765_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_2
X_5434_ _9480_/Q _5430_/A _6067_/B1 _5430_/Y VGND VGND VPWR VPWR _9480_/D sky130_fd_sc_hd__a22o_1
X_8153_ _8153_/A VGND VGND VPWR VPWR _8432_/B sky130_fd_sc_hd__inv_4
XFILLER_126_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput344 _8846_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_2
Xoutput311 _9787_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_2
Xoutput322 _9797_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_2
Xoutput333 _9086_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_2
Xoutput377 _9079_/Q VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput366 _9061_/Q VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7104_ _4794_/Y _7067_/A _4684_/Y _7146_/A VGND VGND VPWR VPWR _7104_/X sky130_fd_sc_hd__o22a_1
Xoutput355 _9810_/Q VGND VGND VPWR VPWR sram_ro_addr[6] sky130_fd_sc_hd__buf_2
X_5365_ _9527_/Q _5361_/A _6067_/B1 _5361_/Y VGND VGND VPWR VPWR _9527_/D sky130_fd_sc_hd__a22o_1
Xoutput388 _9068_/Q VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_2
X_5296_ _9574_/Q _5292_/A _6064_/B1 _5292_/Y VGND VGND VPWR VPWR _9574_/D sky130_fd_sc_hd__a22o_1
X_8084_ _8138_/B _8594_/A _8083_/X VGND VGND VPWR VPWR _8086_/A sky130_fd_sc_hd__o21ai_1
X_7035_ _4987_/B _7039_/A _7039_/B _6053_/B _7034_/X VGND VGND VPWR VPWR _7036_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8986_ hold619/X _4971_/A _9093_/Q VGND VGND VPWR VPWR _8986_/X sky130_fd_sc_hd__mux2_2
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7937_ _8048_/C _7937_/B VGND VGND VPWR VPWR _8567_/C sky130_fd_sc_hd__or2_4
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7868_ _8366_/A VGND VGND VPWR VPWR _7868_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9607_ _9651_/CLK _9607_/D _9563_/SET_B VGND VGND VPWR VPWR _9607_/Q sky130_fd_sc_hd__dfrtp_2
X_6819_ _9571_/Q VGND VGND VPWR VPWR _6819_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7799_ _7933_/B VGND VGND VPWR VPWR _8230_/A sky130_fd_sc_hd__clkinv_2
XFILLER_11_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9538_ _9576_/CLK _9538_/D _9537_/SET_B VGND VGND VPWR VPWR _9538_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9469_ _9577_/CLK _9469_/D _9571_/SET_B VGND VGND VPWR VPWR _9469_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ _9670_/Q _5146_/A _8969_/A1 _5146_/Y VGND VGND VPWR VPWR _9670_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5081_ _7766_/A _5081_/B VGND VGND VPWR VPWR _5081_/X sky130_fd_sc_hd__and2_1
XFILLER_123_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8840_ _8840_/A VGND VGND VPWR VPWR _8840_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5983_ _9154_/Q _5981_/A hold510/X _5981_/Y VGND VGND VPWR VPWR _9154_/D sky130_fd_sc_hd__a22o_1
X_8771_ _8771_/A VGND VGND VPWR VPWR _8771_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4934_ _6189_/A _4947_/A _4931_/Y _4932_/Y _5301_/B VGND VGND VPWR VPWR _4934_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_40_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7722_ _6405_/Y _7507_/A _6418_/Y _7508_/A _7721_/X VGND VGND VPWR VPWR _7729_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_23 _6142_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4865_ _4865_/A _4865_/B VGND VGND VPWR VPWR _4865_/X sky130_fd_sc_hd__or2_4
XFILLER_32_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7653_ _4705_/Y _7521_/X _4910_/Y _7522_/X VGND VGND VPWR VPWR _7653_/X sky130_fd_sc_hd__o22a_1
XANTENNA_12 _4932_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_45 _6706_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7584_ _6499_/Y _7525_/X _7248_/A _7526_/X _7583_/X VGND VGND VPWR VPWR _7585_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA_34 _6380_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _9162_/Q VGND VGND VPWR VPWR _4796_/Y sky130_fd_sc_hd__inv_2
XANTENNA_56 _7095_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6604_ _8831_/A _5340_/B _6600_/Y _4611_/B _6603_/X VGND VGND VPWR VPWR _6617_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_67 _7050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_78 _8843_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9323_ _9728_/CLK _9323_/D _9571_/SET_B VGND VGND VPWR VPWR _9323_/Q sky130_fd_sc_hd__dfrtp_1
X_6535_ _9230_/Q VGND VGND VPWR VPWR _6535_/Y sky130_fd_sc_hd__inv_2
XANTENNA_89 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9254_ _9833_/CLK _9254_/D _9730_/SET_B VGND VGND VPWR VPWR _9254_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8205_ _8205_/A _8209_/A VGND VGND VPWR VPWR _8750_/D sky130_fd_sc_hd__nor2_1
X_6466_ _9678_/Q VGND VGND VPWR VPWR _6466_/Y sky130_fd_sc_hd__inv_2
X_5417_ _5570_/A _5417_/B VGND VGND VPWR VPWR _5418_/A sky130_fd_sc_hd__or2_1
X_6397_ _6384_/Y _5847_/B _6386_/X _6390_/X _6396_/X VGND VGND VPWR VPWR _6506_/B
+ sky130_fd_sc_hd__o2111a_2
X_9185_ _9212_/CLK _9185_/D _9797_/SET_B VGND VGND VPWR VPWR _9185_/Q sky130_fd_sc_hd__dfrtp_1
X_8136_ _8563_/A _8479_/B VGND VGND VPWR VPWR _8602_/A sky130_fd_sc_hd__nor2_1
X_5348_ _9538_/Q _5342_/A hold136/X _5342_/Y VGND VGND VPWR VPWR _5348_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8067_ _8429_/A _8178_/B _8053_/A _8178_/B _8066_/X VGND VGND VPWR VPWR _8067_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7018_ _8852_/A _8851_/A _7005_/A VGND VGND VPWR VPWR _7018_/Y sky130_fd_sc_hd__o21ai_1
X_5279_ _9585_/Q _5276_/A _8965_/A1 _5276_/Y VGND VGND VPWR VPWR _9585_/D sky130_fd_sc_hd__a22o_1
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8969_ _9661_/Q _8969_/A1 _8973_/S VGND VGND VPWR VPWR _8969_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4650_ _9831_/Q _9138_/Q hold35/X VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__or3_4
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR _6116_/A sky130_fd_sc_hd__clkbuf_1
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR _6862_/A sky130_fd_sc_hd__clkbuf_1
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR _6711_/A sky130_fd_sc_hd__clkbuf_1
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR _4775_/A sky130_fd_sc_hd__clkbuf_1
X_6320_ _9795_/Q VGND VGND VPWR VPWR _6320_/Y sky130_fd_sc_hd__inv_2
X_4581_ _4581_/A VGND VGND VPWR VPWR _9799_/D sky130_fd_sc_hd__clkbuf_1
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR _6184_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _8859_/A sky130_fd_sc_hd__buf_4
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _8858_/A sky130_fd_sc_hd__buf_6
XFILLER_143_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput76 qspi_enabled VGND VGND VPWR VPWR _8877_/S sky130_fd_sc_hd__buf_6
Xinput98 sram_ro_data[14] VGND VGND VPWR VPWR _6252_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_182_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6251_ _9796_/Q VGND VGND VPWR VPWR _6251_/Y sky130_fd_sc_hd__inv_2
X_5202_ _5202_/A VGND VGND VPWR VPWR _5203_/A sky130_fd_sc_hd__buf_2
X_6182_ _9386_/Q VGND VGND VPWR VPWR _6182_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5133_ _5378_/A _5133_/B VGND VGND VPWR VPWR _5134_/A sky130_fd_sc_hd__or2_1
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5064_ _9014_/X _4572_/B _9720_/Q _5085_/D VGND VGND VPWR VPWR _9720_/D sky130_fd_sc_hd__a22o_1
X_8823_ _8823_/A VGND VGND VPWR VPWR _8824_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5966_ _5966_/A _5966_/B _5966_/C _5966_/D VGND VGND VPWR VPWR _5969_/B sky130_fd_sc_hd__or4_2
X_8754_ _8780_/A _8754_/B VGND VGND VPWR VPWR _8754_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5897_ _9205_/Q _5895_/X _6064_/B1 _5896_/Y VGND VGND VPWR VPWR _5897_/X sky130_fd_sc_hd__a22o_1
X_8685_ _8027_/Y _8432_/B _8359_/B _8406_/D _8618_/D VGND VGND VPWR VPWR _8717_/D
+ sky130_fd_sc_hd__a2111o_2
X_4917_ _4909_/Y _4611_/B _4910_/Y _5321_/B _4916_/X VGND VGND VPWR VPWR _4918_/D
+ sky130_fd_sc_hd__o221a_1
X_7705_ _6539_/Y _7515_/A _6582_/Y _7516_/A VGND VGND VPWR VPWR _7705_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7636_ _6096_/Y _7519_/X _6110_/Y _7520_/X _7635_/X VGND VGND VPWR VPWR _7639_/C
+ sky130_fd_sc_hd__o221a_1
X_4848_ _6142_/A _4848_/B VGND VGND VPWR VPWR _4848_/X sky130_fd_sc_hd__or2_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7567_ _7567_/A _7567_/B _7567_/C _7567_/D VGND VGND VPWR VPWR _7568_/D sky130_fd_sc_hd__and4_1
X_4779_ _4770_/Y _5628_/B _4772_/Y _5570_/B _4778_/X VGND VGND VPWR VPWR _4811_/A
+ sky130_fd_sc_hd__o221a_1
X_9306_ _9831_/CLK _9306_/D _9727_/SET_B VGND VGND VPWR VPWR _9306_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6518_ _6516_/Y _5609_/B _6517_/Y _4715_/X VGND VGND VPWR VPWR _6518_/X sky130_fd_sc_hd__o22a_1
X_7498_ _7498_/A VGND VGND VPWR VPWR _7498_/X sky130_fd_sc_hd__buf_4
X_9237_ _9421_/CLK _9237_/D _9537_/SET_B VGND VGND VPWR VPWR _9237_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6449_ _9729_/Q VGND VGND VPWR VPWR _6449_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_164_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9168_ _9491_/CLK _9168_/D _9731_/SET_B VGND VGND VPWR VPWR _9168_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_csclk clkbuf_2_0_0_csclk/X VGND VGND VPWR VPWR _9561_/CLK sky130_fd_sc_hd__clkbuf_16
X_8119_ _8119_/A _8714_/B VGND VGND VPWR VPWR _8123_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9099_ _9322_/CLK _9099_/D _9821_/SET_B VGND VGND VPWR VPWR _9099_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_2_0_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5820_ _5820_/A VGND VGND VPWR VPWR _5820_/Y sky130_fd_sc_hd__inv_2
X_5751_ _7113_/A _7108_/C VGND VGND VPWR VPWR _7072_/A sky130_fd_sc_hd__or2_1
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8470_ _8729_/B _8470_/B VGND VGND VPWR VPWR _8472_/A sky130_fd_sc_hd__or2_1
X_4702_ _4808_/A _4898_/B VGND VGND VPWR VPWR _6083_/C sky130_fd_sc_hd__or2_4
XFILLER_187_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5682_ _5752_/B VGND VGND VPWR VPWR _5723_/A sky130_fd_sc_hd__buf_4
X_7421_ _6465_/Y _7070_/A _6394_/Y _7166_/A _7420_/X VGND VGND VPWR VPWR _7428_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4633_ _4883_/A _4900_/A VGND VGND VPWR VPWR _4634_/B sky130_fd_sc_hd__or2_4
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold602 hold602/A VGND VGND VPWR VPWR hold602/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4564_ _9106_/Q VGND VGND VPWR VPWR _8853_/A sky130_fd_sc_hd__inv_2
X_7352_ _6928_/Y _7160_/X _6864_/Y _7071_/B _7351_/X VGND VGND VPWR VPWR _7353_/D
+ sky130_fd_sc_hd__o221a_1
Xhold613 _8967_/X VGND VGND VPWR VPWR hold613/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold635 _5456_/X VGND VGND VPWR VPWR _5457_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7283_ _6221_/Y _7095_/B _6210_/Y _7157_/X VGND VGND VPWR VPWR _7283_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold624 _4534_/D VGND VGND VPWR VPWR _4708_/B sky130_fd_sc_hd__buf_2
X_6303_ _6301_/Y _4883_/X _6302_/Y _5301_/B VGND VGND VPWR VPWR _6303_/X sky130_fd_sc_hd__o22a_1
Xhold668 _5231_/X VGND VGND VPWR VPWR _9615_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_4495_ _6083_/A VGND VGND VPWR VPWR _5250_/A sky130_fd_sc_hd__buf_8
X_6234_ _6232_/Y _6112_/B _6233_/Y _4611_/B VGND VGND VPWR VPWR _6234_/X sky130_fd_sc_hd__o22a_1
Xhold646 _5705_/X VGND VGND VPWR VPWR _9306_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold657 _4641_/X VGND VGND VPWR VPWR _9763_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold679 _5478_/X VGND VGND VPWR VPWR _9451_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_9022_ _9623_/Q _7737_/A VGND VGND VPWR VPWR _9022_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_89_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6165_ _6165_/A VGND VGND VPWR VPWR _8971_/S sky130_fd_sc_hd__inv_8
XFILLER_85_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _9694_/Q _5114_/A hold510/X _5114_/Y VGND VGND VPWR VPWR _5116_/X sky130_fd_sc_hd__a22o_1
X_6096_ _9226_/Q VGND VGND VPWR VPWR _6096_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5047_ _5282_/A _5047_/B VGND VGND VPWR VPWR _5048_/A sky130_fd_sc_hd__or2_1
XFILLER_150_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8806_ _8806_/A VGND VGND VPWR VPWR _8806_/X sky130_fd_sc_hd__clkbuf_1
X_6998_ _6357_/Y _6995_/A _9067_/Q _6995_/Y VGND VGND VPWR VPWR _9067_/D sky130_fd_sc_hd__o22a_1
X_9786_ _9791_/CLK _9786_/D _9821_/SET_B VGND VGND VPWR VPWR _9786_/Q sky130_fd_sc_hd__dfrtp_1
X_8737_ _8737_/A _8737_/B _8737_/C _8737_/D VGND VGND VPWR VPWR _8769_/D sky130_fd_sc_hd__or4_2
XFILLER_13_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5949_ _9166_/Q _5948_/A _8959_/A1 _5948_/Y VGND VGND VPWR VPWR _9166_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8668_ _8443_/A _8666_/X _8158_/A _8667_/Y VGND VGND VPWR VPWR _8671_/B sky130_fd_sc_hd__o22ai_2
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8599_ _8428_/A _8011_/A _8429_/A _7866_/A _8598_/Y VGND VGND VPWR VPWR _8600_/A
+ sky130_fd_sc_hd__o311a_1
X_7619_ _6219_/Y _7527_/X _6210_/Y _7528_/X VGND VGND VPWR VPWR _7619_/X sky130_fd_sc_hd__o22a_1
XFILLER_175_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput200 wb_sel_i[2] VGND VGND VPWR VPWR _7765_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7970_ _7970_/A _7970_/B VGND VGND VPWR VPWR _7970_/X sky130_fd_sc_hd__and2_1
XFILLER_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6921_ _9261_/Q VGND VGND VPWR VPWR _6921_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9640_ _9643_/CLK _9640_/D _9689_/SET_B VGND VGND VPWR VPWR _9640_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6852_ _6850_/Y _5455_/B _6851_/Y _4883_/X VGND VGND VPWR VPWR _6852_/X sky130_fd_sc_hd__o22a_1
X_9571_ _9574_/CLK _9571_/D _9571_/SET_B VGND VGND VPWR VPWR _9571_/Q sky130_fd_sc_hd__dfstp_1
X_5803_ _9269_/Q _5799_/A _6067_/B1 _5799_/Y VGND VGND VPWR VPWR _9269_/D sky130_fd_sc_hd__a22o_1
X_8522_ _8557_/B _8479_/B _8563_/B _8479_/B VGND VGND VPWR VPWR _8748_/A sky130_fd_sc_hd__o22ai_2
X_6783_ _6779_/Y _5647_/B _6780_/Y _6083_/C _6782_/X VGND VGND VPWR VPWR _6790_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5734_ _7436_/B _5732_/Y _9097_/Q _5733_/X VGND VGND VPWR VPWR _9295_/D sky130_fd_sc_hd__a31o_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5665_ _9323_/Q _5660_/A _6008_/B1 _5660_/Y VGND VGND VPWR VPWR _9323_/D sky130_fd_sc_hd__a22o_1
X_8453_ _8776_/B _8616_/A VGND VGND VPWR VPWR _8453_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8384_ _8155_/Y _8156_/Y _8636_/B VGND VGND VPWR VPWR _8398_/A sky130_fd_sc_hd__a21o_1
X_4616_ _9779_/Q _4613_/A hold696/X _4613_/Y VGND VGND VPWR VPWR _9779_/D sky130_fd_sc_hd__a22o_1
X_7404_ _6580_/Y _7182_/A _6640_/Y _7183_/A VGND VGND VPWR VPWR _7404_/X sky130_fd_sc_hd__o22a_1
XFILLER_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold410 hold410/A VGND VGND VPWR VPWR hold411/A sky130_fd_sc_hd__dlygate4sd3_1
X_7335_ _4786_/Y _7171_/X _4942_/Y _7172_/X _7334_/X VGND VGND VPWR VPWR _7340_/B
+ sky130_fd_sc_hd__o221a_1
X_5596_ _9370_/Q _5591_/A _6008_/B1 _5591_/Y VGND VGND VPWR VPWR _9370_/D sky130_fd_sc_hd__a22o_1
Xhold443 hold443/A VGND VGND VPWR VPWR _6060_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold421 hold421/A VGND VGND VPWR VPWR hold422/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 hold432/A VGND VGND VPWR VPWR _9138_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold454 _6117_/B VGND VGND VPWR VPWR _4933_/B sky130_fd_sc_hd__buf_2
XFILLER_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4547_ _4547_/A VGND VGND VPWR VPWR _4547_/Y sky130_fd_sc_hd__clkinv_2
X_7266_ _6351_/Y _7167_/X _6333_/Y _7168_/X VGND VGND VPWR VPWR _7266_/X sky130_fd_sc_hd__o22a_1
Xhold476 _5453_/X VGND VGND VPWR VPWR hold477/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold465 hold465/A VGND VGND VPWR VPWR hold466/A sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _4682_/C _4508_/B _4685_/C VGND VGND VPWR VPWR _4883_/A sky130_fd_sc_hd__or3_4
Xhold487 _5254_/X VGND VGND VPWR VPWR _9601_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_9005_ _7773_/X _9005_/A1 _9017_/S VGND VGND VPWR VPWR _9005_/X sky130_fd_sc_hd__mux2_1
X_6217_ _7292_/A _5636_/B _6213_/Y _5805_/B _6216_/X VGND VGND VPWR VPWR _6218_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7197_ _6670_/Y _7161_/X _6792_/Y _7162_/X VGND VGND VPWR VPWR _7197_/X sky130_fd_sc_hd__o22a_1
XFILLER_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold498 hold498/A VGND VGND VPWR VPWR hold499/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6148_ _6146_/Y _4585_/B _6147_/Y _4511_/B VGND VGND VPWR VPWR _6148_/X sky130_fd_sc_hd__o22a_4
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _6081_/A VGND VGND VPWR VPWR _6080_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_57_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9769_ _9817_/CLK _9769_/D _9821_/SET_B VGND VGND VPWR VPWR _9769_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5450_ _9470_/Q _5446_/A _6064_/B1 _5446_/Y VGND VGND VPWR VPWR _5450_/X sky130_fd_sc_hd__a22o_1
XFILLER_172_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5381_ _9517_/Q _5380_/A hold516/X _5380_/Y VGND VGND VPWR VPWR _5381_/X sky130_fd_sc_hd__a22o_1
XFILLER_160_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7120_ _4737_/Y _7070_/A _4826_/Y _7166_/A _7119_/X VGND VGND VPWR VPWR _7132_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _9322_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_115_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7051_ _9628_/Q _7051_/B VGND VGND VPWR VPWR _7052_/A sky130_fd_sc_hd__and2b_1
X_6002_ _9141_/Q _6000_/A hold510/X _6000_/Y VGND VGND VPWR VPWR _6002_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7953_ _7953_/A _8288_/B VGND VGND VPWR VPWR _8359_/A sky130_fd_sc_hd__nor2_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6904_ _9480_/Q VGND VGND VPWR VPWR _6904_/Y sky130_fd_sc_hd__clkinv_2
X_7884_ _8347_/A VGND VGND VPWR VPWR _8229_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9623_ _9734_/CLK _9623_/D _9731_/SET_B VGND VGND VPWR VPWR _9623_/Q sky130_fd_sc_hd__dfrtp_4
X_6835_ _6830_/Y _5935_/B _6831_/Y _5971_/B _6834_/X VGND VGND VPWR VPWR _6861_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6766_ _9564_/Q VGND VGND VPWR VPWR _6766_/Y sky130_fd_sc_hd__inv_2
X_9554_ _9686_/CLK _9554_/D _7042_/B VGND VGND VPWR VPWR _9554_/Q sky130_fd_sc_hd__dfstp_1
X_8505_ _8505_/A _8727_/A VGND VGND VPWR VPWR _8506_/D sky130_fd_sc_hd__or2_1
XFILLER_10_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5717_ _9095_/Q VGND VGND VPWR VPWR _5718_/A sky130_fd_sc_hd__inv_2
X_9485_ _9491_/CLK _9485_/D _9731_/SET_B VGND VGND VPWR VPWR _9485_/Q sky130_fd_sc_hd__dfstp_1
X_6697_ _6692_/Y _5598_/B _6693_/Y _5581_/B _6696_/X VGND VGND VPWR VPWR _6722_/C
+ sky130_fd_sc_hd__o221a_1
X_5648_ _5648_/A VGND VGND VPWR VPWR _5649_/A sky130_fd_sc_hd__clkbuf_4
X_8436_ _8436_/A _8436_/B _8436_/C _8436_/D VGND VGND VPWR VPWR _8437_/B sky130_fd_sc_hd__or4_1
XFILLER_136_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5579_ _9381_/Q _5572_/A _8969_/A1 _5572_/Y VGND VGND VPWR VPWR _9381_/D sky130_fd_sc_hd__a22o_1
X_8367_ _8367_/A VGND VGND VPWR VPWR _8510_/A sky130_fd_sc_hd__inv_2
Xhold251 _9703_/Q VGND VGND VPWR VPWR hold251/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold262 hold579/X VGND VGND VPWR VPWR hold578/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 hold240/A VGND VGND VPWR VPWR hold241/A sky130_fd_sc_hd__dlygate4sd3_1
X_7318_ _7318_/A _7318_/B _7318_/C _7318_/D VGND VGND VPWR VPWR _7319_/C sky130_fd_sc_hd__and4_1
XFILLER_123_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8298_ _8302_/A _8306_/B VGND VGND VPWR VPWR _8716_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold273 _5614_/X VGND VGND VPWR VPWR hold274/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold295 hold295/A VGND VGND VPWR VPWR hold296/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 hold284/A VGND VGND VPWR VPWR _9463_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_131_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7249_ _6453_/Y _5756_/X _6365_/Y _7071_/A _7248_/X VGND VGND VPWR VPWR _7252_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_124 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_113 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_146 _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 _6295_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_179 _7052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _8813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4950_ _9440_/Q VGND VGND VPWR VPWR _4950_/Y sky130_fd_sc_hd__clkinv_2
X_4881_ _4953_/A _4933_/A VGND VGND VPWR VPWR _5397_/B sky130_fd_sc_hd__or2_4
XFILLER_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6620_ _9508_/Q VGND VGND VPWR VPWR _6620_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_177_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6551_ _9222_/Q VGND VGND VPWR VPWR _8789_/A sky130_fd_sc_hd__inv_4
XFILLER_20_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5502_ _9433_/Q _5495_/A hold593/X _5495_/Y VGND VGND VPWR VPWR _5502_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6482_ _6482_/A VGND VGND VPWR VPWR _6482_/Y sky130_fd_sc_hd__inv_2
X_9270_ _9800_/CLK _9270_/D _9817_/SET_B VGND VGND VPWR VPWR _9270_/Q sky130_fd_sc_hd__dfstp_1
X_8221_ _8586_/A _8133_/Y _8220_/X VGND VGND VPWR VPWR _8221_/Y sky130_fd_sc_hd__a21oi_1
Xoutput301 _9766_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_2
X_5433_ _9481_/Q _5430_/A hold217/X _5430_/Y VGND VGND VPWR VPWR _9481_/D sky130_fd_sc_hd__a22o_1
X_8152_ _8182_/B VGND VGND VPWR VPWR _8586_/B sky130_fd_sc_hd__clkinv_4
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput312 _9788_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_2
Xoutput323 _9798_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_2
Xoutput334 _9087_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_2
X_5364_ _9528_/Q _5361_/A hold217/A _5361_/Y VGND VGND VPWR VPWR _9528_/D sky130_fd_sc_hd__a22o_1
Xoutput345 _7050_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_2
Xoutput378 _9080_/Q VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_2
Xoutput367 _9070_/Q VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_2
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput356 _9811_/Q VGND VGND VPWR VPWR sram_ro_addr[7] sky130_fd_sc_hd__buf_2
X_7103_ _4877_/Y _7135_/A _4872_/Y _7136_/A _7102_/X VGND VGND VPWR VPWR _7133_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_141_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5295_ _9575_/Q _5291_/X hold577/A _5292_/Y VGND VGND VPWR VPWR _5295_/X sky130_fd_sc_hd__a22o_1
Xoutput389 _9069_/Q VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_2
X_8083_ _8429_/A _8594_/A _8082_/Y VGND VGND VPWR VPWR _8083_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7034_ _4973_/B _4981_/Y _7034_/C _9000_/X VGND VGND VPWR VPWR _7034_/X sky130_fd_sc_hd__and4bb_1
XFILLER_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8985_ hold504/X _9130_/Q _9093_/Q VGND VGND VPWR VPWR _8985_/X sky130_fd_sc_hd__mux2_1
X_7936_ _7936_/A VGND VGND VPWR VPWR _8048_/C sky130_fd_sc_hd__inv_2
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7867_ _7942_/C _8570_/A _8625_/A _7904_/D VGND VGND VPWR VPWR _8366_/A sky130_fd_sc_hd__or4_4
XFILLER_70_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9606_ _9651_/CLK _9606_/D _9689_/SET_B VGND VGND VPWR VPWR _9606_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6818_ _9511_/Q VGND VGND VPWR VPWR _6818_/Y sky130_fd_sc_hd__inv_2
X_7798_ _8277_/A VGND VGND VPWR VPWR _8552_/A sky130_fd_sc_hd__buf_8
XFILLER_50_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9537_ _9576_/CLK _9537_/D _9537_/SET_B VGND VGND VPWR VPWR _9537_/Q sky130_fd_sc_hd__dfstp_1
X_6749_ _9403_/Q VGND VGND VPWR VPWR _6749_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9468_ _9514_/CLK _9468_/D _9571_/SET_B VGND VGND VPWR VPWR _9468_/Q sky130_fd_sc_hd__dfrtp_1
X_8419_ _8625_/C _8419_/B _8419_/C VGND VGND VPWR VPWR _8607_/A sky130_fd_sc_hd__or3_1
XFILLER_109_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9399_ _9831_/CLK _9399_/D _9571_/SET_B VGND VGND VPWR VPWR _9399_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5080_ _7766_/A _7766_/B _8855_/A VGND VGND VPWR VPWR _5085_/B sky130_fd_sc_hd__a21oi_1
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5982_ _9155_/Q _5981_/A hold516/X _5981_/Y VGND VGND VPWR VPWR _9155_/D sky130_fd_sc_hd__a22o_1
X_8770_ _8770_/A VGND VGND VPWR VPWR _8770_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4933_ _4933_/A _4933_/B VGND VGND VPWR VPWR _5301_/B sky130_fd_sc_hd__or2_4
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7721_ _6440_/Y _7509_/A _6435_/Y _7510_/A VGND VGND VPWR VPWR _7721_/X sky130_fd_sc_hd__o22a_1
X_4864_ _9135_/Q VGND VGND VPWR VPWR _4864_/Y sky130_fd_sc_hd__inv_2
XANTENNA_13 _5698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7652_ _4782_/Y _7513_/X _4921_/Y _7514_/X _7651_/X VGND VGND VPWR VPWR _7657_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA_57 _8317_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_24 _6148_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _6711_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7583_ _6461_/Y _7527_/X _6408_/Y _7528_/X VGND VGND VPWR VPWR _7583_/X sky130_fd_sc_hd__o22a_1
X_4795_ _4900_/A _4806_/B VGND VGND VPWR VPWR _5068_/B sky130_fd_sc_hd__or2_4
XANTENNA_35 _6380_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ _6601_/Y _4929_/X _8815_/A _5406_/B VGND VGND VPWR VPWR _6603_/X sky130_fd_sc_hd__o22a_1
XANTENNA_68 _7050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6534_ _9425_/Q VGND VGND VPWR VPWR _6534_/Y sky130_fd_sc_hd__inv_2
X_9322_ _9322_/CLK _9322_/D _9797_/SET_B VGND VGND VPWR VPWR _9322_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9253_ _9695_/CLK _9253_/D _9689_/SET_B VGND VGND VPWR VPWR _9253_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6465_ _9205_/Q VGND VGND VPWR VPWR _6465_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5416_ _9492_/Q _5408_/A hold601/A _5408_/Y VGND VGND VPWR VPWR _5416_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8204_ _8750_/B _8204_/B VGND VGND VPWR VPWR _8206_/A sky130_fd_sc_hd__or2_1
X_6396_ _6391_/Y _5598_/B _6392_/Y _5620_/B _6395_/X VGND VGND VPWR VPWR _6396_/X
+ sky130_fd_sc_hd__o221a_1
X_9184_ _9212_/CLK _9184_/D _9797_/SET_B VGND VGND VPWR VPWR _9184_/Q sky130_fd_sc_hd__dfrtp_1
X_8135_ _8135_/A VGND VGND VPWR VPWR _8762_/A sky130_fd_sc_hd__inv_2
X_5347_ _9539_/Q hold630/X _8964_/A1 _5342_/Y VGND VGND VPWR VPWR _9539_/D sky130_fd_sc_hd__a22o_1
XFILLER_133_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8066_ _8053_/A _8171_/B _8063_/X _8449_/A _8496_/B VGND VGND VPWR VPWR _8066_/X
+ sky130_fd_sc_hd__o2111a_1
X_5278_ _9586_/Q _5276_/A _8964_/A1 _5276_/Y VGND VGND VPWR VPWR _9586_/D sky130_fd_sc_hd__a22o_1
X_7017_ _8853_/A _8851_/A _5969_/X VGND VGND VPWR VPWR _7017_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8968_ _9658_/Q hold510/X _8971_/S VGND VGND VPWR VPWR _8968_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7919_ _8436_/D _8314_/A VGND VGND VPWR VPWR _7920_/A sky130_fd_sc_hd__or2_2
X_8899_ _7604_/Y _9679_/Q _9020_/S VGND VGND VPWR VPWR _8899_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4580_ _6067_/B1 _9799_/Q _4582_/S VGND VGND VPWR VPWR _4581_/A sky130_fd_sc_hd__mux2_1
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR _4928_/A sky130_fd_sc_hd__clkbuf_1
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR _6757_/A sky130_fd_sc_hd__clkbuf_1
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR _6562_/A sky130_fd_sc_hd__clkbuf_1
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR _6934_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR _6118_/A sky130_fd_sc_hd__clkbuf_1
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _8860_/A sky130_fd_sc_hd__buf_6
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _7046_/B sky130_fd_sc_hd__buf_6
XFILLER_155_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput99 sram_ro_data[15] VGND VGND VPWR VPWR _6130_/A sky130_fd_sc_hd__clkbuf_1
X_6250_ _6250_/A VGND VGND VPWR VPWR _6250_/Y sky130_fd_sc_hd__inv_2
X_6181_ _6176_/Y _6180_/A _9085_/Q _6180_/Y VGND VGND VPWR VPWR _9085_/D sky130_fd_sc_hd__o22a_1
X_5201_ _5201_/A _5201_/B VGND VGND VPWR VPWR _5202_/A sky130_fd_sc_hd__or2_4
X_5132_ _9682_/Q _5131_/X _7763_/A _5085_/D VGND VGND VPWR VPWR _9682_/D sky130_fd_sc_hd__o211a_1
XFILLER_97_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5063_ _9015_/X _4572_/B _9721_/Q _5085_/D VGND VGND VPWR VPWR _9721_/D sky130_fd_sc_hd__a22o_1
X_8822_ _8822_/A VGND VGND VPWR VPWR _8822_/X sky130_fd_sc_hd__clkbuf_1
X_5965_ _7874_/C _5965_/B _5965_/C _5964_/X VGND VGND VPWR VPWR _5966_/D sky130_fd_sc_hd__or4b_1
X_8753_ _8158_/A _8666_/X _8158_/B _8667_/Y _8752_/Y VGND VGND VPWR VPWR _8754_/B
+ sky130_fd_sc_hd__o221ai_4
XFILLER_80_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5896_ _5896_/A VGND VGND VPWR VPWR _5896_/Y sky130_fd_sc_hd__inv_2
X_8684_ _8684_/A _8684_/B _8684_/C _8684_/D VGND VGND VPWR VPWR _8773_/A sky130_fd_sc_hd__or4_2
X_4916_ _4912_/Y _5474_/B _4914_/Y _4915_/X VGND VGND VPWR VPWR _4916_/X sky130_fd_sc_hd__o22a_1
X_7704_ _6508_/Y _7507_/A _6646_/Y _7508_/A _7703_/X VGND VGND VPWR VPWR _7711_/A
+ sky130_fd_sc_hd__o221a_1
X_7635_ _6152_/Y _7521_/X _6104_/Y _7522_/X VGND VGND VPWR VPWR _7635_/X sky130_fd_sc_hd__o22a_1
X_4847_ _9601_/Q VGND VGND VPWR VPWR _8849_/A sky130_fd_sc_hd__inv_2
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9305_ _9694_/CLK _9305_/D _9689_/SET_B VGND VGND VPWR VPWR _9305_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7566_ _7731_/A _7525_/X _8803_/A _7526_/X _7565_/X VGND VGND VPWR VPWR _7567_/D
+ sky130_fd_sc_hd__o221a_1
X_4778_ _4808_/A _4832_/A _4774_/Y _4775_/Y _6166_/A VGND VGND VPWR VPWR _4778_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6517_ _9204_/Q VGND VGND VPWR VPWR _6517_/Y sky130_fd_sc_hd__inv_2
X_7497_ _7497_/A VGND VGND VPWR VPWR _7497_/X sky130_fd_sc_hd__buf_4
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9236_ _9651_/CLK _9236_/D _9537_/SET_B VGND VGND VPWR VPWR _9236_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6448_ _9478_/Q VGND VGND VPWR VPWR _6448_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9167_ _9225_/CLK _9167_/D _9731_/SET_B VGND VGND VPWR VPWR _9167_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6379_ _9483_/Q VGND VGND VPWR VPWR _6379_/Y sky130_fd_sc_hd__inv_2
X_8118_ _8118_/A _8479_/B VGND VGND VPWR VPWR _8714_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9098_ _9319_/CLK _9098_/D _9797_/SET_B VGND VGND VPWR VPWR _9098_/Q sky130_fd_sc_hd__dfrtp_4
X_8049_ _8049_/A _8101_/A VGND VGND VPWR VPWR _8049_/X sky130_fd_sc_hd__or2_1
XFILLER_102_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5750_ _7068_/A _7081_/B VGND VGND VPWR VPWR _7108_/C sky130_fd_sc_hd__or2_2
XFILLER_148_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _9086_/Q VGND VGND VPWR VPWR _4701_/Y sky130_fd_sc_hd__inv_2
X_5681_ _5675_/B _5673_/X _5685_/A _5680_/X VGND VGND VPWR VPWR _9321_/D sky130_fd_sc_hd__o2bb2a_1
X_4632_ _4750_/C _4642_/B _4750_/A _4708_/B VGND VGND VPWR VPWR _6189_/B sky130_fd_sc_hd__or4_4
X_7420_ _6392_/Y _7167_/A _6472_/Y _7168_/A VGND VGND VPWR VPWR _7420_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold603 _8881_/X VGND VGND VPWR VPWR hold603/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_4563_ _9107_/Q VGND VGND VPWR VPWR _7763_/A sky130_fd_sc_hd__clkinv_2
XFILLER_128_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7351_ _6963_/Y _7161_/X _6836_/Y _7162_/X VGND VGND VPWR VPWR _7351_/X sky130_fd_sc_hd__o22a_1
Xhold614 _5246_/X VGND VGND VPWR VPWR _9606_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_190_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold636 _5414_/X VGND VGND VPWR VPWR _9494_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6302_ _9567_/Q VGND VGND VPWR VPWR _6302_/Y sky130_fd_sc_hd__clkinv_8
X_7282_ _6227_/Y _7149_/X _6214_/Y _7150_/X _7281_/X VGND VGND VPWR VPWR _7287_/B
+ sky130_fd_sc_hd__o221a_1
X_4494_ _5770_/A VGND VGND VPWR VPWR _6083_/A sky130_fd_sc_hd__buf_12
XFILLER_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold625 hold625/A VGND VGND VPWR VPWR hold625/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold669 _5230_/X VGND VGND VPWR VPWR _9616_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6233_ _9780_/Q VGND VGND VPWR VPWR _6233_/Y sky130_fd_sc_hd__clkinv_4
Xhold647 _4516_/X VGND VGND VPWR VPWR _9825_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold658 _5289_/X VGND VGND VPWR VPWR _9578_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_9021_ _9622_/Q _8785_/A VGND VGND VPWR VPWR _9021_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_170_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6164_ _9387_/Q VGND VGND VPWR VPWR _6164_/Y sky130_fd_sc_hd__clkinv_2
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _9695_/Q _5114_/A hold516/X _5114_/Y VGND VGND VPWR VPWR _5115_/X sky130_fd_sc_hd__a22o_1
X_6095_ _6090_/Y _4865_/X _8849_/B _6196_/A _6094_/X VGND VGND VPWR VPWR _6102_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5046_ _9730_/Q _5038_/A _8975_/A1 _5038_/Y VGND VGND VPWR VPWR _9730_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8805_ _8805_/A VGND VGND VPWR VPWR _8806_/A sky130_fd_sc_hd__clkbuf_1
X_6997_ _6268_/Y _6995_/A _9068_/Q _6995_/Y VGND VGND VPWR VPWR _9068_/D sky130_fd_sc_hd__o22a_1
X_9785_ _9791_/CLK _9785_/D _9821_/SET_B VGND VGND VPWR VPWR _9785_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8736_ _8538_/A _8258_/X _8354_/D _7944_/X VGND VGND VPWR VPWR _8737_/B sky130_fd_sc_hd__o211ai_1
XFILLER_13_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5948_ _5948_/A VGND VGND VPWR VPWR _5948_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8667_ _8667_/A _8667_/B VGND VGND VPWR VPWR _8667_/Y sky130_fd_sc_hd__nor2_1
X_5879_ _9218_/Q _8960_/X _8914_/X _5878_/X VGND VGND VPWR VPWR _9218_/D sky130_fd_sc_hd__o22a_1
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7618_ _6225_/Y _7519_/X _6199_/Y _7520_/X _7617_/X VGND VGND VPWR VPWR _7621_/C
+ sky130_fd_sc_hd__o221a_1
X_8598_ _8643_/D VGND VGND VPWR VPWR _8598_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7549_ _7549_/A _7549_/B _7549_/C _7549_/D VGND VGND VPWR VPWR _7550_/D sky130_fd_sc_hd__and4_1
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9219_ _9225_/CLK _9219_/D _9537_/SET_B VGND VGND VPWR VPWR _9219_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_108_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput201 wb_sel_i[3] VGND VGND VPWR VPWR _7766_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6920_ _9194_/Q VGND VGND VPWR VPWR _6920_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_81_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6851_ _6851_/A VGND VGND VPWR VPWR _6851_/Y sky130_fd_sc_hd__inv_2
X_9570_ _9574_/CLK _9570_/D _9571_/SET_B VGND VGND VPWR VPWR _9570_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5802_ _9270_/Q _5799_/A hold217/A _5799_/Y VGND VGND VPWR VPWR _9270_/D sky130_fd_sc_hd__a22o_1
X_8521_ _8746_/B _8521_/B VGND VGND VPWR VPWR _8523_/A sky130_fd_sc_hd__or2_1
X_6782_ input37/X _8971_/S _6781_/Y _5927_/B VGND VGND VPWR VPWR _6782_/X sky130_fd_sc_hd__o2bb2a_1
X_5733_ _5723_/A _7471_/A _5719_/A _9295_/Q VGND VGND VPWR VPWR _5733_/X sky130_fd_sc_hd__o211a_1
XFILLER_148_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5664_ _9324_/Q _5660_/A _6067_/B1 _5660_/Y VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__a22o_1
X_8452_ _8452_/A VGND VGND VPWR VPWR _8776_/B sky130_fd_sc_hd__inv_2
XFILLER_30_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8383_ _8383_/A _8383_/B _8538_/A VGND VGND VPWR VPWR _8636_/B sky130_fd_sc_hd__nor3_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4615_ _9780_/Q _4613_/A hold510/X _4613_/Y VGND VGND VPWR VPWR _9780_/D sky130_fd_sc_hd__a22o_1
X_5595_ _9371_/Q _5591_/A _6067_/B1 _5591_/Y VGND VGND VPWR VPWR _9371_/D sky130_fd_sc_hd__a22o_1
X_7403_ _6574_/Y _5756_/A _6560_/Y _7061_/A _7402_/X VGND VGND VPWR VPWR _7406_/C
+ sky130_fd_sc_hd__o221a_1
Xhold411 hold411/A VGND VGND VPWR VPWR _5515_/A sky130_fd_sc_hd__clkbuf_2
Xhold400 hold400/A VGND VGND VPWR VPWR _4941_/A sky130_fd_sc_hd__clkbuf_2
X_7334_ _4822_/Y _7173_/X _4807_/Y _7174_/X VGND VGND VPWR VPWR _7334_/X sky130_fd_sc_hd__o22a_1
X_4546_ _4546_/A VGND VGND VPWR VPWR _4547_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_145_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold444 _6058_/X VGND VGND VPWR VPWR _6059_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold433 _5999_/X VGND VGND VPWR VPWR hold434/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 hold422/A VGND VGND VPWR VPWR _9205_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7265_ _7265_/A _7265_/B _7265_/C _7265_/D VGND VGND VPWR VPWR _7275_/B sky130_fd_sc_hd__and4_1
Xhold477 hold477/A VGND VGND VPWR VPWR _9467_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold455 _6067_/X VGND VGND VPWR VPWR hold456/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 hold466/A VGND VGND VPWR VPWR _5660_/A sky130_fd_sc_hd__clkbuf_2
X_4477_ _4476_/Y hold691/X hold470/X VGND VGND VPWR VPWR _4477_/X sky130_fd_sc_hd__a21o_1
X_9004_ _7771_/X _9004_/A1 _9017_/S VGND VGND VPWR VPWR _9004_/X sky130_fd_sc_hd__mux2_1
X_6216_ _6214_/Y _5786_/B _6215_/Y _5826_/B VGND VGND VPWR VPWR _6216_/X sky130_fd_sc_hd__o22a_1
XFILLER_131_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7196_ _6779_/Y _7155_/X _6784_/Y _7156_/X _7195_/X VGND VGND VPWR VPWR _7199_/C
+ sky130_fd_sc_hd__o221a_1
Xhold499 hold499/A VGND VGND VPWR VPWR _9831_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold488 _5664_/X VGND VGND VPWR VPWR _9324_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_112_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6147_ _9827_/Q VGND VGND VPWR VPWR _6147_/Y sky130_fd_sc_hd__inv_6
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6078_ _6078_/A VGND VGND VPWR VPWR _6078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5029_ _5029_/A VGND VGND VPWR VPWR _5030_/S sky130_fd_sc_hd__clkbuf_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9768_ _9817_/CLK _9768_/D _9817_/SET_B VGND VGND VPWR VPWR _9768_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8719_ _8719_/A _8719_/B _8719_/C _8719_/D VGND VGND VPWR VPWR _8773_/D sky130_fd_sc_hd__or4_2
XFILLER_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9699_ _9833_/CLK _9699_/D _9730_/SET_B VGND VGND VPWR VPWR _9699_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5380_ _5380_/A VGND VGND VPWR VPWR _5380_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7050_ _7050_/A VGND VGND VPWR VPWR _7050_/X sky130_fd_sc_hd__buf_6
X_6001_ _9142_/Q _6000_/A hold516/X _6000_/Y VGND VGND VPWR VPWR _6001_/X sky130_fd_sc_hd__a22o_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7952_ _8042_/B _8288_/B _7903_/X _8358_/A _7951_/X VGND VGND VPWR VPWR _7956_/B
+ sky130_fd_sc_hd__o221ai_1
XFILLER_39_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6903_ _9428_/Q VGND VGND VPWR VPWR _6903_/Y sky130_fd_sc_hd__clkinv_2
X_7883_ _8436_/A _8421_/B _8436_/C _8236_/A VGND VGND VPWR VPWR _8347_/A sky130_fd_sc_hd__or4_4
X_9622_ _9730_/CLK _9622_/D _9797_/SET_B VGND VGND VPWR VPWR _9622_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6834_ _6832_/Y _5543_/B _6833_/Y _5628_/B _6189_/X VGND VGND VPWR VPWR _6834_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6765_ _6760_/Y _5389_/B _6761_/Y _5321_/B _6764_/X VGND VGND VPWR VPWR _6772_/C
+ sky130_fd_sc_hd__o221a_1
X_9553_ _9561_/CLK _9553_/D _7042_/B VGND VGND VPWR VPWR _9553_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5716_ _9298_/Q _5708_/A _8975_/A1 _5708_/Y VGND VGND VPWR VPWR _9298_/D sky130_fd_sc_hd__a22o_1
X_9484_ _9491_/CLK _9484_/D _9731_/SET_B VGND VGND VPWR VPWR _9484_/Q sky130_fd_sc_hd__dfstp_1
X_8504_ _7873_/B _8341_/B _7901_/Y _8586_/A _8027_/Y VGND VGND VPWR VPWR _8710_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_148_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8435_ _8435_/A VGND VGND VPWR VPWR _8435_/Y sky130_fd_sc_hd__inv_2
X_6696_ _7380_/A _5658_/B _6695_/Y _5706_/B VGND VGND VPWR VPWR _6696_/X sky130_fd_sc_hd__o22a_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _5847_/A _5647_/B VGND VGND VPWR VPWR _5648_/A sky130_fd_sc_hd__or2_1
XFILLER_148_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5578_ _9382_/Q _5572_/A _8965_/A1 _5572_/Y VGND VGND VPWR VPWR _9382_/D sky130_fd_sc_hd__a22o_1
XFILLER_151_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8366_ _8366_/A _8540_/B VGND VGND VPWR VPWR _8548_/C sky130_fd_sc_hd__nor2_1
Xhold230 _5657_/X VGND VGND VPWR VPWR hold231/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _5370_/X VGND VGND VPWR VPWR hold253/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 hold241/A VGND VGND VPWR VPWR _9380_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7317_ _6121_/Y _7180_/X _6092_/Y _7181_/X _7316_/X VGND VGND VPWR VPWR _7318_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8297_ _8297_/A _8535_/B VGND VGND VPWR VPWR _8299_/A sky130_fd_sc_hd__or2_1
X_4529_ _9818_/Q _4527_/A _6065_/B1 _4527_/Y VGND VGND VPWR VPWR _9818_/D sky130_fd_sc_hd__a22o_1
Xhold274 hold274/A VGND VGND VPWR VPWR hold275/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold578/X VGND VGND VPWR VPWR hold577/A sky130_fd_sc_hd__buf_12
Xhold296 hold296/A VGND VGND VPWR VPWR _9549_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold285 _5575_/X VGND VGND VPWR VPWR hold286/A sky130_fd_sc_hd__dlygate4sd3_1
X_7248_ _7248_/A _7380_/B VGND VGND VPWR VPWR _7248_/X sky130_fd_sc_hd__or2_1
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7179_ _6849_/Y _5756_/X _6944_/Y _7071_/A _7178_/X VGND VGND VPWR VPWR _7186_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_125 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _6400_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_147 _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 _8815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4880_ _9500_/Q VGND VGND VPWR VPWR _4880_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6550_ _8791_/A _5847_/B _8801_/A _5687_/B _6549_/X VGND VGND VPWR VPWR _6557_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5501_ _9434_/Q hold632/X _8965_/A1 _5495_/Y VGND VGND VPWR VPWR _9434_/D sky130_fd_sc_hd__a22o_1
XFILLER_118_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6481_ _6481_/A VGND VGND VPWR VPWR _6481_/Y sky130_fd_sc_hd__clkinv_4
X_8220_ _8421_/B _8473_/A _8219_/X VGND VGND VPWR VPWR _8220_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5432_ _9482_/Q _5430_/A _6065_/B1 _5430_/Y VGND VGND VPWR VPWR _9482_/D sky130_fd_sc_hd__a22o_1
XFILLER_145_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8151_ _8667_/A _8324_/B _8151_/C VGND VGND VPWR VPWR _8750_/B sky130_fd_sc_hd__and3_2
XFILLER_126_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput302 _9767_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_2
Xoutput313 _9789_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_2
Xoutput324 _9799_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_2
Xoutput335 _9088_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_2
X_5363_ _9529_/Q _5361_/A _6065_/B1 _5361_/Y VGND VGND VPWR VPWR _9529_/D sky130_fd_sc_hd__a22o_1
Xoutput346 _7052_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_2
Xoutput368 _9071_/Q VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_113_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput357 _9802_/Q VGND VGND VPWR VPWR sram_ro_clk sky130_fd_sc_hd__buf_2
X_7102_ _4741_/Y _7137_/A _4772_/Y _7138_/A _7101_/X VGND VGND VPWR VPWR _7102_/X
+ sky130_fd_sc_hd__o221a_1
Xoutput379 _9081_/Q VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5294_ _9576_/Q _5292_/A hold510/X _5292_/Y VGND VGND VPWR VPWR _5294_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8082_ _8082_/A _8727_/A VGND VGND VPWR VPWR _8082_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7033_ _7033_/A VGND VGND VPWR VPWR _9101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8984_ _8983_/X hold463/X _9629_/Q VGND VGND VPWR VPWR _8984_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7935_ _7935_/A _8383_/B VGND VGND VPWR VPWR _7935_/X sky130_fd_sc_hd__or2_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7866_ _7866_/A VGND VGND VPWR VPWR _8418_/A sky130_fd_sc_hd__inv_2
XFILLER_63_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9605_ _9651_/CLK _9605_/D _9563_/SET_B VGND VGND VPWR VPWR _9605_/Q sky130_fd_sc_hd__dfrtp_1
X_6817_ _6180_/A _6816_/Y _9080_/Q _6180_/Y VGND VGND VPWR VPWR _9080_/D sky130_fd_sc_hd__o22a_1
XFILLER_168_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7797_ _8436_/A _8421_/B _7875_/B VGND VGND VPWR VPWR _8277_/A sky130_fd_sc_hd__or3_4
X_9536_ _9577_/CLK _9536_/D _9571_/SET_B VGND VGND VPWR VPWR _9536_/Q sky130_fd_sc_hd__dfstp_1
X_6748_ _9538_/Q VGND VGND VPWR VPWR _6748_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_136_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9467_ _9514_/CLK _9467_/D _9571_/SET_B VGND VGND VPWR VPWR _9467_/Q sky130_fd_sc_hd__dfstp_1
X_6679_ _6674_/Y _5786_/B _6675_/Y _5847_/B _6678_/X VGND VGND VPWR VPWR _6680_/C
+ sky130_fd_sc_hd__o221a_1
X_8418_ _8418_/A _8581_/A VGND VGND VPWR VPWR _8422_/B sky130_fd_sc_hd__or2_1
XFILLER_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9398_ _9831_/CLK _9398_/D _9571_/SET_B VGND VGND VPWR VPWR _9398_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_136_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8349_ _8347_/B _8306_/B _8483_/A VGND VGND VPWR VPWR _8352_/B sky130_fd_sc_hd__o21ai_1
XFILLER_124_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5981_ _5981_/A VGND VGND VPWR VPWR _5981_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4932_ _9562_/Q VGND VGND VPWR VPWR _4932_/Y sky130_fd_sc_hd__inv_6
XFILLER_92_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7720_ _6489_/Y _7497_/A _7717_/X _7719_/X VGND VGND VPWR VPWR _7730_/C sky130_fd_sc_hd__o211a_1
XFILLER_178_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7651_ _4681_/Y _7515_/X _4845_/Y _7516_/X VGND VGND VPWR VPWR _7651_/X sky130_fd_sc_hd__o22a_1
X_6602_ _9495_/Q VGND VGND VPWR VPWR _8815_/A sky130_fd_sc_hd__clkinv_8
X_4863_ _6142_/A _4922_/B VGND VGND VPWR VPWR _4863_/X sky130_fd_sc_hd__or2_4
XANTENNA_14 _6127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_25 _6233_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7582_ _6488_/Y _7519_/X _6380_/Y _7520_/X _7581_/X VGND VGND VPWR VPWR _7585_/C
+ sky130_fd_sc_hd__o221a_1
X_4794_ _9709_/Q VGND VGND VPWR VPWR _4794_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_36 _6439_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 _6772_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _8417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6533_ _9276_/Q VGND VGND VPWR VPWR _8797_/A sky130_fd_sc_hd__inv_4
XANTENNA_69 _9161_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9321_ _9322_/CLK _9321_/D _9797_/SET_B VGND VGND VPWR VPWR _9321_/Q sky130_fd_sc_hd__dfrtp_1
X_9252_ _9392_/CLK _9252_/D _9563_/SET_B VGND VGND VPWR VPWR _9252_/Q sky130_fd_sc_hd__dfrtp_1
X_6464_ _6464_/A _6464_/B _6464_/C _6464_/D VGND VGND VPWR VPWR _6505_/B sky130_fd_sc_hd__and4_1
X_5415_ _9493_/Q _5408_/A hold593/A _5408_/Y VGND VGND VPWR VPWR _5415_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8203_ _8203_/A _8412_/A VGND VGND VPWR VPWR _8204_/B sky130_fd_sc_hd__or2_1
X_9183_ _9212_/CLK _9183_/D _9797_/SET_B VGND VGND VPWR VPWR _9183_/Q sky130_fd_sc_hd__dfrtp_1
X_6395_ _6393_/Y _5771_/B _6394_/Y _5581_/B VGND VGND VPWR VPWR _6395_/X sky130_fd_sc_hd__o22a_1
X_8134_ _8134_/A _8134_/B VGND VGND VPWR VPWR _8473_/A sky130_fd_sc_hd__nor2_1
X_5346_ _9540_/Q _5342_/A _8959_/A1 _5342_/Y VGND VGND VPWR VPWR _5346_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8065_ _8065_/A _8178_/B VGND VGND VPWR VPWR _8496_/B sky130_fd_sc_hd__or2_1
XFILLER_87_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5277_ _9587_/Q _5276_/A _6064_/B1 _5276_/Y VGND VGND VPWR VPWR _9587_/D sky130_fd_sc_hd__a22o_1
X_7016_ hold698/X hold710/X _9019_/S VGND VGND VPWR VPWR _7016_/Y sky130_fd_sc_hd__o21ai_4
X_8967_ _9647_/Q hold612/X _8975_/S VGND VGND VPWR VPWR _8967_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7918_ _7918_/A _7918_/B VGND VGND VPWR VPWR _7918_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8898_ _8897_/X _9209_/Q _9096_/Q VGND VGND VPWR VPWR _8898_/X sky130_fd_sc_hd__mux2_1
X_7849_ _8288_/A VGND VGND VPWR VPWR _8383_/A sky130_fd_sc_hd__buf_8
XFILLER_62_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9519_ _9550_/CLK _9519_/D _9537_/SET_B VGND VGND VPWR VPWR _9519_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_156_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _9751_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_46_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR _6825_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_190_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_2
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__buf_2
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR _6655_/A sky130_fd_sc_hd__clkbuf_1
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_4
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_8
XFILLER_10_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__buf_8
XFILLER_170_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5200_ _9636_/Q _5192_/A hold601/X _5192_/Y VGND VGND VPWR VPWR _5200_/X sky130_fd_sc_hd__a22o_1
X_6180_ _6180_/A VGND VGND VPWR VPWR _6180_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5131_ _9103_/Q _9104_/Q _9105_/Q _9107_/D VGND VGND VPWR VPWR _5131_/X sky130_fd_sc_hd__or4_2
XFILLER_69_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5062_ _9016_/X _4572_/B _9722_/Q _5085_/D VGND VGND VPWR VPWR _9722_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8821_ _8821_/A VGND VGND VPWR VPWR _8822_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8752_ _8752_/A VGND VGND VPWR VPWR _8752_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5964_ _7874_/A _7789_/B VGND VGND VPWR VPWR _5964_/X sky130_fd_sc_hd__or2_1
X_7703_ _6643_/Y _7509_/A _6618_/Y _7510_/A VGND VGND VPWR VPWR _7703_/X sky130_fd_sc_hd__o22a_1
X_8683_ _8683_/A _8683_/B _8683_/C _8385_/Y VGND VGND VPWR VPWR _8761_/C sky130_fd_sc_hd__or4b_2
X_5895_ _5895_/A VGND VGND VPWR VPWR _5895_/X sky130_fd_sc_hd__clkbuf_2
X_4915_ _6142_/A _4915_/B VGND VGND VPWR VPWR _4915_/X sky130_fd_sc_hd__or2_4
X_7634_ _6171_/Y _7513_/X _6144_/Y _7514_/X _7633_/X VGND VGND VPWR VPWR _7639_/B
+ sky130_fd_sc_hd__o221a_1
X_4846_ _4883_/A _4913_/A VGND VGND VPWR VPWR _5123_/B sky130_fd_sc_hd__or2_4
XFILLER_165_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7565_ _8825_/A _7527_/X _8801_/A _7528_/X VGND VGND VPWR VPWR _7565_/X sky130_fd_sc_hd__o22a_1
X_6516_ _9357_/Q VGND VGND VPWR VPWR _6516_/Y sky130_fd_sc_hd__clkinv_4
X_9304_ _9391_/CLK _9304_/D _9689_/SET_B VGND VGND VPWR VPWR _9304_/Q sky130_fd_sc_hd__dfrtp_1
X_4777_ _4777_/A VGND VGND VPWR VPWR _6166_/A sky130_fd_sc_hd__buf_6
XFILLER_134_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7496_ _6921_/Y _7491_/X _6952_/Y _7492_/X _7495_/X VGND VGND VPWR VPWR _7532_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9235_ _9830_/CLK _9235_/D _9537_/SET_B VGND VGND VPWR VPWR _9235_/Q sky130_fd_sc_hd__dfrtp_1
X_6447_ _9160_/Q VGND VGND VPWR VPWR _6447_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6378_ _9535_/Q VGND VGND VPWR VPWR _6378_/Y sky130_fd_sc_hd__clkinv_4
X_9166_ _9827_/CLK _9166_/D _9730_/SET_B VGND VGND VPWR VPWR _9166_/Q sky130_fd_sc_hd__dfrtp_1
X_8117_ _8557_/B _8479_/B _8116_/Y VGND VGND VPWR VPWR _8119_/A sky130_fd_sc_hd__o21ai_1
X_5329_ _5378_/A _5329_/B VGND VGND VPWR VPWR _5330_/A sky130_fd_sc_hd__or2_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9097_ _9322_/CLK _9097_/D _9797_/SET_B VGND VGND VPWR VPWR _9097_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_180_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8048_ _8260_/A _8260_/B _8048_/C VGND VGND VPWR VPWR _8101_/A sky130_fd_sc_hd__or3_4
XFILLER_75_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4700_ _5201_/B VGND VGND VPWR VPWR _4700_/Y sky130_fd_sc_hd__inv_4
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _5675_/B _5780_/C _5673_/A _5677_/B VGND VGND VPWR VPWR _5680_/X sky130_fd_sc_hd__o31a_1
XFILLER_175_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4631_ _9768_/Q _4625_/A _6008_/B1 _4625_/Y VGND VGND VPWR VPWR _9768_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7350_ _6833_/Y _7155_/X _6871_/Y _7156_/X _7349_/X VGND VGND VPWR VPWR _7353_/C
+ sky130_fd_sc_hd__o221a_1
X_4562_ _4562_/A VGND VGND VPWR VPWR _9802_/D sky130_fd_sc_hd__clkbuf_1
Xhold604 _5377_/X VGND VGND VPWR VPWR _9518_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold615 _5854_/X VGND VGND VPWR VPWR _9235_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_155_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7281_ _6200_/Y _7151_/X _6199_/Y _7152_/X VGND VGND VPWR VPWR _7281_/X sky130_fd_sc_hd__o22a_1
XFILLER_143_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4493_ _4750_/A _4750_/B _4689_/A _4750_/D VGND VGND VPWR VPWR _4832_/A sky130_fd_sc_hd__or4_4
Xhold626 _4648_/X VGND VGND VPWR VPWR _9761_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6301_ _6301_/A VGND VGND VPWR VPWR _6301_/Y sky130_fd_sc_hd__inv_2
Xhold637 _5189_/X VGND VGND VPWR VPWR _9644_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6232_ _9438_/Q VGND VGND VPWR VPWR _6232_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold648 _4513_/A VGND VGND VPWR VPWR hold648/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold659 _4532_/X VGND VGND VPWR VPWR _9815_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_9020_ _7484_/X _4897_/Y _9020_/S VGND VGND VPWR VPWR _9020_/X sky130_fd_sc_hd__mux2_1
X_6163_ _6163_/A VGND VGND VPWR VPWR _6163_/Y sky130_fd_sc_hd__clkinv_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5114_/A VGND VGND VPWR VPWR _5114_/Y sky130_fd_sc_hd__inv_2
X_6094_ _6092_/Y _5609_/B _6093_/Y _5112_/B VGND VGND VPWR VPWR _6094_/X sky130_fd_sc_hd__o22a_1
Xrepeater410 _7042_/B VGND VGND VPWR VPWR _9817_/SET_B sky130_fd_sc_hd__buf_12
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5045_ _9731_/Q _5038_/A _8969_/A1 _5038_/Y VGND VGND VPWR VPWR _9731_/D sky130_fd_sc_hd__a22o_1
XFILLER_97_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8804_ _8804_/A VGND VGND VPWR VPWR _8804_/X sky130_fd_sc_hd__clkbuf_1
X_6996_ _6176_/Y _6995_/A _9069_/Q _6995_/Y VGND VGND VPWR VPWR _9069_/D sky130_fd_sc_hd__o22a_1
X_9784_ _9791_/CLK _9784_/D _9817_/SET_B VGND VGND VPWR VPWR _9784_/Q sky130_fd_sc_hd__dfstp_1
X_8735_ _8735_/A _8735_/B _8735_/C _7968_/A VGND VGND VPWR VPWR _8738_/B sky130_fd_sc_hd__or4b_1
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5947_ _5947_/A VGND VGND VPWR VPWR _5948_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8666_ _8674_/A _8666_/B VGND VGND VPWR VPWR _8666_/X sky130_fd_sc_hd__and2_1
XFILLER_166_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7617_ _6215_/Y _7521_/X _6191_/Y _7522_/X VGND VGND VPWR VPWR _7617_/X sky130_fd_sc_hd__o22a_1
X_5878_ _5889_/A VGND VGND VPWR VPWR _5878_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_193_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8597_ _8160_/A _8439_/B _8209_/A _8443_/B _8210_/A VGND VGND VPWR VPWR _8673_/B
+ sky130_fd_sc_hd__o221ai_1
X_4829_ _4829_/A VGND VGND VPWR VPWR _4830_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7548_ _6786_/Y _7525_/X _7204_/A _7526_/X _7547_/X VGND VGND VPWR VPWR _7549_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_146_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7479_ _7479_/A _9293_/Q _7479_/C _9297_/Q VGND VGND VPWR VPWR _7528_/A sky130_fd_sc_hd__or4_4
XFILLER_161_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9218_ _9322_/CLK _9218_/D _9797_/SET_B VGND VGND VPWR VPWR _9218_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput202 wb_we_i VGND VGND VPWR VPWR _7766_/A sky130_fd_sc_hd__clkbuf_2
X_9149_ _9734_/CLK _9149_/D _9731_/SET_B VGND VGND VPWR VPWR _9149_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 hold1/A VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dlymetal6s4s_1
XFILLER_39_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6850_ _9459_/Q VGND VGND VPWR VPWR _6850_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6781_ _9177_/Q VGND VGND VPWR VPWR _6781_/Y sky130_fd_sc_hd__clkinv_2
X_5801_ _9271_/Q _5799_/A _6065_/B1 _5799_/Y VGND VGND VPWR VPWR _9271_/D sky130_fd_sc_hd__a22o_1
X_8520_ _8745_/D _8520_/B VGND VGND VPWR VPWR _8521_/B sky130_fd_sc_hd__or2_1
X_5732_ _7471_/A VGND VGND VPWR VPWR _5732_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_1_mgmt_gpio_in[4] clkbuf_1_1_1_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR clkbuf_2_3_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_2
X_5663_ _9325_/Q _5660_/A hold217/X _5660_/Y VGND VGND VPWR VPWR _9325_/D sky130_fd_sc_hd__a22o_1
X_8451_ _8178_/B _8443_/B _8448_/X _8450_/Y VGND VGND VPWR VPWR _8451_/X sky130_fd_sc_hd__o211a_1
X_8382_ _8120_/C _8382_/B _8382_/C _8436_/A VGND VGND VPWR VPWR _8764_/A sky130_fd_sc_hd__and4b_1
XFILLER_135_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5594_ _9372_/Q _5591_/A hold217/A _5591_/Y VGND VGND VPWR VPWR _9372_/D sky130_fd_sc_hd__a22o_1
X_4614_ _9781_/Q _4613_/A hold516/X _4613_/Y VGND VGND VPWR VPWR _9781_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7402_ _7402_/A _7424_/B VGND VGND VPWR VPWR _7402_/X sky130_fd_sc_hd__or2_1
XFILLER_190_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7333_ _4714_/Y _7071_/D _4681_/Y _7166_/X _7332_/X VGND VGND VPWR VPWR _7340_/A
+ sky130_fd_sc_hd__o221a_1
X_4545_ _5201_/A _4545_/B VGND VGND VPWR VPWR _4546_/A sky130_fd_sc_hd__or2_1
Xhold401 _9127_/Q VGND VGND VPWR VPWR hold402/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 hold434/A VGND VGND VPWR VPWR _6000_/A sky130_fd_sc_hd__buf_2
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold423 _5895_/X VGND VGND VPWR VPWR hold424/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _5513_/X VGND VGND VPWR VPWR _5514_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold445 _6189_/B VGND VGND VPWR VPWR _4900_/A sky130_fd_sc_hd__buf_2
X_9003_ _7769_/X _9003_/A1 _9017_/S VGND VGND VPWR VPWR _9003_/X sky130_fd_sc_hd__mux2_1
X_7264_ _6319_/Y _7160_/X _6345_/Y _7071_/B _7263_/X VGND VGND VPWR VPWR _7265_/D
+ sky130_fd_sc_hd__o221a_1
Xhold456 hold456/A VGND VGND VPWR VPWR _9113_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold478 _5901_/X VGND VGND VPWR VPWR _9201_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold467 _5658_/X VGND VGND VPWR VPWR _5659_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4476_ _9629_/Q VGND VGND VPWR VPWR _4476_/Y sky130_fd_sc_hd__inv_2
X_6215_ _9252_/Q VGND VGND VPWR VPWR _6215_/Y sky130_fd_sc_hd__clkinv_2
X_7195_ _6751_/Y _7095_/B _6664_/Y _7157_/X VGND VGND VPWR VPWR _7195_/X sky130_fd_sc_hd__o22a_1
Xhold489 _8980_/X VGND VGND VPWR VPWR hold490/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6146_ _9797_/Q VGND VGND VPWR VPWR _6146_/Y sky130_fd_sc_hd__inv_2
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _6081_/A VGND VGND VPWR VPWR _6078_/A sky130_fd_sc_hd__clkbuf_1
X_5028_ _9133_/Q _6053_/C _9134_/Q _6053_/B VGND VGND VPWR VPWR _5029_/A sky130_fd_sc_hd__or4_1
XFILLER_166_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6979_ _4958_/Y _6180_/A _9078_/Q _6180_/Y VGND VGND VPWR VPWR _9078_/D sky130_fd_sc_hd__o22a_1
X_9767_ _9817_/CLK _9767_/D _9817_/SET_B VGND VGND VPWR VPWR _9767_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8718_ _8718_/A _8718_/B VGND VGND VPWR VPWR _8719_/B sky130_fd_sc_hd__or2_1
X_9698_ _9833_/CLK _9698_/D _9730_/SET_B VGND VGND VPWR VPWR _9698_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8649_ _8649_/A _8649_/B _8649_/C _7949_/X VGND VGND VPWR VPWR _8777_/A sky130_fd_sc_hd__or4b_1
XFILLER_21_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6000_ _6000_/A VGND VGND VPWR VPWR _6000_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7951_ _8280_/A _7903_/X _7948_/X _7949_/X _8496_/A VGND VGND VPWR VPWR _7951_/X
+ sky130_fd_sc_hd__o2111a_1
X_7882_ _8557_/B _7887_/A VGND VGND VPWR VPWR _7970_/A sky130_fd_sc_hd__or2_2
X_6902_ _9441_/Q VGND VGND VPWR VPWR _6902_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9621_ _9730_/CLK _9621_/D _9797_/SET_B VGND VGND VPWR VPWR _9621_/Q sky130_fd_sc_hd__dfrtp_4
X_6833_ _9345_/Q VGND VGND VPWR VPWR _6833_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6764_ _6762_/Y _5990_/B _6763_/Y _5103_/B VGND VGND VPWR VPWR _6764_/X sky130_fd_sc_hd__o22a_1
X_9552_ _9579_/CLK _9552_/D _7042_/B VGND VGND VPWR VPWR _9552_/Q sky130_fd_sc_hd__dfrtp_1
X_5715_ _9299_/Q _5708_/A hold593/X _5708_/Y VGND VGND VPWR VPWR _9299_/D sky130_fd_sc_hd__a22o_1
X_6695_ _9300_/Q VGND VGND VPWR VPWR _6695_/Y sky130_fd_sc_hd__inv_2
X_8503_ _8503_/A _8669_/A VGND VGND VPWR VPWR _8506_/B sky130_fd_sc_hd__or2_1
X_9483_ _9483_/CLK _9483_/D _9727_/SET_B VGND VGND VPWR VPWR _9483_/Q sky130_fd_sc_hd__dfrtp_1
X_5646_ _9336_/Q _5638_/A _8975_/A1 _5638_/Y VGND VGND VPWR VPWR _9336_/D sky130_fd_sc_hd__a22o_1
X_8434_ _8434_/A VGND VGND VPWR VPWR _8750_/A sky130_fd_sc_hd__inv_2
XFILLER_191_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5577_ _9383_/Q _5572_/A _8964_/A1 _5572_/Y VGND VGND VPWR VPWR _9383_/D sky130_fd_sc_hd__a22o_1
Xhold220 hold220/A VGND VGND VPWR VPWR _9512_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_8365_ _8505_/A _8687_/B VGND VGND VPWR VPWR _8641_/C sky130_fd_sc_hd__or2_2
Xhold231 hold231/A VGND VGND VPWR VPWR hold232/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 _9749_/Q VGND VGND VPWR VPWR hold243/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold253/A VGND VGND VPWR VPWR hold254/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7316_ _6135_/Y _7182_/X _6147_/Y _7183_/X VGND VGND VPWR VPWR _7316_/X sky130_fd_sc_hd__o22a_1
X_8296_ _8383_/A _8296_/B VGND VGND VPWR VPWR _8535_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4528_ _9819_/Q _4527_/A _6064_/B1 _4527_/Y VGND VGND VPWR VPWR _9819_/D sky130_fd_sc_hd__a22o_1
Xhold275 hold275/A VGND VGND VPWR VPWR _9359_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold264 _5306_/X VGND VGND VPWR VPWR hold265/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A VGND VGND VPWR VPWR hold287/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7247_ _6487_/Y _7171_/X _6452_/Y _7172_/X _7246_/X VGND VGND VPWR VPWR _7252_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_172_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold297 _6003_/X VGND VGND VPWR VPWR hold298/A sky130_fd_sc_hd__dlygate4sd3_1
X_7178_ _7178_/A _7380_/B VGND VGND VPWR VPWR _7178_/X sky130_fd_sc_hd__or2_1
X_6129_ _9395_/Q VGND VGND VPWR VPWR _6129_/Y sky130_fd_sc_hd__inv_4
XFILLER_100_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_104 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _4784_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _6444_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9819_ _9819_/CLK _9819_/D _7042_/B VGND VGND VPWR VPWR _9819_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5500_ _9435_/Q hold632/X _8964_/A1 _5495_/Y VGND VGND VPWR VPWR _9435_/D sky130_fd_sc_hd__a22o_1
XFILLER_158_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6480_ _9778_/Q VGND VGND VPWR VPWR _6480_/Y sky130_fd_sc_hd__inv_2
X_5431_ _9483_/Q _5430_/A _6064_/B1 _5430_/Y VGND VGND VPWR VPWR _9483_/D sky130_fd_sc_hd__a22o_1
X_8150_ _8264_/C VGND VGND VPWR VPWR _8151_/C sky130_fd_sc_hd__inv_2
XFILLER_114_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput325 _9776_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_2
Xoutput303 _9761_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_2
Xoutput314 _9790_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_2
X_5362_ _9530_/Q _5361_/A _6064_/B1 _5361_/Y VGND VGND VPWR VPWR _9530_/D sky130_fd_sc_hd__a22o_1
Xoutput347 _8859_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_2
XFILLER_160_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput369 _9072_/Q VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_2
X_8081_ _8666_/B _8594_/A VGND VGND VPWR VPWR _8727_/A sky130_fd_sc_hd__nor2_1
Xoutput358 _9803_/Q VGND VGND VPWR VPWR sram_ro_csb sky130_fd_sc_hd__buf_2
Xoutput336 _9089_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_2
X_7101_ _4938_/Y _7139_/A _4936_/Y _7140_/A VGND VGND VPWR VPWR _7101_/X sky130_fd_sc_hd__o22a_1
X_7032_ _9107_/Q _7032_/B VGND VGND VPWR VPWR _7033_/A sky130_fd_sc_hd__or2_1
X_5293_ _9577_/Q _5292_/A hold516/X _5292_/Y VGND VGND VPWR VPWR _5293_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8983_ _9130_/Q _9129_/Q _9093_/Q VGND VGND VPWR VPWR _8983_/X sky130_fd_sc_hd__mux2_1
X_7934_ _8258_/B VGND VGND VPWR VPWR _8383_/B sky130_fd_sc_hd__buf_4
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7865_ _8138_/B _8702_/B _8702_/C VGND VGND VPWR VPWR _7866_/A sky130_fd_sc_hd__or3_1
XFILLER_82_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9604_ _9651_/CLK _9604_/D _9563_/SET_B VGND VGND VPWR VPWR _9604_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7796_ _7996_/B VGND VGND VPWR VPWR _8436_/A sky130_fd_sc_hd__clkbuf_4
X_6816_ _6816_/A _6816_/B _6816_/C VGND VGND VPWR VPWR _6816_/Y sky130_fd_sc_hd__nand3_4
XFILLER_149_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6747_ _6747_/A _6747_/B _6747_/C _6747_/D VGND VGND VPWR VPWR _6815_/A sky130_fd_sc_hd__and4_1
XFILLER_11_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9535_ _9582_/CLK _9535_/D _7042_/B VGND VGND VPWR VPWR _9535_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9466_ _9514_/CLK _9466_/D _9571_/SET_B VGND VGND VPWR VPWR _9466_/Q sky130_fd_sc_hd__dfstp_1
X_6678_ _6676_/Y _5771_/B _6677_/Y _5839_/B VGND VGND VPWR VPWR _6678_/X sky130_fd_sc_hd__o22a_1
X_8417_ _8417_/A _8624_/A _8720_/A _8688_/A VGND VGND VPWR VPWR _8422_/A sky130_fd_sc_hd__or4_1
X_9397_ _9514_/CLK _9397_/D _9571_/SET_B VGND VGND VPWR VPWR _9397_/Q sky130_fd_sc_hd__dfrtp_1
X_5629_ _5629_/A VGND VGND VPWR VPWR _5630_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8348_ _8563_/B _7924_/B _8489_/B _8257_/X _8439_/A VGND VGND VPWR VPWR _8348_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8279_ _8279_/A _8400_/B _8684_/B _8401_/B VGND VGND VPWR VPWR _8283_/A sky130_fd_sc_hd__or4_1
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5980_ _5980_/A VGND VGND VPWR VPWR _5981_/A sky130_fd_sc_hd__clkbuf_4
X_4931_ _9800_/Q VGND VGND VPWR VPWR _4931_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4862_ _4862_/A VGND VGND VPWR VPWR _4862_/Y sky130_fd_sc_hd__clkinv_2
X_7650_ _4743_/Y _7507_/X _4887_/Y _7508_/X _7649_/X VGND VGND VPWR VPWR _7657_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6601_ _6601_/A VGND VGND VPWR VPWR _6601_/Y sky130_fd_sc_hd__inv_2
XANTENNA_26 _6242_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7581_ _6398_/Y _7521_/X _6458_/Y _7522_/X VGND VGND VPWR VPWR _7581_/X sky130_fd_sc_hd__o22a_1
X_4793_ _4808_/A _4933_/B VGND VGND VPWR VPWR _5609_/B sky130_fd_sc_hd__or2_4
XANTENNA_48 _6777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 _6127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9320_ _9322_/CLK _9320_/D _9797_/SET_B VGND VGND VPWR VPWR _9320_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_37 _6439_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_59 _8807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6532_ _6532_/A _6532_/B _6532_/C _6532_/D VGND VGND VPWR VPWR _6660_/A sky130_fd_sc_hd__and4_1
XFILLER_173_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9251_ _9695_/CLK _9251_/D _9563_/SET_B VGND VGND VPWR VPWR _9251_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6463_ _6458_/Y _5340_/B _6459_/Y _5455_/B _6462_/X VGND VGND VPWR VPWR _6464_/D
+ sky130_fd_sc_hd__o221a_1
X_5414_ _9494_/Q _5408_/A _8965_/A1 _5408_/Y VGND VGND VPWR VPWR _5414_/X sky130_fd_sc_hd__a22o_1
X_8202_ _8596_/A _8420_/B VGND VGND VPWR VPWR _8412_/A sky130_fd_sc_hd__nor2_1
X_9182_ _9212_/CLK _9182_/D _9797_/SET_B VGND VGND VPWR VPWR _9182_/Q sky130_fd_sc_hd__dfrtp_1
X_8133_ _8134_/B VGND VGND VPWR VPWR _8133_/Y sky130_fd_sc_hd__inv_2
X_6394_ _9379_/Q VGND VGND VPWR VPWR _6394_/Y sky130_fd_sc_hd__clkinv_2
X_5345_ _9541_/Q _5342_/A hold577/A _5342_/Y VGND VGND VPWR VPWR _5345_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8064_ _8068_/A _8178_/B VGND VGND VPWR VPWR _8449_/A sky130_fd_sc_hd__or2_1
XFILLER_87_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5276_ _5276_/A VGND VGND VPWR VPWR _5276_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7015_ _4958_/Y _7007_/A _9054_/Q _7007_/Y VGND VGND VPWR VPWR _9054_/D sky130_fd_sc_hd__o22a_1
XFILLER_68_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8966_ _9652_/Q _8975_/A1 _8971_/S VGND VGND VPWR VPWR _8966_/X sky130_fd_sc_hd__mux2_1
X_7917_ _7917_/A _8288_/A VGND VGND VPWR VPWR _7918_/B sky130_fd_sc_hd__or2_1
XFILLER_102_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8897_ _7586_/Y _9678_/Q _9020_/S VGND VGND VPWR VPWR _8897_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7848_ _7848_/A VGND VGND VPWR VPWR _8288_/A sky130_fd_sc_hd__buf_4
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7779_ _9110_/Q _7779_/A2 _9109_/Q _7779_/B2 _7778_/X VGND VGND VPWR VPWR _7779_/X
+ sky130_fd_sc_hd__a221o_1
X_9518_ _9550_/CLK _9518_/D _9563_/SET_B VGND VGND VPWR VPWR _9518_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9449_ _9582_/CLK _9449_/D _9727_/SET_B VGND VGND VPWR VPWR _9449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR _6797_/A sky130_fd_sc_hd__clkbuf_1
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR _6552_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_155_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR _6880_/A sky130_fd_sc_hd__clkbuf_1
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR _6442_/A sky130_fd_sc_hd__clkbuf_1
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput79 spi_enabled VGND VGND VPWR VPWR _8875_/S sky130_fd_sc_hd__buf_6
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _8843_/A sky130_fd_sc_hd__buf_8
XFILLER_69_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5130_ _9683_/Q _5125_/A _6008_/B1 _5125_/Y VGND VGND VPWR VPWR _5130_/X sky130_fd_sc_hd__a22o_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5061_ _9017_/X _4572_/B _9723_/Q _5085_/D VGND VGND VPWR VPWR _9723_/D sky130_fd_sc_hd__a22o_1
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8820_ _8820_/A VGND VGND VPWR VPWR _8820_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5963_ _7874_/B VGND VGND VPWR VPWR _7789_/B sky130_fd_sc_hd__inv_2
X_8751_ _8751_/A _8751_/B _8751_/C _8751_/D VGND VGND VPWR VPWR _8780_/A sky130_fd_sc_hd__or4_1
XFILLER_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_opt_4_0_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_4_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4914_ _4914_/A VGND VGND VPWR VPWR _4914_/Y sky130_fd_sc_hd__clkinv_2
X_7702_ _6547_/Y _7497_/A _7699_/X _7701_/X VGND VGND VPWR VPWR _7712_/C sky130_fd_sc_hd__o211a_1
X_8682_ _8682_/A _8682_/B _8682_/C VGND VGND VPWR VPWR _8683_/C sky130_fd_sc_hd__nor3_1
X_5894_ _5990_/A _5894_/B VGND VGND VPWR VPWR _5894_/X sky130_fd_sc_hd__or2_1
XFILLER_52_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7633_ _6129_/Y _7515_/X _6093_/Y _7516_/X VGND VGND VPWR VPWR _7633_/X sky130_fd_sc_hd__o22a_1
X_4845_ _9683_/Q VGND VGND VPWR VPWR _4845_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7564_ _8789_/A _7519_/X _8829_/A _7520_/X _7563_/X VGND VGND VPWR VPWR _7567_/C
+ sky130_fd_sc_hd__o221a_1
X_4776_ _4803_/A _4776_/B VGND VGND VPWR VPWR _4777_/A sky130_fd_sc_hd__or2_1
X_9303_ _9392_/CLK _9303_/D _9689_/SET_B VGND VGND VPWR VPWR _9303_/Q sky130_fd_sc_hd__dfrtp_1
X_6515_ _9352_/Q VGND VGND VPWR VPWR _6515_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7495_ _6941_/Y _7493_/X _6875_/Y _7494_/X VGND VGND VPWR VPWR _7495_/X sky130_fd_sc_hd__o22a_1
X_6446_ _9496_/Q VGND VGND VPWR VPWR _6446_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_173_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9234_ _9830_/CLK _9234_/D _9537_/SET_B VGND VGND VPWR VPWR _9234_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6377_ _9574_/Q VGND VGND VPWR VPWR _6377_/Y sky130_fd_sc_hd__clkinv_4
X_9165_ _9833_/CLK _9165_/D _9730_/SET_B VGND VGND VPWR VPWR _9165_/Q sky130_fd_sc_hd__dfrtp_1
X_8116_ _8627_/B _8116_/B VGND VGND VPWR VPWR _8116_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9096_ _9319_/CLK _9096_/D _9797_/SET_B VGND VGND VPWR VPWR _9096_/Q sky130_fd_sc_hd__dfrtp_4
X_5328_ _9552_/Q _5323_/A _6008_/B1 _5323_/Y VGND VGND VPWR VPWR _9552_/D sky130_fd_sc_hd__a22o_1
X_8047_ _8043_/Y _8608_/B _8105_/C VGND VGND VPWR VPWR _8056_/A sky130_fd_sc_hd__o21a_1
XFILLER_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5259_ _9599_/Q _5257_/A _8964_/A1 _5257_/Y VGND VGND VPWR VPWR _9599_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8949_ _7740_/Y _4971_/A _9093_/Q VGND VGND VPWR VPWR _8949_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _9769_/Q _4625_/A _6067_/B1 _4625_/Y VGND VGND VPWR VPWR _9769_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4561_ _6067_/B1 _9802_/Q _4561_/S VGND VGND VPWR VPWR _4562_/A sky130_fd_sc_hd__mux2_1
X_6300_ _9445_/Q VGND VGND VPWR VPWR _6300_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_183_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold616 _5605_/X VGND VGND VPWR VPWR _9365_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold605 _9629_/Q VGND VGND VPWR VPWR _8987_/S sky130_fd_sc_hd__buf_8
XFILLER_143_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7280_ _6206_/Y _7144_/X _6246_/Y _7145_/X _7279_/X VGND VGND VPWR VPWR _7287_/A
+ sky130_fd_sc_hd__o221a_1
X_4492_ _4642_/B VGND VGND VPWR VPWR _4750_/D sky130_fd_sc_hd__clkinv_2
Xhold627 _4647_/S VGND VGND VPWR VPWR _4645_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xhold638 _5655_/X VGND VGND VPWR VPWR _9330_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6231_ _9490_/Q VGND VGND VPWR VPWR _6231_/Y sky130_fd_sc_hd__clkinv_2
Xhold649 _4511_/X VGND VGND VPWR VPWR _4512_/A sky130_fd_sc_hd__clkdlybuf4s25_1
X_6162_ _6157_/Y _5805_/B _6158_/Y _5979_/B _6161_/X VGND VGND VPWR VPWR _6175_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5113_/A VGND VGND VPWR VPWR _5114_/A sky130_fd_sc_hd__clkbuf_4
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _9695_/Q VGND VGND VPWR VPWR _6093_/Y sky130_fd_sc_hd__inv_2
Xrepeater400 hold601/X VGND VGND VPWR VPWR _6008_/B1 sky130_fd_sc_hd__buf_12
Xrepeater411 _7042_/B VGND VGND VPWR VPWR _9821_/SET_B sky130_fd_sc_hd__buf_12
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _9732_/Q _5038_/A _8965_/A1 _5038_/Y VGND VGND VPWR VPWR _9732_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8803_ _8803_/A VGND VGND VPWR VPWR _8804_/A sky130_fd_sc_hd__clkbuf_1
X_6995_ _6995_/A VGND VGND VPWR VPWR _6995_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9783_ _9791_/CLK _9783_/D _9817_/SET_B VGND VGND VPWR VPWR _9783_/Q sky130_fd_sc_hd__dfstp_1
X_8734_ _8713_/Y _8715_/X _8722_/Y _8724_/X _8733_/Y VGND VGND VPWR VPWR _8734_/Y
+ sky130_fd_sc_hd__o221ai_1
X_5946_ _5990_/A _5946_/B VGND VGND VPWR VPWR _5947_/A sky130_fd_sc_hd__or2_1
X_8665_ _8139_/A _8664_/X _8589_/X VGND VGND VPWR VPWR _8752_/A sky130_fd_sc_hd__o21ai_2
X_5877_ _8960_/X VGND VGND VPWR VPWR _5889_/A sky130_fd_sc_hd__clkinv_4
XFILLER_193_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7616_ _6206_/Y _7513_/X _6190_/Y _7514_/X _7615_/X VGND VGND VPWR VPWR _7621_/B
+ sky130_fd_sc_hd__o221a_1
X_4828_ _9812_/Q _9750_/Q _9668_/Q VGND VGND VPWR VPWR _4829_/A sky130_fd_sc_hd__or3_1
XFILLER_138_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8596_ _8596_/A _8596_/B VGND VGND VPWR VPWR _8751_/A sky130_fd_sc_hd__nor2_1
XFILLER_193_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7547_ _6681_/Y _7527_/X _6664_/Y _7528_/X VGND VGND VPWR VPWR _7547_/X sky130_fd_sc_hd__o22a_1
X_4759_ _4803_/A _4949_/A VGND VGND VPWR VPWR _4760_/A sky130_fd_sc_hd__or2_1
XFILLER_107_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7478_ _7479_/A _9293_/Q _7478_/C _7478_/D VGND VGND VPWR VPWR _7527_/A sky130_fd_sc_hd__or4_4
X_6429_ _9392_/Q VGND VGND VPWR VPWR _6429_/Y sky130_fd_sc_hd__inv_4
XFILLER_146_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9217_ _9322_/CLK _9217_/D _9797_/SET_B VGND VGND VPWR VPWR _9217_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9148_ _9736_/CLK _9148_/D _9731_/SET_B VGND VGND VPWR VPWR _9148_/Q sky130_fd_sc_hd__dfstp_1
X_9079_ _9705_/CLK _9079_/D VGND VGND VPWR VPWR _9079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2 hold2/A VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6780_ _9088_/Q VGND VGND VPWR VPWR _6780_/Y sky130_fd_sc_hd__inv_2
X_5800_ _9272_/Q _5799_/A _6064_/B1 _5799_/Y VGND VGND VPWR VPWR _9272_/D sky130_fd_sc_hd__a22o_1
X_5731_ _9295_/Q VGND VGND VPWR VPWR _7436_/B sky130_fd_sc_hd__inv_2
XFILLER_50_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8450_ _8649_/B _8615_/A VGND VGND VPWR VPWR _8450_/Y sky130_fd_sc_hd__nor2_1
X_5662_ _9326_/Q _5660_/A _6065_/B1 _5660_/Y VGND VGND VPWR VPWR _5662_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8381_ _8693_/A _8714_/C VGND VGND VPWR VPWR _8747_/A sky130_fd_sc_hd__or2_2
XFILLER_136_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4613_ _4613_/A VGND VGND VPWR VPWR _4613_/Y sky130_fd_sc_hd__clkinv_2
X_5593_ _9373_/Q _5591_/A _8964_/A1 _5591_/Y VGND VGND VPWR VPWR _9373_/D sky130_fd_sc_hd__a22o_1
X_7401_ _6547_/Y _7171_/A _6586_/Y _7172_/A _7400_/X VGND VGND VPWR VPWR _7406_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_175_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7332_ _4739_/Y _7167_/X _4719_/Y _7168_/X VGND VGND VPWR VPWR _7332_/X sky130_fd_sc_hd__o22a_1
X_4544_ _4883_/A _6142_/B VGND VGND VPWR VPWR _4545_/B sky130_fd_sc_hd__or2_4
Xhold402 hold402/A VGND VGND VPWR VPWR hold403/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold413 _9718_/Q VGND VGND VPWR VPWR hold414/A sky130_fd_sc_hd__dlygate4sd3_1
X_7263_ _6332_/Y _7161_/X _6294_/Y _7162_/X VGND VGND VPWR VPWR _7263_/X sky130_fd_sc_hd__o22a_1
Xhold435 _5998_/X VGND VGND VPWR VPWR _5999_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold424 hold424/A VGND VGND VPWR VPWR _5896_/A sky130_fd_sc_hd__clkbuf_2
X_9002_ _7767_/X _5083_/X _9002_/S VGND VGND VPWR VPWR _9002_/X sky130_fd_sc_hd__mux2_1
X_6214_ _9279_/Q VGND VGND VPWR VPWR _6214_/Y sky130_fd_sc_hd__inv_2
Xhold457 _5898_/X VGND VGND VPWR VPWR _9204_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold446 _5450_/X VGND VGND VPWR VPWR hold447/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 _8984_/X VGND VGND VPWR VPWR hold469/A sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _4823_/A VGND VGND VPWR VPWR _4682_/C sky130_fd_sc_hd__inv_2
XFILLER_171_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7194_ _6767_/Y _7149_/X _6674_/Y _7150_/X _7193_/X VGND VGND VPWR VPWR _7199_/B
+ sky130_fd_sc_hd__o221a_1
Xhold479 _5252_/X VGND VGND VPWR VPWR hold480/A sky130_fd_sc_hd__dlygate4sd3_1
X_6145_ _9517_/Q VGND VGND VPWR VPWR _6145_/Y sky130_fd_sc_hd__clkinv_2
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6076_/A VGND VGND VPWR VPWR _6076_/X sky130_fd_sc_hd__clkbuf_1
X_5027_ _5027_/A VGND VGND VPWR VPWR _5027_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9766_ _9817_/CLK _9766_/D _9821_/SET_B VGND VGND VPWR VPWR _9766_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6978_ _6180_/A _6977_/Y _9079_/Q _6180_/Y VGND VGND VPWR VPWR _9079_/D sky130_fd_sc_hd__o22a_1
X_8717_ _8717_/A _8717_/B _8717_/C _8717_/D VGND VGND VPWR VPWR _8758_/D sky130_fd_sc_hd__or4_4
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5929_ _5929_/A VGND VGND VPWR VPWR _5929_/Y sky130_fd_sc_hd__inv_2
X_9697_ _9833_/CLK _9697_/D _9730_/SET_B VGND VGND VPWR VPWR _9697_/Q sky130_fd_sc_hd__dfrtp_1
X_8648_ _8714_/B _8648_/B VGND VGND VPWR VPWR _8747_/B sky130_fd_sc_hd__or2_1
XFILLER_139_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8579_ _7873_/A _8341_/B _8102_/C _8578_/Y _8516_/B VGND VGND VPWR VPWR _8659_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7950_ _7953_/A _8281_/B VGND VGND VPWR VPWR _8496_/A sky130_fd_sc_hd__or2_2
XFILLER_54_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7881_ _8702_/B _8538_/A VGND VGND VPWR VPWR _7887_/A sky130_fd_sc_hd__or2_2
X_6901_ _6896_/Y _5367_/B _6897_/Y _5389_/B _6900_/X VGND VGND VPWR VPWR _6908_/C
+ sky130_fd_sc_hd__o221a_1
X_9620_ _9734_/CLK _9620_/D _9731_/SET_B VGND VGND VPWR VPWR _9620_/Q sky130_fd_sc_hd__dfrtp_1
X_6832_ _9402_/Q VGND VGND VPWR VPWR _6832_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_62_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9551_ _9576_/CLK _9551_/D _9537_/SET_B VGND VGND VPWR VPWR _9551_/Q sky130_fd_sc_hd__dfrtp_1
X_6763_ _9698_/Q VGND VGND VPWR VPWR _6763_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5714_ _9300_/Q _5708_/A _8965_/A1 _5708_/Y VGND VGND VPWR VPWR _9300_/D sky130_fd_sc_hd__a22o_1
X_6694_ _9325_/Q VGND VGND VPWR VPWR _7380_/A sky130_fd_sc_hd__clkinv_2
X_8502_ _8502_/A VGND VGND VPWR VPWR _8669_/A sky130_fd_sc_hd__inv_2
X_9482_ _9483_/CLK _9482_/D _9727_/SET_B VGND VGND VPWR VPWR _9482_/Q sky130_fd_sc_hd__dfrtp_1
X_5645_ _9337_/Q _5638_/A _8969_/A1 _5638_/Y VGND VGND VPWR VPWR _9337_/D sky130_fd_sc_hd__a22o_1
X_8433_ _8586_/C VGND VGND VPWR VPWR _8443_/B sky130_fd_sc_hd__clkinv_4
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold210 hold210/A VGND VGND VPWR VPWR _9234_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5576_ _9384_/Q _5572_/A _8959_/A1 _5572_/Y VGND VGND VPWR VPWR _5576_/X sky130_fd_sc_hd__a22o_1
X_8364_ _7901_/Y _8344_/Y _8360_/X _8535_/C _8699_/A VGND VGND VPWR VPWR _8369_/A
+ sky130_fd_sc_hd__a2111o_2
Xhold232 hold232/A VGND VGND VPWR VPWR _9328_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold243 hold243/A VGND VGND VPWR VPWR hold244/A sky130_fd_sc_hd__dlygate4sd3_1
X_7315_ _6103_/Y _5756_/X _6090_/Y _7071_/A _7314_/X VGND VGND VPWR VPWR _7318_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold221 _5452_/X VGND VGND VPWR VPWR hold222/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4527_ _4527_/A VGND VGND VPWR VPWR _4527_/Y sky130_fd_sc_hd__inv_2
X_8295_ _8295_/A _8619_/B VGND VGND VPWR VPWR _8297_/A sky130_fd_sc_hd__or2_1
Xhold265 hold265/A VGND VGND VPWR VPWR hold266/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 hold254/A VGND VGND VPWR VPWR _9525_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold287 hold287/A VGND VGND VPWR VPWR _9385_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold276 _5498_/X VGND VGND VPWR VPWR hold277/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7246_ _6377_/Y _7173_/X _6467_/Y _7174_/X VGND VGND VPWR VPWR _7246_/X sky130_fd_sc_hd__o22a_1
Xhold298 hold298/A VGND VGND VPWR VPWR hold299/A sky130_fd_sc_hd__dlygate4sd3_1
X_7177_ _7424_/B VGND VGND VPWR VPWR _7380_/B sky130_fd_sc_hd__buf_4
X_6128_ _6128_/A VGND VGND VPWR VPWR _6128_/Y sky130_fd_sc_hd__clkinv_2
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6059_/A VGND VGND VPWR VPWR _6059_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_105 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9818_ _9819_/CLK _9818_/D _9817_/SET_B VGND VGND VPWR VPWR _9818_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_149 _4919_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9749_ _4467_/A1 _9749_/D _4986_/X VGND VGND VPWR VPWR _9749_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5430_ _5430_/A VGND VGND VPWR VPWR _5430_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput326 _9777_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_2
Xoutput304 _9768_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_2
Xoutput315 _9791_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_2
X_5361_ _5361_/A VGND VGND VPWR VPWR _5361_/Y sky130_fd_sc_hd__inv_2
Xoutput348 _8860_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_2
XFILLER_141_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5292_ _5292_/A VGND VGND VPWR VPWR _5292_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput359 _9161_/Q VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_2
X_8080_ _8080_/A _8458_/A VGND VGND VPWR VPWR _8082_/A sky130_fd_sc_hd__nand2_1
Xoutput337 _4830_/A VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_2
X_7100_ _7127_/A _7100_/B VGND VGND VPWR VPWR _7140_/A sky130_fd_sc_hd__or2_2
X_7031_ _9098_/Q _5782_/B _7027_/Y _7030_/Y VGND VGND VPWR VPWR _9098_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8982_ _9752_/Q hold341/X _9629_/Q VGND VGND VPWR VPWR _8982_/X sky130_fd_sc_hd__mux2_8
XFILLER_55_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7933_ _8005_/A _7933_/B _7942_/C _8234_/A VGND VGND VPWR VPWR _8258_/B sky130_fd_sc_hd__or4_2
X_7864_ _8216_/A VGND VGND VPWR VPWR _8518_/A sky130_fd_sc_hd__inv_2
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9603_ _9651_/CLK _9603_/D _9563_/SET_B VGND VGND VPWR VPWR _9603_/Q sky130_fd_sc_hd__dfrtp_1
X_7795_ _8421_/D VGND VGND VPWR VPWR _7996_/B sky130_fd_sc_hd__inv_2
X_6815_ _6815_/A _6815_/B _6815_/C _6815_/D VGND VGND VPWR VPWR _6816_/C sky130_fd_sc_hd__and4_1
X_6746_ _6741_/Y _4937_/X _6742_/Y _5282_/B _6745_/X VGND VGND VPWR VPWR _6747_/D
+ sky130_fd_sc_hd__o221a_1
X_9534_ _9812_/CLK _9534_/D _7042_/B VGND VGND VPWR VPWR _9534_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9465_ _9550_/CLK _9465_/D _9571_/SET_B VGND VGND VPWR VPWR _9465_/Q sky130_fd_sc_hd__dfrtp_1
X_6677_ _9242_/Q VGND VGND VPWR VPWR _6677_/Y sky130_fd_sc_hd__inv_2
X_8416_ _8246_/A _8321_/C _8322_/C VGND VGND VPWR VPWR _8688_/A sky130_fd_sc_hd__o21ai_1
X_9396_ _9831_/CLK _9396_/D _9727_/SET_B VGND VGND VPWR VPWR _9396_/Q sky130_fd_sc_hd__dfrtp_1
X_5628_ _5698_/A _5628_/B VGND VGND VPWR VPWR _5629_/A sky130_fd_sc_hd__or2_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5559_ _5570_/A _5559_/B VGND VGND VPWR VPWR _5560_/A sky130_fd_sc_hd__or2_1
X_8347_ _8347_/A _8347_/B VGND VGND VPWR VPWR _8489_/B sky130_fd_sc_hd__or2_1
XFILLER_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8278_ _8278_/A VGND VGND VPWR VPWR _8401_/B sky130_fd_sc_hd__inv_2
X_7229_ _8811_/A _7180_/X _6516_/Y _7181_/X _7228_/X VGND VGND VPWR VPWR _7230_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _9212_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_14_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4930_ _9782_/Q VGND VGND VPWR VPWR _4930_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4861_ _4853_/Y _4854_/X _4855_/Y _5455_/B _4860_/X VGND VGND VPWR VPWR _4886_/A
+ sky130_fd_sc_hd__o221a_1
X_6600_ _9777_/Q VGND VGND VPWR VPWR _6600_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4792_ _9354_/Q VGND VGND VPWR VPWR _4792_/Y sky130_fd_sc_hd__inv_4
X_7580_ _6384_/Y _7513_/X _6446_/Y _7514_/X _7579_/X VGND VGND VPWR VPWR _7585_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA_27 _6244_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 _6127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_38 _6427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6531_ _7402_/A _5658_/B _7733_/A _5935_/B _6530_/X VGND VGND VPWR VPWR _6532_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA_49 _6780_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9250_ _9420_/CLK _9250_/D _9537_/SET_B VGND VGND VPWR VPWR _9250_/Q sky130_fd_sc_hd__dfrtp_1
X_6462_ _6460_/Y _4525_/B _6461_/Y _6058_/B VGND VGND VPWR VPWR _6462_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5413_ _9495_/Q _5408_/A hold42/X _5408_/Y VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__a22o_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6393_ _9286_/Q VGND VGND VPWR VPWR _6393_/Y sky130_fd_sc_hd__inv_2
X_8201_ _8201_/A _8687_/A VGND VGND VPWR VPWR _8203_/A sky130_fd_sc_hd__or2_1
X_9181_ _9212_/CLK _9181_/D _9730_/SET_B VGND VGND VPWR VPWR _9181_/Q sky130_fd_sc_hd__dfrtp_1
X_8132_ _8567_/A _8132_/B _8428_/A VGND VGND VPWR VPWR _8134_/B sky130_fd_sc_hd__or3_1
X_5344_ _9542_/Q _5342_/A hold510/X _5342_/Y VGND VGND VPWR VPWR _5344_/X sky130_fd_sc_hd__a22o_1
X_8063_ _8431_/A _8171_/B _8060_/X _8445_/A _8492_/A VGND VGND VPWR VPWR _8063_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_101_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5275_ _5275_/A VGND VGND VPWR VPWR _5276_/A sky130_fd_sc_hd__clkbuf_2
X_7014_ _6977_/Y _7007_/A _9055_/Q _7007_/Y VGND VGND VPWR VPWR _9055_/D sky130_fd_sc_hd__o22a_1
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8965_ _9654_/Q _8965_/A1 _8971_/S VGND VGND VPWR VPWR _8965_/X sky130_fd_sc_hd__mux2_1
X_7916_ _7957_/A _8274_/B VGND VGND VPWR VPWR _7916_/X sky130_fd_sc_hd__or2_1
X_8896_ _8895_/X _9208_/Q _9096_/Q VGND VGND VPWR VPWR _8896_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7847_ _8421_/D _8421_/B _7875_/B VGND VGND VPWR VPWR _7848_/A sky130_fd_sc_hd__or3_1
XFILLER_62_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7778_ _9108_/Q _7778_/B VGND VGND VPWR VPWR _7778_/X sky130_fd_sc_hd__and2_1
XFILLER_168_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9517_ _9577_/CLK _9517_/D _9571_/SET_B VGND VGND VPWR VPWR _9517_/Q sky130_fd_sc_hd__dfrtp_1
X_6729_ _9120_/Q VGND VGND VPWR VPWR _6729_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_109_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9448_ _9582_/CLK _9448_/D _9727_/SET_B VGND VGND VPWR VPWR _9448_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9379_ _9561_/CLK _9379_/D _7042_/B VGND VGND VPWR VPWR _9379_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _8847_/A sky130_fd_sc_hd__buf_6
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR _6601_/A sky130_fd_sc_hd__clkbuf_1
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR _6276_/A sky130_fd_sc_hd__clkbuf_1
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_4
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__buf_4
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR _4971_/A sky130_fd_sc_hd__buf_12
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5060_ _9091_/Q _5057_/Y _6015_/B _9724_/Q VGND VGND VPWR VPWR _9724_/D sky130_fd_sc_hd__a31o_1
XFILLER_111_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5962_ _7869_/A VGND VGND VPWR VPWR _7874_/A sky130_fd_sc_hd__inv_2
X_8750_ _8750_/A _8750_/B _8750_/C _8750_/D VGND VGND VPWR VPWR _8751_/B sky130_fd_sc_hd__or4_1
XFILLER_80_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4913_ _4913_/A _4913_/B VGND VGND VPWR VPWR _5474_/B sky130_fd_sc_hd__or2_4
XFILLER_18_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7701_ _6510_/Y _7500_/A _6628_/Y _7501_/A _7700_/X VGND VGND VPWR VPWR _7701_/X
+ sky130_fd_sc_hd__o221a_1
X_8681_ _8156_/Y _8432_/B _8637_/C _8398_/A _8614_/C VGND VGND VPWR VPWR _8719_/D
+ sky130_fd_sc_hd__a2111o_1
X_5893_ _8960_/X _7028_/A _5892_/Y _5889_/A _9206_/Q VGND VGND VPWR VPWR _9206_/D
+ sky130_fd_sc_hd__a32o_1
X_7632_ _6153_/Y _7507_/X _6145_/Y _7508_/X _7631_/X VGND VGND VPWR VPWR _7639_/A
+ sky130_fd_sc_hd__o221a_1
X_4844_ _6117_/A _4865_/A VGND VGND VPWR VPWR _4844_/X sky130_fd_sc_hd__or2_4
XFILLER_193_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4775_ _4775_/A VGND VGND VPWR VPWR _4775_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7563_ _8793_/A _7521_/X _8831_/A _7522_/X VGND VGND VPWR VPWR _7563_/X sky130_fd_sc_hd__o22a_1
X_6514_ _9339_/Q VGND VGND VPWR VPWR _8803_/A sky130_fd_sc_hd__inv_4
X_9302_ _9392_/CLK hold77/X _9689_/SET_B VGND VGND VPWR VPWR _9302_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9233_ _9830_/CLK _9233_/D _9537_/SET_B VGND VGND VPWR VPWR _9233_/Q sky130_fd_sc_hd__dfstp_1
X_7494_ _7494_/A VGND VGND VPWR VPWR _7494_/X sky130_fd_sc_hd__buf_4
XFILLER_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6445_ _6440_/Y _5466_/B _6441_/Y _5609_/B _6444_/X VGND VGND VPWR VPWR _6464_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6376_ _6371_/Y _5282_/B _6372_/Y _5274_/B _6375_/X VGND VGND VPWR VPWR _6383_/C
+ sky130_fd_sc_hd__o221a_2
X_9164_ _9833_/CLK _9164_/D _9730_/SET_B VGND VGND VPWR VPWR _9164_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_161_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8115_ _8115_/A _8746_/A VGND VGND VPWR VPWR _8116_/B sky130_fd_sc_hd__or2_1
XFILLER_114_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9095_ _9322_/CLK _9095_/D _9797_/SET_B VGND VGND VPWR VPWR _9095_/Q sky130_fd_sc_hd__dfstp_1
X_5327_ _9553_/Q _5323_/A _6067_/B1 _5323_/Y VGND VGND VPWR VPWR _9553_/D sky130_fd_sc_hd__a22o_1
X_8046_ _8567_/C VGND VGND VPWR VPWR _8105_/C sky130_fd_sc_hd__clkinv_2
XFILLER_102_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5258_ _9600_/Q _5257_/A _6064_/B1 _5257_/Y VGND VGND VPWR VPWR _9600_/D sky130_fd_sc_hd__a22o_1
X_5189_ _9644_/Q _5181_/A _8975_/A1 _5181_/Y VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8948_ _7757_/X _9130_/Q _9093_/Q VGND VGND VPWR VPWR _8948_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8879_ input83/X _8879_/A1 _9628_/Q VGND VGND VPWR VPWR _8879_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4560_ _4560_/A VGND VGND VPWR VPWR _4560_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold617 _5643_/X VGND VGND VPWR VPWR _9339_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold606 _5339_/X VGND VGND VPWR VPWR _9544_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_128_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4491_ _4750_/C VGND VGND VPWR VPWR _4689_/A sky130_fd_sc_hd__clkinv_2
XFILLER_6_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold639 _5649_/A VGND VGND VPWR VPWR hold639/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold628 _4915_/B VGND VGND VPWR VPWR _4939_/A sky130_fd_sc_hd__clkbuf_2
X_6230_ _9594_/Q VGND VGND VPWR VPWR _6230_/Y sky130_fd_sc_hd__inv_6
X_6161_ _6159_/Y _5902_/B _6160_/Y _5068_/B VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__o22a_1
XFILLER_131_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5112_ _5378_/A _5112_/B VGND VGND VPWR VPWR _5113_/A sky130_fd_sc_hd__or2_1
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater401 hold601/X VGND VGND VPWR VPWR _8975_/A1 sky130_fd_sc_hd__buf_12
X_6092_ _9361_/Q VGND VGND VPWR VPWR _6092_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_97_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _9733_/Q _5038_/A _8964_/A1 _5038_/Y VGND VGND VPWR VPWR _9733_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8802_ _8802_/A VGND VGND VPWR VPWR _8802_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6994_ _6994_/A VGND VGND VPWR VPWR _6995_/A sky130_fd_sc_hd__clkbuf_4
X_9782_ _9791_/CLK _9782_/D _9821_/SET_B VGND VGND VPWR VPWR _9782_/Q sky130_fd_sc_hd__dfstp_1
X_5945_ _9167_/Q _5937_/A _8975_/A1 _5937_/Y VGND VGND VPWR VPWR _9167_/D sky130_fd_sc_hd__a22o_1
X_8733_ _8755_/A _8731_/X _8677_/Y _8732_/Y VGND VGND VPWR VPWR _8733_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5876_ _9219_/Q _5868_/A _8975_/A1 _5868_/Y VGND VGND VPWR VPWR _9219_/D sky130_fd_sc_hd__a22o_1
X_8664_ _8011_/A _8157_/B _8666_/B _8439_/A _8437_/B VGND VGND VPWR VPWR _8664_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7615_ _6185_/Y _7515_/X _6188_/Y _7516_/X VGND VGND VPWR VPWR _7615_/X sky130_fd_sc_hd__o22a_1
XFILLER_138_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4827_ _4827_/A _4951_/B VGND VGND VPWR VPWR _5559_/B sky130_fd_sc_hd__or2_4
X_8595_ _8595_/A _8669_/D _8728_/C _8672_/D VGND VGND VPWR VPWR _8601_/A sky130_fd_sc_hd__or4_2
XFILLER_193_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7546_ _6718_/Y _7519_/X _6766_/Y _7520_/X _7545_/X VGND VGND VPWR VPWR _7549_/C
+ sky130_fd_sc_hd__o221a_1
X_4758_ _4758_/A VGND VGND VPWR VPWR _4758_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4689_ _4689_/A _4750_/D _4689_/C _4708_/B VGND VGND VPWR VPWR _4848_/B sky130_fd_sc_hd__or4_4
X_7477_ _7477_/A _7479_/C _9297_/Q VGND VGND VPWR VPWR _7526_/A sky130_fd_sc_hd__or3_4
XFILLER_161_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6428_ _9556_/Q VGND VGND VPWR VPWR _6428_/Y sky130_fd_sc_hd__inv_2
X_9216_ _9319_/CLK _9216_/D _9797_/SET_B VGND VGND VPWR VPWR _9216_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9147_ _9833_/CLK _9147_/D _9730_/SET_B VGND VGND VPWR VPWR _9147_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6359_ _9444_/Q VGND VGND VPWR VPWR _6359_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9078_ _9705_/CLK _9078_/D VGND VGND VPWR VPWR _9078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8029_ _8139_/A _8428_/B VGND VGND VPWR VPWR _8091_/B sky130_fd_sc_hd__or2_2
XFILLER_124_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3 hold3/A VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5730_ _5723_/Y _5729_/X _5719_/A VGND VGND VPWR VPWR _9296_/D sky130_fd_sc_hd__o21a_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5661_ _9327_/Q _5660_/A _6064_/B1 _5660_/Y VGND VGND VPWR VPWR _5661_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7400_ _6637_/Y _7173_/A _6534_/Y _7174_/A VGND VGND VPWR VPWR _7400_/X sky130_fd_sc_hd__o22a_1
X_8380_ _8380_/A VGND VGND VPWR VPWR _8380_/X sky130_fd_sc_hd__clkbuf_1
X_5592_ _9374_/Q _5591_/A _6064_/B1 _5591_/Y VGND VGND VPWR VPWR _9374_/D sky130_fd_sc_hd__a22o_1
X_4612_ _4612_/A VGND VGND VPWR VPWR _4613_/A sky130_fd_sc_hd__buf_2
XFILLER_190_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4543_ _4689_/C _4750_/B _4750_/C _4750_/D VGND VGND VPWR VPWR _6142_/B sky130_fd_sc_hd__or4_4
X_7331_ _7331_/A _7331_/B _7331_/C _7331_/D VGND VGND VPWR VPWR _7341_/B sky130_fd_sc_hd__and4_1
X_7262_ _6327_/Y _7155_/X _6341_/Y _7156_/X _7261_/X VGND VGND VPWR VPWR _7265_/C
+ sky130_fd_sc_hd__o221a_1
Xhold414 hold414/A VGND VGND VPWR VPWR hold415/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 _5894_/X VGND VGND VPWR VPWR _5895_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold436 _4865_/X VGND VGND VPWR VPWR _5998_/B sky130_fd_sc_hd__clkbuf_2
Xhold403 hold403/A VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_6213_ _9266_/Q VGND VGND VPWR VPWR _6213_/Y sky130_fd_sc_hd__inv_2
Xhold447 hold447/A VGND VGND VPWR VPWR hold448/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 _5661_/X VGND VGND VPWR VPWR hold459/A sky130_fd_sc_hd__dlygate4sd3_1
X_4474_ _5770_/A VGND VGND VPWR VPWR _5201_/A sky130_fd_sc_hd__buf_6
Xhold469 hold469/A VGND VGND VPWR VPWR hold470/A sky130_fd_sc_hd__dlygate4sd3_1
X_9001_ _7134_/X _4897_/Y _9001_/S VGND VGND VPWR VPWR _9001_/X sky130_fd_sc_hd__mux2_1
X_7193_ _6791_/Y _7151_/X _6766_/Y _7152_/X VGND VGND VPWR VPWR _7193_/X sky130_fd_sc_hd__o22a_1
X_6144_ _9499_/Q VGND VGND VPWR VPWR _6144_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6075_ _6081_/A VGND VGND VPWR VPWR _6076_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5026_ _6017_/A VGND VGND VPWR VPWR _5027_/A sky130_fd_sc_hd__clkbuf_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _6977_/A _6977_/B _6977_/C VGND VGND VPWR VPWR _6977_/Y sky130_fd_sc_hd__nand3_4
X_9765_ _9817_/CLK _9765_/D _9817_/SET_B VGND VGND VPWR VPWR _9765_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5928_ _5928_/A VGND VGND VPWR VPWR _5929_/A sky130_fd_sc_hd__clkbuf_2
X_8716_ _8716_/A _8716_/B VGND VGND VPWR VPWR _8717_/B sky130_fd_sc_hd__or2_1
XFILLER_41_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9696_ _9833_/CLK _9696_/D _9730_/SET_B VGND VGND VPWR VPWR _9696_/Q sky130_fd_sc_hd__dfrtp_1
X_8647_ _8647_/A _8647_/B VGND VGND VPWR VPWR _8749_/B sky130_fd_sc_hd__or2_1
X_5859_ _5859_/A VGND VGND VPWR VPWR _5860_/A sky130_fd_sc_hd__clkbuf_2
X_8578_ _8578_/A VGND VGND VPWR VPWR _8578_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7529_ _6854_/Y _7527_/X _6957_/Y _7528_/X VGND VGND VPWR VPWR _7529_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7880_ _8489_/A VGND VGND VPWR VPWR _8538_/A sky130_fd_sc_hd__buf_4
XFILLER_94_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6900_ _6898_/Y _5466_/B _6899_/Y _5274_/B VGND VGND VPWR VPWR _6900_/X sky130_fd_sc_hd__o22a_1
X_6831_ _9157_/Q VGND VGND VPWR VPWR _6831_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9550_ _9550_/CLK _9550_/D _9537_/SET_B VGND VGND VPWR VPWR _9550_/Q sky130_fd_sc_hd__dfrtp_1
X_8501_ _8501_/A _8776_/C _8501_/C _8656_/C VGND VGND VPWR VPWR _8506_/A sky130_fd_sc_hd__or4_1
X_6762_ _9145_/Q VGND VGND VPWR VPWR _6762_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5713_ _9301_/Q _5708_/A hold42/X _5708_/Y VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__a22o_1
XFILLER_148_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6693_ _9377_/Q VGND VGND VPWR VPWR _6693_/Y sky130_fd_sc_hd__inv_2
X_9481_ _9483_/CLK _9481_/D _9727_/SET_B VGND VGND VPWR VPWR _9481_/Q sky130_fd_sc_hd__dfstp_1
X_5644_ _9338_/Q _5638_/A hold136/X _5638_/Y VGND VGND VPWR VPWR _5644_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8432_ _8560_/B _8432_/B VGND VGND VPWR VPWR _8586_/C sky130_fd_sc_hd__or2_1
XFILLER_31_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8363_ _8503_/A _8716_/B VGND VGND VPWR VPWR _8699_/A sky130_fd_sc_hd__or2_1
Xhold200 _5247_/X VGND VGND VPWR VPWR hold201/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 _5311_/X VGND VGND VPWR VPWR hold212/A sky130_fd_sc_hd__dlygate4sd3_1
X_5575_ _9385_/Q _5572_/A hold577/A _5572_/Y VGND VGND VPWR VPWR _5575_/X sky130_fd_sc_hd__a22o_1
XFILLER_156_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7314_ _7314_/A _7380_/B VGND VGND VPWR VPWR _7314_/X sky130_fd_sc_hd__or2_1
Xhold233 _5619_/X VGND VGND VPWR VPWR hold234/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 hold244/A VGND VGND VPWR VPWR hold245/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 hold222/A VGND VGND VPWR VPWR hold223/A sky130_fd_sc_hd__dlygate4sd3_1
X_8294_ _8361_/A _8302_/B VGND VGND VPWR VPWR _8619_/B sky130_fd_sc_hd__nor2_1
X_4526_ _4526_/A VGND VGND VPWR VPWR _4527_/A sky130_fd_sc_hd__clkbuf_2
Xhold266 hold266/A VGND VGND VPWR VPWR _9567_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold277 hold277/A VGND VGND VPWR VPWR hold278/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold255 _5300_/X VGND VGND VPWR VPWR hold256/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7245_ _6488_/Y _7071_/D _6429_/Y _7166_/X _7244_/X VGND VGND VPWR VPWR _7252_/A
+ sky130_fd_sc_hd__o221a_1
Xhold288 _5711_/X VGND VGND VPWR VPWR hold289/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold299 hold299/A VGND VGND VPWR VPWR _9140_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7176_ _6950_/Y _7171_/X _6890_/Y _7172_/X _7175_/X VGND VGND VPWR VPWR _7186_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6127_ _6127_/A _6127_/B _6127_/C _6127_/D VGND VGND VPWR VPWR _6176_/B sky130_fd_sc_hd__and4_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6083_/A _6058_/B VGND VGND VPWR VPWR _6058_/X sky130_fd_sc_hd__or2_1
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_106 _5998_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5009_ _5017_/A VGND VGND VPWR VPWR _5010_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_139 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_128 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9817_ _9817_/CLK _9817_/D _9817_/SET_B VGND VGND VPWR VPWR _9817_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9748_ _4467_/A1 _9748_/D _4992_/X VGND VGND VPWR VPWR _9748_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9679_ _9679_/CLK _9679_/D _9730_/SET_B VGND VGND VPWR VPWR _9679_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput305 _9769_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_2
Xoutput316 _9792_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_2
X_5360_ _5360_/A VGND VGND VPWR VPWR _5361_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5291_ _5291_/A VGND VGND VPWR VPWR _5291_/X sky130_fd_sc_hd__clkbuf_4
Xoutput338 _8844_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_2
Xoutput327 _9778_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_2
Xoutput349 _9804_/Q VGND VGND VPWR VPWR sram_ro_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_141_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7030_ _7030_/A VGND VGND VPWR VPWR _7030_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8981_ hold491/X hold385/X _8987_/S VGND VGND VPWR VPWR _8981_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7932_ _8042_/B _8274_/B _8483_/A _7931_/X VGND VGND VPWR VPWR _7932_/X sky130_fd_sc_hd__o211a_1
XFILLER_55_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7863_ _8557_/A _8314_/A VGND VGND VPWR VPWR _8216_/A sky130_fd_sc_hd__or2_1
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7794_ _8341_/A _8324_/C _7873_/A VGND VGND VPWR VPWR _8678_/A sky130_fd_sc_hd__and3_2
XFILLER_90_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6814_ _6814_/A _6814_/B _6814_/C _6814_/D VGND VGND VPWR VPWR _6815_/D sky130_fd_sc_hd__and4_1
XFILLER_23_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9602_ _9686_/CLK _9602_/D _7042_/B VGND VGND VPWR VPWR _9602_/Q sky130_fd_sc_hd__dfrtp_1
X_6745_ _6743_/Y _5397_/B _6744_/Y _5406_/B VGND VGND VPWR VPWR _6745_/X sky130_fd_sc_hd__o22a_1
XFILLER_23_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9533_ _9582_/CLK _9533_/D _7042_/B VGND VGND VPWR VPWR _9533_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_51_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9464_ _9516_/CLK _9464_/D _9571_/SET_B VGND VGND VPWR VPWR _9464_/Q sky130_fd_sc_hd__dfrtp_1
X_8415_ _8415_/A _8735_/B VGND VGND VPWR VPWR _8624_/A sky130_fd_sc_hd__or2_2
XFILLER_109_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6676_ _9284_/Q VGND VGND VPWR VPWR _6676_/Y sky130_fd_sc_hd__clkinv_2
X_9395_ _9694_/CLK _9395_/D _9689_/SET_B VGND VGND VPWR VPWR _9395_/Q sky130_fd_sc_hd__dfrtp_1
X_5627_ _9349_/Q _5622_/A _8975_/A1 _5622_/Y VGND VGND VPWR VPWR _9349_/D sky130_fd_sc_hd__a22o_1
X_8346_ _8493_/A _8684_/B VGND VGND VPWR VPWR _8346_/Y sky130_fd_sc_hd__nor2_2
X_5558_ _9396_/Q _5553_/A _6008_/B1 _5553_/Y VGND VGND VPWR VPWR _9396_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8277_ _8277_/A _8281_/B VGND VGND VPWR VPWR _8278_/A sky130_fd_sc_hd__or2_1
X_4509_ _4750_/C _4642_/B _4689_/C _4708_/B VGND VGND VPWR VPWR _4827_/A sky130_fd_sc_hd__or4_4
X_7228_ _8825_/A _7182_/X _8823_/A _7183_/X VGND VGND VPWR VPWR _7228_/X sky130_fd_sc_hd__o22a_1
X_5489_ _9443_/Q _5484_/A _6065_/B1 _5484_/Y VGND VGND VPWR VPWR _9443_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7159_ _6945_/Y _7155_/X _6936_/Y _7156_/X _7158_/X VGND VGND VPWR VPWR _7165_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4860_ _4857_/Y _4502_/B _4858_/Y _5255_/B VGND VGND VPWR VPWR _4860_/X sky130_fd_sc_hd__o22a_1
XFILLER_82_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_17 _6127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _6427_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _6528_/Y _5771_/B _6529_/Y _5839_/B VGND VGND VPWR VPWR _6530_/X sky130_fd_sc_hd__o22a_1
XANTENNA_28 _6246_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4791_ _4827_/A _4865_/B VGND VGND VPWR VPWR _5112_/B sky130_fd_sc_hd__or2_4
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6461_ _9116_/Q VGND VGND VPWR VPWR _6461_/Y sky130_fd_sc_hd__clkinv_2
X_5412_ _9496_/Q _5408_/A hold53/X _5408_/Y VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__a22o_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6392_ _9353_/Q VGND VGND VPWR VPWR _6392_/Y sky130_fd_sc_hd__clkinv_2
X_8200_ _8596_/A _8682_/B VGND VGND VPWR VPWR _8687_/A sky130_fd_sc_hd__nor2_1
X_9180_ _9319_/CLK _9180_/D _9797_/SET_B VGND VGND VPWR VPWR _9180_/Q sky130_fd_sc_hd__dfrtp_1
X_8131_ _8260_/A _8137_/B _8008_/A _8161_/A VGND VGND VPWR VPWR _8428_/A sky130_fd_sc_hd__or4bb_4
X_5343_ _9543_/Q _5342_/A hold516/X _5342_/Y VGND VGND VPWR VPWR _5343_/X sky130_fd_sc_hd__a22o_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8062_ _8065_/A _8171_/B VGND VGND VPWR VPWR _8492_/A sky130_fd_sc_hd__or2_1
X_5274_ _5282_/A _5274_/B VGND VGND VPWR VPWR _5275_/A sky130_fd_sc_hd__or2_1
X_7013_ _6816_/Y _7007_/A _9056_/Q _7007_/Y VGND VGND VPWR VPWR _9056_/D sky130_fd_sc_hd__o22a_1
XFILLER_114_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8964_ _9655_/Q _8964_/A1 _8971_/S VGND VGND VPWR VPWR _8964_/X sky130_fd_sc_hd__mux2_1
X_7915_ _8268_/C _8272_/A VGND VGND VPWR VPWR _8274_/B sky130_fd_sc_hd__or2_2
X_8895_ _7568_/Y _9677_/Q _9020_/S VGND VGND VPWR VPWR _8895_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7846_ _7846_/A VGND VGND VPWR VPWR _8243_/A sky130_fd_sc_hd__buf_4
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7777_ _9110_/Q _7777_/A2 _9109_/Q _7777_/B2 _7776_/X VGND VGND VPWR VPWR _7777_/X
+ sky130_fd_sc_hd__a221o_1
X_4989_ _4989_/A VGND VGND VPWR VPWR _4989_/Y sky130_fd_sc_hd__clkinv_2
X_9516_ _9516_/CLK _9516_/D _9571_/SET_B VGND VGND VPWR VPWR _9516_/Q sky130_fd_sc_hd__dfrtp_1
X_6728_ _6723_/Y _4511_/B _6724_/Y _5570_/B _6727_/X VGND VGND VPWR VPWR _6747_/A
+ sky130_fd_sc_hd__o221a_1
X_9447_ _9686_/CLK _9447_/D _9817_/SET_B VGND VGND VPWR VPWR _9447_/Q sky130_fd_sc_hd__dfrtp_1
X_6070__1 _8879_/A1 VGND VGND VPWR VPWR _9100_/CLK sky130_fd_sc_hd__inv_4
X_6659_ _6659_/A _6659_/B _6659_/C _6659_/D VGND VGND VPWR VPWR _6660_/D sky130_fd_sc_hd__and4_2
XFILLER_191_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9378_ _9561_/CLK _9378_/D _7042_/B VGND VGND VPWR VPWR _9378_/Q sky130_fd_sc_hd__dfrtp_1
X_8329_ _8755_/A _8329_/B VGND VGND VPWR VPWR _8329_/X sky130_fd_sc_hd__or2_1
XFILLER_152_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_2
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR _6844_/A sky130_fd_sc_hd__clkbuf_1
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR _6737_/A sky130_fd_sc_hd__clkbuf_1
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR _6481_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR _6224_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_155_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5961_ _5961_/A _5961_/B input164/X VGND VGND VPWR VPWR _5965_/C sky130_fd_sc_hd__or3b_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8680_ _8763_/B VGND VGND VPWR VPWR _8680_/Y sky130_fd_sc_hd__inv_2
X_7700_ _6637_/Y _7502_/A _6635_/Y _7503_/A VGND VGND VPWR VPWR _7700_/X sky130_fd_sc_hd__o22a_1
X_4912_ _9448_/Q VGND VGND VPWR VPWR _4912_/Y sky130_fd_sc_hd__clkinv_2
X_7631_ _6105_/Y _7509_/X _6121_/Y _7510_/X VGND VGND VPWR VPWR _7631_/X sky130_fd_sc_hd__o22a_1
X_5892_ _9020_/X VGND VGND VPWR VPWR _5892_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4843_ _4843_/A VGND VGND VPWR VPWR _4843_/Y sky130_fd_sc_hd__inv_2
X_7562_ _8791_/A _7513_/X _8815_/A _7514_/X _7561_/X VGND VGND VPWR VPWR _7567_/B
+ sky130_fd_sc_hd__o221a_1
X_4774_ _9831_/Q VGND VGND VPWR VPWR _4774_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9301_ _9392_/CLK hold95/X _9689_/SET_B VGND VGND VPWR VPWR _9301_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_119_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6513_ _6508_/Y _5797_/B _8799_/A _5706_/B _6512_/X VGND VGND VPWR VPWR _6532_/A
+ sky130_fd_sc_hd__o221a_1
X_7493_ _7493_/A VGND VGND VPWR VPWR _7493_/X sky130_fd_sc_hd__buf_4
X_9232_ _9830_/CLK _9232_/D _9537_/SET_B VGND VGND VPWR VPWR _9232_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6444_ _6442_/Y _4844_/X _6443_/Y _5255_/B VGND VGND VPWR VPWR _6444_/X sky130_fd_sc_hd__o22a_4
XFILLER_106_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6375_ _6373_/Y _4634_/B _6374_/Y _5589_/B VGND VGND VPWR VPWR _6375_/X sky130_fd_sc_hd__o22a_1
X_9163_ _9833_/CLK _9163_/D _9730_/SET_B VGND VGND VPWR VPWR _9163_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8114_ _8755_/A _8582_/A VGND VGND VPWR VPWR _8746_/A sky130_fd_sc_hd__or2_1
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9094_ _8879_/A1 _9094_/D _6074_/X VGND VGND VPWR VPWR _9094_/Q sky130_fd_sc_hd__dfrtp_2
X_5326_ _9554_/Q _5323_/A hold217/X _5323_/Y VGND VGND VPWR VPWR _9554_/D sky130_fd_sc_hd__a22o_1
X_8045_ _8045_/A VGND VGND VPWR VPWR _8608_/B sky130_fd_sc_hd__inv_2
XFILLER_114_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5257_ _5257_/A VGND VGND VPWR VPWR _5257_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5188_ _9645_/Q _5181_/A hold593/X _5181_/Y VGND VGND VPWR VPWR _9645_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8947_ _7752_/X _9128_/Q _9093_/Q VGND VGND VPWR VPWR _8947_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8878_ input84/X hold23/A _9668_/Q VGND VGND VPWR VPWR _8878_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7829_ _7904_/D _7827_/B _7828_/B VGND VGND VPWR VPWR _8580_/B sky130_fd_sc_hd__a21o_2
XFILLER_157_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold607 _5569_/X VGND VGND VPWR VPWR _9388_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold618 _5298_/X VGND VGND VPWR VPWR _9572_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_4490_ _4803_/A VGND VGND VPWR VPWR _4808_/A sky130_fd_sc_hd__clkbuf_4
Xhold629 _5346_/X VGND VGND VPWR VPWR _9540_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6160_ _9716_/Q VGND VGND VPWR VPWR _6160_/Y sky130_fd_sc_hd__inv_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5770_/A VGND VGND VPWR VPWR _5378_/A sky130_fd_sc_hd__buf_8
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater402 _9730_/SET_B VGND VGND VPWR VPWR _9731_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6091_ _6091_/A VGND VGND VPWR VPWR _8849_/B sky130_fd_sc_hd__clkinv_4
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _9734_/Q _5038_/A _8959_/A1 _5038_/Y VGND VGND VPWR VPWR _9734_/D sky130_fd_sc_hd__a22o_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8801_ _8801_/A VGND VGND VPWR VPWR _8802_/A sky130_fd_sc_hd__clkbuf_1
X_6993_ _7005_/B _6993_/B VGND VGND VPWR VPWR _6994_/A sky130_fd_sc_hd__or2_4
X_9781_ _9819_/CLK _9781_/D _9821_/SET_B VGND VGND VPWR VPWR _9781_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8732_ _8756_/C VGND VGND VPWR VPWR _8732_/Y sky130_fd_sc_hd__inv_2
X_5944_ _9168_/Q _5937_/A _8969_/A1 _5937_/Y VGND VGND VPWR VPWR _9168_/D sky130_fd_sc_hd__a22o_1
XFILLER_159_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5875_ _9220_/Q _5868_/A _8969_/A1 _5868_/Y VGND VGND VPWR VPWR _9220_/D sky130_fd_sc_hd__a22o_1
X_8663_ _8755_/D VGND VGND VPWR VPWR _8663_/Y sky130_fd_sc_hd__inv_2
X_4826_ _9388_/Q VGND VGND VPWR VPWR _4826_/Y sky130_fd_sc_hd__inv_6
X_7614_ _6214_/Y _7507_/X _6226_/Y _7508_/X _7613_/X VGND VGND VPWR VPWR _7621_/A
+ sky130_fd_sc_hd__o221a_1
X_8594_ _8594_/A _8596_/B VGND VGND VPWR VPWR _8672_/D sky130_fd_sc_hd__nor2_1
XFILLER_138_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7545_ _6668_/Y _7521_/X _6748_/Y _7522_/X VGND VGND VPWR VPWR _7545_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4757_ _4753_/Y _5647_/B _4755_/Y _5826_/B VGND VGND VPWR VPWR _4757_/X sky130_fd_sc_hd__o22a_1
X_4688_ _9193_/Q VGND VGND VPWR VPWR _4688_/Y sky130_fd_sc_hd__inv_2
X_7476_ _7477_/A _7476_/B _9297_/Q VGND VGND VPWR VPWR _7525_/A sky130_fd_sc_hd__or3_4
X_6427_ _9522_/Q VGND VGND VPWR VPWR _6427_/Y sky130_fd_sc_hd__inv_4
XFILLER_107_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9215_ _9322_/CLK _9215_/D _9797_/SET_B VGND VGND VPWR VPWR _9215_/Q sky130_fd_sc_hd__dfrtp_1
X_6358_ _6180_/A _6357_/Y _9083_/Q _6180_/Y VGND VGND VPWR VPWR _9083_/D sky130_fd_sc_hd__o22a_1
X_9146_ _9833_/CLK _9146_/D _9730_/SET_B VGND VGND VPWR VPWR _9146_/Q sky130_fd_sc_hd__dfrtp_1
X_5309_ _9564_/Q _5303_/A hold136/X _5303_/Y VGND VGND VPWR VPWR _5309_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9077_ _9705_/CLK _9077_/D VGND VGND VPWR VPWR _9077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6289_ _9779_/Q VGND VGND VPWR VPWR _6289_/Y sky130_fd_sc_hd__inv_2
X_8028_ _8028_/A _8132_/B VGND VGND VPWR VPWR _8428_/B sky130_fd_sc_hd__or2b_1
XFILLER_124_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9695_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold4 hold4/A VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xnet399_2 net399_3/A VGND VGND VPWR VPWR _7053_/A sky130_fd_sc_hd__inv_4
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5660_ _5660_/A VGND VGND VPWR VPWR _5660_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4611_ _5201_/A _4611_/B VGND VGND VPWR VPWR _4612_/A sky130_fd_sc_hd__or2_1
X_5591_ _5591_/A VGND VGND VPWR VPWR _5591_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4542_ _4542_/A VGND VGND VPWR VPWR _9812_/D sky130_fd_sc_hd__clkbuf_1
X_7330_ _4705_/Y _7160_/X _4845_/Y _7071_/B _7329_/X VGND VGND VPWR VPWR _7331_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7261_ _6295_/Y _7095_/B _6347_/Y _7157_/X VGND VGND VPWR VPWR _7261_/X sky130_fd_sc_hd__o22a_1
XFILLER_128_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold415 hold415/A VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4473_ _4473_/A VGND VGND VPWR VPWR _5770_/A sky130_fd_sc_hd__inv_6
Xhold426 _4715_/X VGND VGND VPWR VPWR _5894_/B sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold404 _8978_/X VGND VGND VPWR VPWR hold404/X sky130_fd_sc_hd__clkbuf_2
X_6212_ _9342_/Q VGND VGND VPWR VPWR _7292_/A sky130_fd_sc_hd__inv_2
XFILLER_131_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold448 hold448/A VGND VGND VPWR VPWR _9470_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold459 hold459/A VGND VGND VPWR VPWR hold460/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 _4865_/A VGND VGND VPWR VPWR _4951_/A sky130_fd_sc_hd__clkbuf_2
X_9000_ _9132_/Q _9134_/Q _9133_/Q VGND VGND VPWR VPWR _9000_/X sky130_fd_sc_hd__mux2_1
X_7192_ _6675_/Y _7144_/X _6712_/Y _7145_/X _7191_/X VGND VGND VPWR VPWR _7199_/A
+ sky130_fd_sc_hd__o221a_1
X_6143_ _6140_/Y _4869_/X _6141_/Y _5329_/B _6142_/X VGND VGND VPWR VPWR _6150_/C
+ sky130_fd_sc_hd__o221a_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6074_ _6074_/A VGND VGND VPWR VPWR _6074_/X sky130_fd_sc_hd__clkbuf_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5025_/A VGND VGND VPWR VPWR _9740_/D sky130_fd_sc_hd__clkbuf_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9833_ _9833_/CLK _9833_/D _9730_/SET_B VGND VGND VPWR VPWR _9833_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6976_ _6976_/A _6976_/B _6976_/C VGND VGND VPWR VPWR _6977_/C sky130_fd_sc_hd__and3_2
XFILLER_65_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9764_ _9817_/CLK _9764_/D _9821_/SET_B VGND VGND VPWR VPWR _9764_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8715_ _8715_/A _8748_/A _8715_/C _8749_/B VGND VGND VPWR VPWR _8715_/X sky130_fd_sc_hd__or4_1
XFILLER_110_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5927_ _5990_/A _5927_/B VGND VGND VPWR VPWR _5928_/A sky130_fd_sc_hd__or2_1
XFILLER_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9695_ _9695_/CLK _9695_/D _9689_/SET_B VGND VGND VPWR VPWR _9695_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8646_ _8646_/A VGND VGND VPWR VPWR _8646_/X sky130_fd_sc_hd__clkbuf_1
X_5858_ _5990_/A _5858_/B VGND VGND VPWR VPWR _5859_/A sky130_fd_sc_hd__or2_1
X_5789_ _9280_/Q _5788_/A hold516/X _5788_/Y VGND VGND VPWR VPWR _5789_/X sky130_fd_sc_hd__a22o_1
X_8577_ _8577_/A _8710_/C _8657_/D _8741_/A VGND VGND VPWR VPWR _8583_/A sky130_fd_sc_hd__or4_2
X_4809_ _4805_/Y _5971_/B _4807_/Y _5513_/B VGND VGND VPWR VPWR _4809_/X sky130_fd_sc_hd__o22a_1
XFILLER_135_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7528_ _7528_/A VGND VGND VPWR VPWR _7528_/X sky130_fd_sc_hd__buf_4
XFILLER_174_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7459_ _7479_/A _9293_/Q _7479_/C _7471_/C VGND VGND VPWR VPWR _7508_/A sky130_fd_sc_hd__or4_4
XFILLER_162_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9129_ _8879_/A1 _9129_/D _6032_/X VGND VGND VPWR VPWR _9129_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6830_ _9168_/Q VGND VGND VPWR VPWR _6830_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6761_ _9554_/Q VGND VGND VPWR VPWR _6761_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_176_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5712_ _9302_/Q _5708_/A hold53/X _5708_/Y VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__a22o_1
X_8500_ _7903_/X _8361_/A _8138_/B _8592_/A VGND VGND VPWR VPWR _8656_/C sky130_fd_sc_hd__o22ai_2
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6692_ _9364_/Q VGND VGND VPWR VPWR _6692_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9480_ _9483_/CLK _9480_/D _9727_/SET_B VGND VGND VPWR VPWR _9480_/Q sky130_fd_sc_hd__dfrtp_1
X_5643_ _9339_/Q _5638_/A hold612/X _5638_/Y VGND VGND VPWR VPWR _5643_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8431_ _8431_/A VGND VGND VPWR VPWR _8560_/B sky130_fd_sc_hd__inv_2
XFILLER_163_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5574_ _9386_/Q _5572_/A hold510/X _5572_/Y VGND VGND VPWR VPWR _5574_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8362_ _8362_/A VGND VGND VPWR VPWR _8503_/A sky130_fd_sc_hd__inv_2
Xhold201 hold201/A VGND VGND VPWR VPWR hold202/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_129_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7313_ _6158_/Y _7171_/X _6122_/Y _7172_/X _7312_/X VGND VGND VPWR VPWR _7318_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4525_ _5282_/A _4525_/B VGND VGND VPWR VPWR _4526_/A sky130_fd_sc_hd__or2_1
Xhold212 hold212/A VGND VGND VPWR VPWR hold213/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 hold234/A VGND VGND VPWR VPWR hold235/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 hold223/A VGND VGND VPWR VPWR _9468_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_8293_ _8293_/A _8639_/B VGND VGND VPWR VPWR _8295_/A sky130_fd_sc_hd__or2_1
Xhold267 _5411_/X VGND VGND VPWR VPWR hold268/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 hold245/A VGND VGND VPWR VPWR hold245/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold278 hold278/A VGND VGND VPWR VPWR _9437_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold256 hold256/A VGND VGND VPWR VPWR hold257/A sky130_fd_sc_hd__dlygate4sd3_1
X_7244_ _6391_/Y _7167_/X _6499_/Y _7168_/X VGND VGND VPWR VPWR _7244_/X sky130_fd_sc_hd__o22a_1
XFILLER_49_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold289 hold289/A VGND VGND VPWR VPWR hold290/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7175_ _6819_/Y _7173_/X _6946_/Y _7174_/X VGND VGND VPWR VPWR _7175_/X sky130_fd_sc_hd__o22a_1
XFILLER_104_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6126_ _6121_/Y _5482_/B _6122_/Y _5521_/B _6125_/X VGND VGND VPWR VPWR _6127_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6057_ _9120_/Q _4485_/A _8965_/A1 _4485_/Y VGND VGND VPWR VPWR _9120_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5008_ _9743_/Q _4989_/A _4971_/A _4989_/Y VGND VGND VPWR VPWR _9743_/D sky130_fd_sc_hd__a22o_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_107 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _7046_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9816_ _9819_/CLK _9816_/D _9817_/SET_B VGND VGND VPWR VPWR _9816_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9747_ _4467_/A1 _9747_/D _4995_/X VGND VGND VPWR VPWR _9747_/Q sky130_fd_sc_hd__dfrtp_1
X_6959_ _9307_/Q VGND VGND VPWR VPWR _6959_/Y sky130_fd_sc_hd__inv_2
X_9678_ _9678_/CLK _9678_/D _9730_/SET_B VGND VGND VPWR VPWR _9678_/Q sky130_fd_sc_hd__dfrtp_1
X_8629_ _8629_/A _8648_/B VGND VGND VPWR VPWR _8723_/A sky130_fd_sc_hd__or2_1
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput306 _9770_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_2
Xoutput317 _9793_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_2
X_5290_ _5378_/A _5290_/B VGND VGND VPWR VPWR _5290_/X sky130_fd_sc_hd__or2_1
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput328 _9779_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_2
Xoutput339 _8861_/X VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_2
XFILLER_153_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8980_ _9128_/Q hold403/X _9093_/Q VGND VGND VPWR VPWR _8980_/X sky130_fd_sc_hd__mux2_1
X_7931_ _7957_/A _8347_/A _8489_/A _8347_/B VGND VGND VPWR VPWR _7931_/X sky130_fd_sc_hd__a211o_1
X_7862_ _7862_/A VGND VGND VPWR VPWR _8557_/A sky130_fd_sc_hd__clkbuf_4
X_9601_ _9686_/CLK _9601_/D _9817_/SET_B VGND VGND VPWR VPWR _9601_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7793_ _8436_/D VGND VGND VPWR VPWR _7873_/A sky130_fd_sc_hd__inv_2
X_6813_ _6809_/Y _4915_/X _4971_/Y _6196_/A _6812_/X VGND VGND VPWR VPWR _6814_/D
+ sky130_fd_sc_hd__o221a_1
X_6744_ _9494_/Q VGND VGND VPWR VPWR _6744_/Y sky130_fd_sc_hd__inv_4
X_9532_ _9582_/CLK _9532_/D _7042_/B VGND VGND VPWR VPWR _9532_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6675_ _9234_/Q VGND VGND VPWR VPWR _6675_/Y sky130_fd_sc_hd__inv_2
X_9463_ _9550_/CLK _9463_/D _9571_/SET_B VGND VGND VPWR VPWR _9463_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5626_ _9350_/Q _5622_/A _8969_/A1 _5622_/Y VGND VGND VPWR VPWR _9350_/D sky130_fd_sc_hd__a22o_1
X_8414_ _8414_/A _8687_/C _8621_/C _8757_/C VGND VGND VPWR VPWR _8417_/A sky130_fd_sc_hd__or4_4
X_9394_ _9694_/CLK _9394_/D _9689_/SET_B VGND VGND VPWR VPWR _9394_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5557_ _9397_/Q _5553_/A _6067_/B1 _5553_/Y VGND VGND VPWR VPWR _5557_/X sky130_fd_sc_hd__a22o_1
X_8345_ _8345_/A VGND VGND VPWR VPWR _8493_/A sky130_fd_sc_hd__inv_2
X_8276_ _8280_/A _8306_/B VGND VGND VPWR VPWR _8684_/B sky130_fd_sc_hd__nor2_1
X_4508_ _4682_/C _4508_/B _4823_/C VGND VGND VPWR VPWR _4913_/B sky130_fd_sc_hd__or3_4
XFILLER_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5488_ _9444_/Q _5484_/A _6064_/B1 _5484_/Y VGND VGND VPWR VPWR _9444_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7227_ _8835_/A _5756_/X _7737_/A _7071_/A _7226_/X VGND VGND VPWR VPWR _7230_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7158_ _6850_/Y _7095_/B _6957_/Y _7157_/X VGND VGND VPWR VPWR _7158_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6109_ _9525_/Q VGND VGND VPWR VPWR _6109_/Y sky130_fd_sc_hd__inv_2
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _7091_/C _7099_/B VGND VGND VPWR VPWR _7145_/A sky130_fd_sc_hd__or2_2
XFILLER_100_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4790_ _9688_/Q VGND VGND VPWR VPWR _4790_/Y sky130_fd_sc_hd__inv_4
XFILLER_82_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_18 _6127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _6282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6460_ _9819_/Q VGND VGND VPWR VPWR _6460_/Y sky130_fd_sc_hd__inv_4
X_5411_ _9497_/Q _5408_/A hold577/A _5408_/Y VGND VGND VPWR VPWR _5411_/X sky130_fd_sc_hd__a22o_1
X_6391_ _9366_/Q VGND VGND VPWR VPWR _6391_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_146_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8130_ _8260_/B _7874_/A _8144_/B VGND VGND VPWR VPWR _8161_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5342_ _5342_/A VGND VGND VPWR VPWR _5342_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8061_ _8068_/A _8171_/B VGND VGND VPWR VPWR _8445_/A sky130_fd_sc_hd__or2_1
X_7012_ _6660_/Y _7007_/A _9057_/Q _7007_/Y VGND VGND VPWR VPWR _9057_/D sky130_fd_sc_hd__o22a_1
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5273_ _9588_/Q _5265_/A _8975_/A1 _5265_/Y VGND VGND VPWR VPWR _9588_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8963_ _9648_/Q hold53/X _8975_/S VGND VGND VPWR VPWR _8963_/X sky130_fd_sc_hd__mux2_1
X_7914_ _8567_/A _7933_/B _7942_/C _8234_/A VGND VGND VPWR VPWR _8272_/A sky130_fd_sc_hd__or4_4
X_8894_ _8893_/X _9207_/Q _9096_/Q VGND VGND VPWR VPWR _8894_/X sky130_fd_sc_hd__mux2_1
X_7845_ _8702_/C _7917_/A VGND VGND VPWR VPWR _7846_/A sky130_fd_sc_hd__or2_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7776_ _9108_/Q _7776_/B VGND VGND VPWR VPWR _7776_/X sky130_fd_sc_hd__and2_1
XFILLER_184_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9515_ _9516_/CLK _9515_/D _9571_/SET_B VGND VGND VPWR VPWR _9515_/Q sky130_fd_sc_hd__dfrtp_2
X_4988_ _4988_/A VGND VGND VPWR VPWR _4989_/A sky130_fd_sc_hd__buf_8
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6727_ _6725_/Y _4869_/X _6726_/Y _5466_/B VGND VGND VPWR VPWR _6727_/X sky130_fd_sc_hd__o22a_1
XFILLER_176_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9446_ _9686_/CLK _9446_/D _9817_/SET_B VGND VGND VPWR VPWR _9446_/Q sky130_fd_sc_hd__dfrtp_1
X_6658_ _6658_/A _6658_/B _6658_/C _6658_/D VGND VGND VPWR VPWR _6659_/D sky130_fd_sc_hd__and4_1
XFILLER_191_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5609_ _5847_/A _5609_/B VGND VGND VPWR VPWR _5610_/A sky130_fd_sc_hd__or2_1
X_9377_ _9561_/CLK _9377_/D _7042_/B VGND VGND VPWR VPWR _9377_/Q sky130_fd_sc_hd__dfstp_1
X_8328_ _8627_/B _8763_/A _8328_/C VGND VGND VPWR VPWR _8329_/B sky130_fd_sc_hd__or3_1
XFILLER_152_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6589_ _6589_/A VGND VGND VPWR VPWR _6589_/Y sky130_fd_sc_hd__inv_2
X_8259_ _8288_/A _8258_/B _8049_/A _8257_/X _8258_/X VGND VGND VPWR VPWR _8259_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR _6416_/A sky130_fd_sc_hd__clkbuf_1
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR _6238_/A sky130_fd_sc_hd__clkbuf_1
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR _6536_/A sky130_fd_sc_hd__buf_4
XFILLER_108_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5960_ _5960_/A _5960_/B input150/X input153/X VGND VGND VPWR VPWR _5965_/B sky130_fd_sc_hd__or4bb_1
X_4911_ _4933_/A _4922_/B VGND VGND VPWR VPWR _5321_/B sky130_fd_sc_hd__or2_4
X_5891_ _5889_/X _8892_/X _8960_/X _9207_/Q VGND VGND VPWR VPWR _9207_/D sky130_fd_sc_hd__o22a_1
X_7630_ _6158_/Y _7497_/X _7627_/X _7629_/X VGND VGND VPWR VPWR _7640_/C sky130_fd_sc_hd__o211a_1
XFILLER_33_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4842_ _4835_/Y _4558_/B _4836_/Y _6058_/B _4841_/X VGND VGND VPWR VPWR _4852_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7561_ _8807_/A _7515_/X _6548_/Y _7516_/X VGND VGND VPWR VPWR _7561_/X sky130_fd_sc_hd__o22a_1
X_4773_ _4808_/A _4951_/A VGND VGND VPWR VPWR _5570_/B sky130_fd_sc_hd__or2_4
X_9300_ _9392_/CLK _9300_/D _9689_/SET_B VGND VGND VPWR VPWR _9300_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_158_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7492_ _7492_/A VGND VGND VPWR VPWR _7492_/X sky130_fd_sc_hd__buf_4
XFILLER_20_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6512_ _6510_/Y _5946_/B _6511_/Y _5589_/B VGND VGND VPWR VPWR _6512_/X sky130_fd_sc_hd__o22a_2
XFILLER_146_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9231_ _9679_/CLK _9231_/D _9730_/SET_B VGND VGND VPWR VPWR _9231_/Q sky130_fd_sc_hd__dfrtp_1
X_6443_ _9600_/Q VGND VGND VPWR VPWR _6443_/Y sky130_fd_sc_hd__clkinv_2
X_6374_ _9374_/Q VGND VGND VPWR VPWR _6374_/Y sky130_fd_sc_hd__inv_2
X_9162_ _9833_/CLK _9162_/D _9730_/SET_B VGND VGND VPWR VPWR _9162_/Q sky130_fd_sc_hd__dfrtp_1
X_8113_ _8229_/A _8479_/B VGND VGND VPWR VPWR _8582_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5325_ _9555_/Q _5323_/A _6065_/B1 _5323_/Y VGND VGND VPWR VPWR _9555_/D sky130_fd_sc_hd__a22o_1
X_9093_ _9751_/CLK _9093_/D _6076_/X VGND VGND VPWR VPWR _9093_/Q sky130_fd_sc_hd__dfrtp_4
X_8044_ _8436_/D _8179_/A VGND VGND VPWR VPWR _8045_/A sky130_fd_sc_hd__or2_1
XFILLER_142_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5256_ _5256_/A VGND VGND VPWR VPWR _5257_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5187_ _9646_/Q _5181_/A hold136/X _5181_/Y VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8946_ _7749_/X _9127_/Q _9093_/Q VGND VGND VPWR VPWR _8946_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8877_ _6613_/Y input92/X _8877_/S VGND VGND VPWR VPWR _8877_/X sky130_fd_sc_hd__mux2_2
XFILLER_12_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7828_ _8567_/A _7828_/B VGND VGND VPWR VPWR _7860_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7759_ _9741_/Q VGND VGND VPWR VPWR _7759_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9429_ _9800_/CLK _9429_/D _9797_/SET_B VGND VGND VPWR VPWR _9429_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_98_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold608 _5350_/X VGND VGND VPWR VPWR _9536_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold619 _9124_/Q VGND VGND VPWR VPWR hold619/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_170_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6090_ _9142_/Q VGND VGND VPWR VPWR _6090_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_69_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5110_ _9696_/Q _5105_/A _8975_/A1 _5105_/Y VGND VGND VPWR VPWR _9696_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5041_ _9735_/Q _5038_/A hold696/A _5038_/Y VGND VGND VPWR VPWR _5041_/X sky130_fd_sc_hd__a22o_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater403 _9797_/SET_B VGND VGND VPWR VPWR _9730_/SET_B sky130_fd_sc_hd__buf_12
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8800_ _8800_/A VGND VGND VPWR VPWR _8800_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_9780_ _9819_/CLK _9780_/D _9817_/SET_B VGND VGND VPWR VPWR _9780_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6992_ _9104_/Q VGND VGND VPWR VPWR _6993_/B sky130_fd_sc_hd__inv_2
X_8731_ _8731_/A _8751_/D _8755_/C _8756_/D VGND VGND VPWR VPWR _8731_/X sky130_fd_sc_hd__or4_1
XFILLER_25_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5943_ _9169_/Q _5937_/A _8965_/A1 _5937_/Y VGND VGND VPWR VPWR _9169_/D sky130_fd_sc_hd__a22o_1
X_5874_ _9221_/Q _5868_/A _8965_/A1 _5868_/Y VGND VGND VPWR VPWR _9221_/D sky130_fd_sc_hd__a22o_1
X_8662_ _8748_/A _8747_/B _8745_/B _8662_/D VGND VGND VPWR VPWR _8662_/Y sky130_fd_sc_hd__nor4_1
XFILLER_61_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7613_ _6256_/Y _7509_/X _6195_/Y _7510_/X VGND VGND VPWR VPWR _7613_/X sky130_fd_sc_hd__o22a_1
X_8593_ _8593_/A _8596_/B VGND VGND VPWR VPWR _8728_/C sky130_fd_sc_hd__nor2_1
XFILLER_21_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4825_ _4925_/B _4953_/B VGND VGND VPWR VPWR _5313_/B sky130_fd_sc_hd__or2_2
XFILLER_193_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7544_ _6675_/Y _7513_/X _6744_/Y _7514_/X _7543_/X VGND VGND VPWR VPWR _7549_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4756_ _4900_/A _4801_/B VGND VGND VPWR VPWR _5826_/B sky130_fd_sc_hd__or2_4
XFILLER_175_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4687_ _4920_/A _4865_/B VGND VGND VPWR VPWR _5935_/B sky130_fd_sc_hd__or2_4
X_7475_ _4737_/Y _7519_/A _4932_/Y _7520_/A _7474_/X VGND VGND VPWR VPWR _7482_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_108_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6426_ _6421_/Y _5378_/B _6422_/Y _5397_/B _6425_/X VGND VGND VPWR VPWR _6439_/B
+ sky130_fd_sc_hd__o221a_2
X_9214_ _9322_/CLK _9214_/D _9797_/SET_B VGND VGND VPWR VPWR _9214_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6357_ _6357_/A _6357_/B _6357_/C _6357_/D VGND VGND VPWR VPWR _6357_/Y sky130_fd_sc_hd__nand4_4
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9145_ _9679_/CLK _9145_/D _9730_/SET_B VGND VGND VPWR VPWR _9145_/Q sky130_fd_sc_hd__dfstp_1
X_5308_ _9565_/Q _5303_/A hold42/X _5303_/Y VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__a22o_1
XFILLER_161_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9076_ _9705_/CLK _9076_/D VGND VGND VPWR VPWR _9076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6288_ _6288_/A VGND VGND VPWR VPWR _6288_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_124_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8027_ _8593_/A VGND VGND VPWR VPWR _8027_/Y sky130_fd_sc_hd__inv_2
X_5239_ _9611_/Q _5237_/Y _6015_/B _5238_/Y VGND VGND VPWR VPWR _9611_/D sky130_fd_sc_hd__o22a_1
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8929_ _7341_/Y _9669_/Q _9001_/S VGND VGND VPWR VPWR _8929_/X sky130_fd_sc_hd__mux2_1
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold5 hold5/A VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_74_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xnet399_3 net399_3/A VGND VGND VPWR VPWR _6390_/A1 sky130_fd_sc_hd__inv_4
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4610_ _6189_/A _4818_/B VGND VGND VPWR VPWR _4611_/B sky130_fd_sc_hd__or2_4
X_5590_ _5590_/A VGND VGND VPWR VPWR _5591_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4541_ _6008_/B1 _9812_/Q _4541_/S VGND VGND VPWR VPWR _4541_/X sky130_fd_sc_hd__mux2_1
X_7260_ _6321_/Y _7149_/X _6339_/Y _7150_/X _7259_/X VGND VGND VPWR VPWR _7265_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4472_ _9617_/Q _4923_/A _9123_/Q VGND VGND VPWR VPWR _9032_/A sky130_fd_sc_hd__mux2_1
Xhold427 _4818_/B VGND VGND VPWR VPWR _4925_/B sky130_fd_sc_hd__clkbuf_2
Xhold416 _8989_/X VGND VGND VPWR VPWR hold417/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold405 _9126_/Q VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_6211_ _6209_/Y _5706_/B _6210_/Y _5687_/B VGND VGND VPWR VPWR _6218_/B sky130_fd_sc_hd__o22a_1
Xhold449 _5445_/X VGND VGND VPWR VPWR hold450/A sky130_fd_sc_hd__dlygate4sd3_1
X_7191_ _6698_/Y _7071_/C _6785_/Y _7146_/X VGND VGND VPWR VPWR _7191_/X sky130_fd_sc_hd__o22a_1
Xhold438 _6064_/X VGND VGND VPWR VPWR hold439/A sky130_fd_sc_hd__dlygate4sd3_1
X_6142_ _6142_/A _6142_/B _9811_/Q VGND VGND VPWR VPWR _6142_/X sky130_fd_sc_hd__or3b_4
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6073_ _6081_/A VGND VGND VPWR VPWR _6074_/A sky130_fd_sc_hd__clkbuf_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _8953_/X _9740_/Q _5024_/S VGND VGND VPWR VPWR _5025_/A sky130_fd_sc_hd__mux2_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9832_ _9832_/CLK _9832_/D _9821_/SET_B VGND VGND VPWR VPWR _9832_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6975_ _6975_/A _6975_/B _6975_/C VGND VGND VPWR VPWR _6976_/C sky130_fd_sc_hd__and3_1
X_9763_ _9817_/CLK _9763_/D _9821_/SET_B VGND VGND VPWR VPWR _9763_/Q sky130_fd_sc_hd__dfrtp_1
X_9694_ _9694_/CLK _9694_/D _9689_/SET_B VGND VGND VPWR VPWR _9694_/Q sky130_fd_sc_hd__dfrtp_1
X_8714_ _8745_/B _8714_/B _8714_/C VGND VGND VPWR VPWR _8715_/C sky130_fd_sc_hd__or3_1
XFILLER_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5926_ _8960_/X _7028_/A _5925_/Y _5889_/A _9180_/Q VGND VGND VPWR VPWR _9180_/D
+ sky130_fd_sc_hd__a32o_1
X_8645_ _8645_/A _8645_/B _8645_/C _8645_/D VGND VGND VPWR VPWR _8646_/A sky130_fd_sc_hd__or4_1
XFILLER_110_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5857_ _9232_/Q _5849_/A _8975_/A1 _5849_/Y VGND VGND VPWR VPWR _9232_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5788_ _5788_/A VGND VGND VPWR VPWR _5788_/Y sky130_fd_sc_hd__inv_2
X_8576_ _8513_/Y _8565_/Y _8560_/X _8512_/B VGND VGND VPWR VPWR _8741_/A sky130_fd_sc_hd__a31o_1
X_4808_ _4808_/A _4808_/B VGND VGND VPWR VPWR _5513_/B sky130_fd_sc_hd__or2_4
XFILLER_119_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4739_ _9349_/Q VGND VGND VPWR VPWR _4739_/Y sky130_fd_sc_hd__clkinv_2
X_7527_ _7527_/A VGND VGND VPWR VPWR _7527_/X sky130_fd_sc_hd__buf_4
XFILLER_134_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7458_ _7471_/A _7479_/C _9297_/Q VGND VGND VPWR VPWR _7507_/A sky130_fd_sc_hd__or3_2
XFILLER_162_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6409_ _9327_/Q VGND VGND VPWR VPWR _7424_/A sky130_fd_sc_hd__clkinv_2
XFILLER_122_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7389_ _6564_/Y _7067_/A _6510_/Y _7146_/A VGND VGND VPWR VPWR _7389_/X sky130_fd_sc_hd__o22a_1
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9128_ _9751_/CLK _9128_/D _6035_/X VGND VGND VPWR VPWR _9128_/Q sky130_fd_sc_hd__dfrtp_2
X_9059_ _9718_/CLK _9059_/D VGND VGND VPWR VPWR _9059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6760_ _9507_/Q VGND VGND VPWR VPWR _6760_/Y sky130_fd_sc_hd__clkinv_2
X_5711_ _9303_/Q _5708_/A hold577/A _5708_/Y VGND VGND VPWR VPWR _5711_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6691_ _6687_/Y _4545_/B _6688_/Y _5436_/B _6690_/X VGND VGND VPWR VPWR _6722_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_188_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5642_ _9340_/Q _5638_/A hold53/X _5638_/Y VGND VGND VPWR VPWR _9340_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8430_ _8139_/B _8439_/B _8212_/X VGND VGND VPWR VPWR _8673_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5573_ _9387_/Q _5572_/A hold516/X _5572_/Y VGND VGND VPWR VPWR _5573_/X sky130_fd_sc_hd__a22o_1
X_8361_ _8361_/A _8540_/B VGND VGND VPWR VPWR _8535_/C sky130_fd_sc_hd__nor2_1
Xhold202 hold202/A VGND VGND VPWR VPWR _9605_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7312_ _6140_/Y _7173_/X _6099_/Y _7174_/X VGND VGND VPWR VPWR _7312_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4524_ _4925_/A _4943_/A VGND VGND VPWR VPWR _4525_/B sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_18_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9694_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold213 hold213/A VGND VGND VPWR VPWR _9562_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold235 hold235/A VGND VGND VPWR VPWR _9354_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold224 _6066_/X VGND VGND VPWR VPWR hold225/A sky130_fd_sc_hd__dlygate4sd3_1
X_8292_ _8292_/A VGND VGND VPWR VPWR _8639_/B sky130_fd_sc_hd__inv_2
Xhold268 hold268/A VGND VGND VPWR VPWR hold269/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 hold518/X VGND VGND VPWR VPWR hold517/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold257 hold257/A VGND VGND VPWR VPWR _9570_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7243_ _7243_/A _7243_/B _7243_/C _7243_/D VGND VGND VPWR VPWR _7253_/B sky130_fd_sc_hd__and4_1
Xhold279 _5184_/X VGND VGND VPWR VPWR hold280/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7174_ _7174_/A VGND VGND VPWR VPWR _7174_/X sky130_fd_sc_hd__buf_4
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6125_ _6123_/Y _4598_/B _6124_/Y _4929_/X VGND VGND VPWR VPWR _6125_/X sky130_fd_sc_hd__o22a_4
XFILLER_98_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6056_ _9121_/Q _4485_/A hold696/X _4485_/Y VGND VGND VPWR VPWR _9121_/D sky130_fd_sc_hd__a22o_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _5007_/A VGND VGND VPWR VPWR _5007_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9815_ _9817_/CLK _9815_/D _7042_/B VGND VGND VPWR VPWR _9815_/Q sky130_fd_sc_hd__dfrtp_1
X_9746_ _4467_/A1 _9746_/D _4998_/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfrtp_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6958_ _9283_/Q VGND VGND VPWR VPWR _6958_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5909_ _9196_/Q _5904_/A _8964_/A1 _5904_/Y VGND VGND VPWR VPWR _9196_/D sky130_fd_sc_hd__a22o_1
X_6889_ _6884_/Y _5406_/B _6885_/Y _5329_/B _6888_/X VGND VGND VPWR VPWR _6908_/A
+ sky130_fd_sc_hd__o221a_2
X_9677_ _9730_/CLK _9677_/D _9730_/SET_B VGND VGND VPWR VPWR _9677_/Q sky130_fd_sc_hd__dfrtp_1
X_8628_ _8628_/A _8688_/B _8720_/B _8763_/B VGND VGND VPWR VPWR _8630_/B sky130_fd_sc_hd__or4_1
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8559_ _8559_/A VGND VGND VPWR VPWR _8559_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput307 _9774_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_2
XFILLER_153_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput318 _9775_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_2
Xoutput329 _9780_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_2
XFILLER_113_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7930_ _7935_/A _8347_/B VGND VGND VPWR VPWR _8483_/A sky130_fd_sc_hd__or2_1
XFILLER_82_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7861_ _8580_/C _7938_/A _8125_/A VGND VGND VPWR VPWR _7862_/A sky130_fd_sc_hd__or3_1
XFILLER_82_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9600_ _9600_/CLK _9600_/D _9821_/SET_B VGND VGND VPWR VPWR _9600_/Q sky130_fd_sc_hd__dfrtp_1
X_6812_ _6810_/Y _5313_/B _6811_/Y _5351_/B VGND VGND VPWR VPWR _6812_/X sky130_fd_sc_hd__o22a_1
X_7792_ _8567_/A _7933_/B _7942_/C _8570_/A VGND VGND VPWR VPWR _8436_/D sky130_fd_sc_hd__or4_4
XFILLER_90_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6743_ _9502_/Q VGND VGND VPWR VPWR _6743_/Y sky130_fd_sc_hd__clkinv_2
X_9531_ _9812_/CLK _9531_/D _9727_/SET_B VGND VGND VPWR VPWR _9531_/Q sky130_fd_sc_hd__dfrtp_1
X_6674_ _9275_/Q VGND VGND VPWR VPWR _6674_/Y sky130_fd_sc_hd__clkinv_2
X_9462_ _9550_/CLK _9462_/D _9571_/SET_B VGND VGND VPWR VPWR _9462_/Q sky130_fd_sc_hd__dfrtp_1
X_5625_ _9351_/Q _5622_/A _8965_/A1 _5622_/Y VGND VGND VPWR VPWR _9351_/D sky130_fd_sc_hd__a22o_1
X_8413_ _8750_/D _8548_/B VGND VGND VPWR VPWR _8757_/C sky130_fd_sc_hd__or2_1
XFILLER_191_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9393_ _9694_/CLK _9393_/D _9689_/SET_B VGND VGND VPWR VPWR _9393_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5556_ _9398_/Q _5553_/A hold217/X _5553_/Y VGND VGND VPWR VPWR _9398_/D sky130_fd_sc_hd__a22o_1
X_8344_ _8540_/B VGND VGND VPWR VPWR _8344_/Y sky130_fd_sc_hd__inv_2
X_4507_ _4507_/A VGND VGND VPWR VPWR _9828_/D sky130_fd_sc_hd__clkbuf_1
X_8275_ _8275_/A VGND VGND VPWR VPWR _8400_/B sky130_fd_sc_hd__inv_2
X_5487_ _9445_/Q _5484_/A hold696/X _5484_/Y VGND VGND VPWR VPWR _9445_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7226_ _8803_/A _7380_/B VGND VGND VPWR VPWR _7226_/X sky130_fd_sc_hd__or2_1
XFILLER_116_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7157_ _7157_/A VGND VGND VPWR VPWR _7157_/X sky130_fd_sc_hd__buf_4
X_6108_ _6103_/Y _5417_/B _6104_/Y _5340_/B _6107_/X VGND VGND VPWR VPWR _6127_/A
+ sky130_fd_sc_hd__o221a_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7161_/A _7181_/A _7156_/A _7150_/A VGND VGND VPWR VPWR _7094_/C sky130_fd_sc_hd__and4_1
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6039_ _9127_/Q _6026_/A _8952_/X _6026_/Y VGND VGND VPWR VPWR _9127_/D sky130_fd_sc_hd__a22o_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9729_ _9729_/CLK _9729_/D _9727_/SET_B VGND VGND VPWR VPWR _9729_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 _6127_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5410_ _9498_/Q _5408_/A hold510/X _5408_/Y VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__a22o_1
X_6390_ _6390_/A1 _6196_/A _6387_/Y _5647_/B _6389_/X VGND VGND VPWR VPWR _6390_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5341_ _5341_/A VGND VGND VPWR VPWR _5342_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8060_ _8443_/A _8431_/A _8053_/A _8443_/A _8059_/X VGND VGND VPWR VPWR _8060_/X
+ sky130_fd_sc_hd__o221a_1
X_7011_ _6506_/Y _7007_/A _9058_/Q _7007_/Y VGND VGND VPWR VPWR _9058_/D sky130_fd_sc_hd__o22a_2
X_5272_ _9589_/Q _5265_/A _8969_/A1 _5265_/Y VGND VGND VPWR VPWR _9589_/D sky130_fd_sc_hd__a22o_1
X_8962_ _9665_/Q hold696/A _8973_/S VGND VGND VPWR VPWR _8962_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7913_ _8280_/A _8268_/C VGND VGND VPWR VPWR _8281_/B sky130_fd_sc_hd__or2_4
X_8893_ _7550_/Y _9676_/Q _9020_/S VGND VGND VPWR VPWR _8893_/X sky130_fd_sc_hd__mux2_1
X_7844_ _7942_/C _8570_/A _8567_/A _7904_/D VGND VGND VPWR VPWR _7917_/A sky130_fd_sc_hd__or4_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7775_ _9110_/Q _7775_/A2 _9109_/Q _7775_/B2 _7774_/X VGND VGND VPWR VPWR _7775_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9514_ _9514_/CLK _9514_/D _9571_/SET_B VGND VGND VPWR VPWR _9514_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4987_ _9090_/Q _4987_/B _9093_/Q VGND VGND VPWR VPWR _4988_/A sky130_fd_sc_hd__or3_1
X_6726_ _9455_/Q VGND VGND VPWR VPWR _6726_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9445_ _9686_/CLK _9445_/D _9817_/SET_B VGND VGND VPWR VPWR _9445_/Q sky130_fd_sc_hd__dfrtp_1
X_6657_ _6652_/Y _4545_/B _8829_/A _5301_/B _6656_/X VGND VGND VPWR VPWR _6658_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_164_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5608_ _9362_/Q _5600_/A _8975_/A1 _5600_/Y VGND VGND VPWR VPWR _9362_/D sky130_fd_sc_hd__a22o_1
X_6588_ _9451_/Q VGND VGND VPWR VPWR _6588_/Y sky130_fd_sc_hd__inv_2
X_9376_ _9561_/CLK _9376_/D _7042_/B VGND VGND VPWR VPWR _9376_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5539_ _9409_/Q _5534_/A hold42/X _5534_/Y VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__a22o_1
X_8327_ _8518_/B _8327_/B VGND VGND VPWR VPWR _8328_/C sky130_fd_sc_hd__or2_1
XFILLER_105_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8258_ _8277_/A _8258_/B VGND VGND VPWR VPWR _8258_/X sky130_fd_sc_hd__or2_2
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7209_ _7209_/A _7209_/B _7209_/C VGND VGND VPWR VPWR _7209_/Y sky130_fd_sc_hd__nand3_4
X_8189_ _8189_/A _8619_/A VGND VGND VPWR VPWR _8191_/A sky130_fd_sc_hd__or2_1
XFILLER_19_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR _6293_/A sky130_fd_sc_hd__clkbuf_1
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR _6137_/A sky130_fd_sc_hd__clkbuf_1
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _6486_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_182_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5890_ _5889_/X _8894_/X _8960_/X _9208_/Q VGND VGND VPWR VPWR _9208_/D sky130_fd_sc_hd__o22a_1
X_4910_ _9552_/Q VGND VGND VPWR VPWR _4910_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4841_ _4838_/Y _5417_/B _4840_/Y _4644_/B VGND VGND VPWR VPWR _4841_/X sky130_fd_sc_hd__o22a_1
X_4772_ _9380_/Q VGND VGND VPWR VPWR _4772_/Y sky130_fd_sc_hd__clkinv_4
X_7560_ _8797_/A _7507_/X _8833_/A _7508_/X _7559_/X VGND VGND VPWR VPWR _7567_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_158_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7491_ _7491_/A VGND VGND VPWR VPWR _7491_/X sky130_fd_sc_hd__buf_4
X_6511_ _9373_/Q VGND VGND VPWR VPWR _6511_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9230_ _9679_/CLK _9230_/D _9730_/SET_B VGND VGND VPWR VPWR _9230_/Q sky130_fd_sc_hd__dfrtp_1
X_6442_ _6442_/A VGND VGND VPWR VPWR _6442_/Y sky130_fd_sc_hd__clkinv_2
X_9161_ _4471_/A1 _9161_/D _6177_/A VGND VGND VPWR VPWR _9161_/Q sky130_fd_sc_hd__dfrtp_4
X_8112_ _8243_/A _8118_/A VGND VGND VPWR VPWR _8755_/A sky130_fd_sc_hd__nor2_4
X_6373_ _9767_/Q VGND VGND VPWR VPWR _6373_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _9319_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_161_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5324_ _9556_/Q _5323_/A _6064_/B1 _5323_/Y VGND VGND VPWR VPWR _9556_/D sky130_fd_sc_hd__a22o_1
X_9092_ _9751_/CLK _9092_/D _6078_/X VGND VGND VPWR VPWR _9092_/Q sky130_fd_sc_hd__dfrtp_2
X_8043_ _8049_/A VGND VGND VPWR VPWR _8043_/Y sky130_fd_sc_hd__inv_2
X_5255_ _5282_/A _5255_/B VGND VGND VPWR VPWR _5256_/A sky130_fd_sc_hd__or2_1
XFILLER_114_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5186_ _9647_/Q _5181_/A hold42/X _5181_/Y VGND VGND VPWR VPWR _5186_/X sky130_fd_sc_hd__a22o_1
XFILLER_56_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8945_ _9653_/Q _8969_/A1 _8971_/S VGND VGND VPWR VPWR _8945_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8876_ _6516_/Y input90/X _8877_/S VGND VGND VPWR VPWR _8876_/X sky130_fd_sc_hd__mux2_2
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7827_ _7904_/D _7827_/B VGND VGND VPWR VPWR _7828_/B sky130_fd_sc_hd__nor2_1
XFILLER_156_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7758_ _9740_/Q VGND VGND VPWR VPWR _7758_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_184_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6709_ _6704_/Y _4865_/X _6705_/Y _4715_/X _6708_/X VGND VGND VPWR VPWR _6721_/B
+ sky130_fd_sc_hd__o221a_1
X_7689_ _6677_/Y _7521_/X _6761_/Y _7522_/X VGND VGND VPWR VPWR _7689_/X sky130_fd_sc_hd__o22a_1
XFILLER_137_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9428_ _9800_/CLK _9428_/D _9817_/SET_B VGND VGND VPWR VPWR _9428_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9359_ _9391_/CLK _9359_/D _9563_/SET_B VGND VGND VPWR VPWR _9359_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold609 _5465_/X VGND VGND VPWR VPWR _9458_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _9736_/Q _5038_/A hold510/X _5038_/Y VGND VGND VPWR VPWR _9736_/D sky130_fd_sc_hd__a22o_1
XFILLER_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater404 _9817_/SET_B VGND VGND VPWR VPWR _9797_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6991_ _4958_/Y _6983_/A _9070_/Q _6983_/Y VGND VGND VPWR VPWR _9070_/D sky130_fd_sc_hd__o22a_1
XFILLER_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8730_ _8730_/A _8730_/B _8730_/C VGND VGND VPWR VPWR _8756_/D sky130_fd_sc_hd__or3_1
X_5942_ _9170_/Q _5937_/A _8964_/A1 _5937_/Y VGND VGND VPWR VPWR _9170_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5873_ _9222_/Q _5868_/A _8964_/A1 _5868_/Y VGND VGND VPWR VPWR _9222_/D sky130_fd_sc_hd__a22o_1
X_8661_ _8661_/A _8749_/A _8748_/B _8661_/D VGND VGND VPWR VPWR _8662_/D sky130_fd_sc_hd__or4_1
X_7612_ _6249_/Y _7497_/X _7609_/X _7611_/X VGND VGND VPWR VPWR _7622_/C sky130_fd_sc_hd__o211a_1
X_8592_ _8592_/A _8596_/B VGND VGND VPWR VPWR _8669_/D sky130_fd_sc_hd__nor2_1
X_4824_ _4951_/B VGND VGND VPWR VPWR _4953_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4755_ _9246_/Q VGND VGND VPWR VPWR _4755_/Y sky130_fd_sc_hd__clkinv_4
X_7543_ _6768_/Y _7515_/X _6804_/Y _7516_/X VGND VGND VPWR VPWR _7543_/X sky130_fd_sc_hd__o22a_1
XFILLER_162_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4686_ _4806_/B VGND VGND VPWR VPWR _4865_/B sky130_fd_sc_hd__buf_2
X_7474_ _4755_/Y _7521_/A _4877_/Y _7522_/A VGND VGND VPWR VPWR _7474_/X sky130_fd_sc_hd__o22a_1
X_9213_ _9319_/CLK _9213_/D _9797_/SET_B VGND VGND VPWR VPWR _9213_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6425_ _6423_/Y _6112_/B _6424_/Y _5628_/B VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__o22a_1
XFILLER_161_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6356_ _6356_/A _6356_/B _6356_/C VGND VGND VPWR VPWR _6357_/D sky130_fd_sc_hd__and3_2
X_9144_ _9679_/CLK _9144_/D _9730_/SET_B VGND VGND VPWR VPWR _9144_/Q sky130_fd_sc_hd__dfrtp_1
X_9075_ _9705_/CLK _9075_/D VGND VGND VPWR VPWR _9075_/Q sky130_fd_sc_hd__dfxtp_1
X_5307_ _9566_/Q _5303_/A hold53/X _5303_/Y VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__a22o_1
XFILLER_115_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6287_ _9515_/Q VGND VGND VPWR VPWR _6287_/Y sky130_fd_sc_hd__inv_6
X_8026_ _8026_/A VGND VGND VPWR VPWR _8593_/A sky130_fd_sc_hd__buf_2
XFILLER_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5238_ _9090_/Q _7039_/A VGND VGND VPWR VPWR _5238_/Y sky130_fd_sc_hd__nor2_1
X_5169_ _5169_/A VGND VGND VPWR VPWR _5170_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_124_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8928_ _8927_/X _9186_/Q _9096_/Q VGND VGND VPWR VPWR _8928_/X sky130_fd_sc_hd__mux2_1
X_8859_ _8859_/A VGND VGND VPWR VPWR _8859_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_169_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold6 hold6/A VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4540_ _4953_/A _6189_/A _5250_/A VGND VGND VPWR VPWR _4541_/S sky130_fd_sc_hd__or3_2
X_4471_ _9618_/Q _4471_/A1 _9830_/Q VGND VGND VPWR VPWR _9033_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold406 _5517_/X VGND VGND VPWR VPWR hold407/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 hold417/A VGND VGND VPWR VPWR hold418/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6210_ _9317_/Q VGND VGND VPWR VPWR _6210_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7190_ _6748_/Y _7135_/X _6735_/Y _7136_/X _7189_/X VGND VGND VPWR VPWR _7209_/A
+ sky130_fd_sc_hd__o221a_1
Xhold428 _5519_/X VGND VGND VPWR VPWR _9423_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold439 hold439/A VGND VGND VPWR VPWR hold440/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6141_ _9551_/Q VGND VGND VPWR VPWR _6141_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6072_/A VGND VGND VPWR VPWR _6072_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5023_ _5023_/A VGND VGND VPWR VPWR _5023_/X sky130_fd_sc_hd__clkbuf_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9831_ _9831_/CLK _9831_/D _9727_/SET_B VGND VGND VPWR VPWR _9831_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6974_ _6969_/Y _5620_/B _6970_/Y _5786_/B _6973_/X VGND VGND VPWR VPWR _6975_/C
+ sky130_fd_sc_hd__o221a_1
X_9762_ _9810_/CLK _9762_/D _7042_/B VGND VGND VPWR VPWR _9762_/Q sky130_fd_sc_hd__dfstp_1
X_9693_ _9695_/CLK _9693_/D _9689_/SET_B VGND VGND VPWR VPWR _9693_/Q sky130_fd_sc_hd__dfrtp_1
X_8713_ _8777_/D _8741_/D _8713_/C _8745_/A VGND VGND VPWR VPWR _8713_/Y sky130_fd_sc_hd__nor4_1
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5925_ _9001_/X VGND VGND VPWR VPWR _5925_/Y sky130_fd_sc_hd__inv_2
X_5856_ _9233_/Q _5849_/A _8969_/A1 _5849_/Y VGND VGND VPWR VPWR _9233_/D sky130_fd_sc_hd__a22o_1
X_8644_ _8243_/A _8383_/A _8702_/C _7920_/A _8376_/X VGND VGND VPWR VPWR _8645_/D
+ sky130_fd_sc_hd__o221ai_2
XFILLER_179_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4807_ _9422_/Q VGND VGND VPWR VPWR _4807_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_166_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5787_ _5787_/A VGND VGND VPWR VPWR _5788_/A sky130_fd_sc_hd__clkbuf_4
X_8575_ _8558_/Y _8570_/Y _8560_/X _8506_/D VGND VGND VPWR VPWR _8657_/D sky130_fd_sc_hd__a31o_1
X_4738_ _4898_/B _4806_/B VGND VGND VPWR VPWR _5866_/B sky130_fd_sc_hd__or2_4
X_7526_ _7526_/A VGND VGND VPWR VPWR _7526_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_134_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4669_ _4669_/A VGND VGND VPWR VPWR _4669_/X sky130_fd_sc_hd__clkbuf_1
X_7457_ _4707_/Y _7497_/A _7450_/X _7456_/X VGND VGND VPWR VPWR _7483_/C sky130_fd_sc_hd__o211a_1
X_6408_ _9315_/Q VGND VGND VPWR VPWR _6408_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_79_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7388_ _6605_/Y _7135_/A _6646_/Y _7136_/A _7387_/X VGND VGND VPWR VPWR _7407_/A
+ sky130_fd_sc_hd__o221a_1
X_9127_ _8879_/A1 _9127_/D _6038_/X VGND VGND VPWR VPWR _9127_/Q sky130_fd_sc_hd__dfrtp_2
X_6339_ _9278_/Q VGND VGND VPWR VPWR _6339_/Y sky130_fd_sc_hd__inv_2
X_9058_ _9718_/CLK _9058_/D VGND VGND VPWR VPWR _9058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8009_ _8009_/A _8161_/B VGND VGND VPWR VPWR _8010_/A sky130_fd_sc_hd__or2_1
XFILLER_88_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5710_ _9304_/Q _5708_/A hold510/X _5708_/Y VGND VGND VPWR VPWR _5710_/X sky130_fd_sc_hd__a22o_1
X_6690_ _4808_/B _6189_/A _6689_/Y _4502_/B _6189_/X VGND VGND VPWR VPWR _6690_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_176_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5641_ _9341_/Q _5638_/A hold696/A _5638_/Y VGND VGND VPWR VPWR _5641_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5572_ _5572_/A VGND VGND VPWR VPWR _5572_/Y sky130_fd_sc_hd__clkinv_2
X_8360_ _8360_/A _8532_/C _8639_/C VGND VGND VPWR VPWR _8360_/X sky130_fd_sc_hd__or3_1
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7311_ _6096_/Y _7071_/D _6129_/Y _7166_/X _7310_/X VGND VGND VPWR VPWR _7318_/A
+ sky130_fd_sc_hd__o221a_1
X_4523_ _4750_/C _4642_/B _4689_/C _4750_/B VGND VGND VPWR VPWR _4808_/B sky130_fd_sc_hd__or4_4
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_2
X_8291_ _8552_/A _8296_/B VGND VGND VPWR VPWR _8292_/A sky130_fd_sc_hd__or2_1
Xhold214 _5416_/X VGND VGND VPWR VPWR hold215/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _5198_/X VGND VGND VPWR VPWR hold204/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 hold225/A VGND VGND VPWR VPWR hold226/A sky130_fd_sc_hd__dlygate4sd3_1
X_7242_ _6398_/Y _7160_/X _6470_/Y _7071_/B _7241_/X VGND VGND VPWR VPWR _7243_/D
+ sky130_fd_sc_hd__o221a_1
Xhold269 hold269/A VGND VGND VPWR VPWR _9497_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold258 _9747_/Q VGND VGND VPWR VPWR hold259/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold517/X VGND VGND VPWR VPWR hold516/A sky130_fd_sc_hd__buf_12
Xhold236 _5697_/X VGND VGND VPWR VPWR hold237/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7173_ _7173_/A VGND VGND VPWR VPWR _7173_/X sky130_fd_sc_hd__buf_4
XFILLER_131_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6124_/A VGND VGND VPWR VPWR _6124_/Y sky130_fd_sc_hd__clkinv_2
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _9751_/Q _6054_/Y _9122_/Q _6054_/A VGND VGND VPWR VPWR _9122_/D sky130_fd_sc_hd__a22o_1
X_5006_ _5017_/A VGND VGND VPWR VPWR _5007_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_100_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9814_ _9832_/CLK _9814_/D _9797_/SET_B VGND VGND VPWR VPWR _9814_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_109 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9745_ _4467_/A1 _9745_/D _5001_/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__dfrtp_1
X_6957_ _9312_/Q VGND VGND VPWR VPWR _6957_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5908_ _9197_/Q _5904_/A _8959_/A1 _5904_/Y VGND VGND VPWR VPWR _9197_/D sky130_fd_sc_hd__a22o_1
X_6888_ _6886_/Y _4937_/X _6887_/Y _5397_/B VGND VGND VPWR VPWR _6888_/X sky130_fd_sc_hd__o22a_1
X_9676_ _9833_/CLK _9676_/D _9730_/SET_B VGND VGND VPWR VPWR _9676_/Q sky130_fd_sc_hd__dfrtp_1
X_8627_ _8627_/A _8627_/B VGND VGND VPWR VPWR _8763_/B sky130_fd_sc_hd__or2_1
X_5839_ _5990_/A _5839_/B VGND VGND VPWR VPWR _5840_/A sky130_fd_sc_hd__or2_1
X_8558_ _8567_/C _8558_/B VGND VGND VPWR VPWR _8558_/Y sky130_fd_sc_hd__nor2_2
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7509_ _7509_/A VGND VGND VPWR VPWR _7509_/X sky130_fd_sc_hd__buf_4
X_8489_ _8489_/A _8489_/B VGND VGND VPWR VPWR _8489_/X sky130_fd_sc_hd__or2_1
XFILLER_190_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput308 _9784_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_2
XFILLER_141_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput319 _9794_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_2
X_7860_ _7860_/A _7860_/B _8580_/B VGND VGND VPWR VPWR _7938_/A sky130_fd_sc_hd__or3b_1
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6811_ _9533_/Q VGND VGND VPWR VPWR _6811_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7791_ _8702_/C VGND VGND VPWR VPWR _8324_/C sky130_fd_sc_hd__clkinv_2
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9530_ _9800_/CLK _9530_/D _9817_/SET_B VGND VGND VPWR VPWR _9530_/Q sky130_fd_sc_hd__dfrtp_1
X_6742_ _9580_/Q VGND VGND VPWR VPWR _6742_/Y sky130_fd_sc_hd__inv_2
X_9461_ _9550_/CLK _9461_/D _9563_/SET_B VGND VGND VPWR VPWR _9461_/Q sky130_fd_sc_hd__dfrtp_1
X_6673_ _6668_/Y _5826_/B _6669_/Y _5797_/B _6672_/X VGND VGND VPWR VPWR _6680_/B
+ sky130_fd_sc_hd__o221a_1
X_9392_ _9392_/CLK hold71/X _9689_/SET_B VGND VGND VPWR VPWR _9392_/Q sky130_fd_sc_hd__dfrtp_1
X_5624_ _9352_/Q _5622_/A _8964_/A1 _5622_/Y VGND VGND VPWR VPWR _9352_/D sky130_fd_sc_hd__a22o_1
X_8412_ _8412_/A _8641_/B VGND VGND VPWR VPWR _8621_/C sky130_fd_sc_hd__or2_1
XFILLER_164_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8343_ _8343_/A VGND VGND VPWR VPWR _8540_/B sky130_fd_sc_hd__buf_6
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5555_ _9399_/Q _5553_/A _6065_/B1 _5553_/Y VGND VGND VPWR VPWR _9399_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4506_ _8969_/A1 _9828_/Q _6049_/S VGND VGND VPWR VPWR _4507_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8274_ _8288_/A _8274_/B VGND VGND VPWR VPWR _8275_/A sky130_fd_sc_hd__or2_1
X_5486_ _9446_/Q _5484_/A hold510/X _5484_/Y VGND VGND VPWR VPWR _9446_/D sky130_fd_sc_hd__a22o_1
X_7225_ _7735_/A _7171_/X _8809_/A _7172_/X _7224_/X VGND VGND VPWR VPWR _7230_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7156_ _7156_/A VGND VGND VPWR VPWR _7156_/X sky130_fd_sc_hd__buf_4
X_6107_ _6105_/Y _4937_/X _6106_/Y _4883_/X VGND VGND VPWR VPWR _6107_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _9288_/Q _9287_/Q _7108_/C _7091_/C VGND VGND VPWR VPWR _7150_/A sky130_fd_sc_hd__or4_4
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6038_ _6038_/A VGND VGND VPWR VPWR _6038_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7989_ _8229_/B _8420_/B VGND VGND VPWR VPWR _8226_/A sky130_fd_sc_hd__or2_1
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9728_ _9728_/CLK _9728_/D _9727_/SET_B VGND VGND VPWR VPWR _9728_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9659_ _9830_/CLK _9659_/D _9537_/SET_B VGND VGND VPWR VPWR _9659_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9392_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_185_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5340_ _5378_/A _5340_/B VGND VGND VPWR VPWR _5341_/A sky130_fd_sc_hd__or2_1
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5271_ _9590_/Q _5265_/A _8965_/A1 _5265_/Y VGND VGND VPWR VPWR _9590_/D sky130_fd_sc_hd__a22o_1
X_7010_ _6357_/Y _7007_/A _9059_/Q _7007_/Y VGND VGND VPWR VPWR _9059_/D sky130_fd_sc_hd__o22a_1
XFILLER_114_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8961_ _9662_/Q _8965_/A1 _8973_/S VGND VGND VPWR VPWR _8961_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7912_ _7912_/A VGND VGND VPWR VPWR _8280_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8892_ _8891_/X _9206_/Q _9096_/Q VGND VGND VPWR VPWR _8892_/X sky130_fd_sc_hd__mux2_1
X_7843_ _8702_/C _8160_/A VGND VGND VPWR VPWR _8629_/A sky130_fd_sc_hd__nor2_2
XFILLER_102_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7774_ _9108_/Q _7774_/B VGND VGND VPWR VPWR _7774_/X sky130_fd_sc_hd__and2_1
X_4986_ _4986_/A VGND VGND VPWR VPWR _4986_/X sky130_fd_sc_hd__clkbuf_1
X_9513_ _9516_/CLK _9513_/D _9571_/SET_B VGND VGND VPWR VPWR _9513_/Q sky130_fd_sc_hd__dfrtp_2
X_6725_ _9572_/Q VGND VGND VPWR VPWR _6725_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6656_ _8823_/A _4511_/B _6655_/Y _4844_/X VGND VGND VPWR VPWR _6656_/X sky130_fd_sc_hd__o22a_1
X_9444_ _9561_/CLK _9444_/D _9817_/SET_B VGND VGND VPWR VPWR _9444_/Q sky130_fd_sc_hd__dfrtp_1
X_5607_ _9363_/Q _5600_/A hold593/X _5600_/Y VGND VGND VPWR VPWR _9363_/D sky130_fd_sc_hd__a22o_1
X_6587_ _9482_/Q VGND VGND VPWR VPWR _6587_/Y sky130_fd_sc_hd__clkinv_2
X_9375_ _9561_/CLK _9375_/D _9727_/SET_B VGND VGND VPWR VPWR _9375_/Q sky130_fd_sc_hd__dfrtp_1
X_5538_ _9410_/Q _5534_/A hold53/X _5534_/Y VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__a22o_1
X_8326_ _8581_/A _8326_/B VGND VGND VPWR VPWR _8327_/B sky130_fd_sc_hd__or2_1
XFILLER_117_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8257_ _8702_/A _8540_/A VGND VGND VPWR VPWR _8257_/X sky130_fd_sc_hd__or2_1
XFILLER_132_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7208_ _7208_/A _7208_/B _7208_/C _7208_/D VGND VGND VPWR VPWR _7209_/C sky130_fd_sc_hd__and4_1
X_5469_ _9457_/Q _5468_/A _6064_/B1 _5468_/Y VGND VGND VPWR VPWR _9457_/D sky130_fd_sc_hd__a22o_1
X_8188_ _8243_/B _8593_/A VGND VGND VPWR VPWR _8619_/A sky130_fd_sc_hd__nor2_1
X_7139_ _7139_/A VGND VGND VPWR VPWR _7139_/X sky130_fd_sc_hd__buf_4
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR _6239_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR _6649_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_155_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4840_ _9761_/Q VGND VGND VPWR VPWR _4840_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4771_ _4808_/A _4922_/B VGND VGND VPWR VPWR _5628_/B sky130_fd_sc_hd__or2_4
X_6510_ _9165_/Q VGND VGND VPWR VPWR _6510_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7490_ _6890_/Y _7485_/X _6922_/Y _7486_/X _7489_/X VGND VGND VPWR VPWR _7532_/A
+ sky130_fd_sc_hd__o221a_1
X_6441_ _9358_/Q VGND VGND VPWR VPWR _6441_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9160_ _9730_/CLK _9160_/D _9730_/SET_B VGND VGND VPWR VPWR _9160_/Q sky130_fd_sc_hd__dfrtp_1
X_6372_ _9587_/Q VGND VGND VPWR VPWR _6372_/Y sky130_fd_sc_hd__inv_2
X_8111_ _8557_/A _8229_/A _8110_/Y VGND VGND VPWR VPWR _8115_/A sky130_fd_sc_hd__o21bai_1
XFILLER_127_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5323_ _5323_/A VGND VGND VPWR VPWR _5323_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9091_ _9751_/CLK _9091_/D _6080_/X VGND VGND VPWR VPWR _9091_/Q sky130_fd_sc_hd__dfrtp_1
X_8042_ _8436_/D _8042_/B VGND VGND VPWR VPWR _8049_/A sky130_fd_sc_hd__or2_1
X_5254_ _5254_/A VGND VGND VPWR VPWR _5254_/X sky130_fd_sc_hd__clkbuf_1
X_5185_ _9648_/Q _5181_/A hold53/X _5181_/Y VGND VGND VPWR VPWR _5185_/X sky130_fd_sc_hd__a22o_1
XFILLER_83_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8944_ _9667_/Q hold516/X _8973_/S VGND VGND VPWR VPWR _8944_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8875_ _6522_/Y input82/X _8875_/S VGND VGND VPWR VPWR _8875_/X sky130_fd_sc_hd__mux2_2
XFILLER_83_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7826_ _8570_/B _7939_/A VGND VGND VPWR VPWR _8580_/C sky130_fd_sc_hd__nand2_2
XFILLER_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4969_ _4969_/A VGND VGND VPWR VPWR _4970_/A sky130_fd_sc_hd__clkbuf_1
X_7757_ _9130_/Q _7754_/B _7756_/Y _9131_/Q _7754_/Y VGND VGND VPWR VPWR _7757_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6708_ _6706_/Y _4634_/B _6707_/Y _4890_/X VGND VGND VPWR VPWR _6708_/X sky130_fd_sc_hd__o22a_1
X_7688_ _6713_/Y _7513_/X _6754_/Y _7514_/X _7687_/X VGND VGND VPWR VPWR _7693_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_164_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9427_ _9431_/CLK _9427_/D _9817_/SET_B VGND VGND VPWR VPWR _9427_/Q sky130_fd_sc_hd__dfrtp_1
X_6639_ _8817_/A _5367_/B _6635_/Y _5351_/B _6638_/X VGND VGND VPWR VPWR _6658_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9358_ _9391_/CLK hold92/X _9563_/SET_B VGND VGND VPWR VPWR _9358_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8309_ _8309_/A _8641_/B VGND VGND VPWR VPWR _8311_/A sky130_fd_sc_hd__or2_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9289_ _9297_/CLK _9289_/D _9797_/SET_B VGND VGND VPWR VPWR _9289_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater405 _9563_/SET_B VGND VGND VPWR VPWR _9689_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_93_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6990_ _6977_/Y _6983_/A _9071_/Q _6983_/Y VGND VGND VPWR VPWR _9071_/D sky130_fd_sc_hd__o22a_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5941_ _9171_/Q _5937_/A _8959_/A1 _5937_/Y VGND VGND VPWR VPWR _9171_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5872_ _9223_/Q _5868_/A _8959_/A1 _5868_/Y VGND VGND VPWR VPWR _5872_/X sky130_fd_sc_hd__a22o_1
X_8660_ _8557_/A _8229_/A _8563_/A _8557_/A VGND VGND VPWR VPWR _8748_/B sky130_fd_sc_hd__o22ai_2
XFILLER_178_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7611_ _6255_/Y _7500_/X _6230_/Y _7501_/X _7610_/X VGND VGND VPWR VPWR _7611_/X
+ sky130_fd_sc_hd__o221a_1
X_8591_ _8171_/B _8596_/B _8178_/B _8596_/B _8590_/X VGND VGND VPWR VPWR _8595_/A
+ sky130_fd_sc_hd__o221ai_1
X_4823_ _4823_/A _4823_/B _4823_/C VGND VGND VPWR VPWR _4937_/B sky130_fd_sc_hd__or3_4
XFILLER_193_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7542_ _6674_/Y _7507_/X _6735_/Y _7508_/X _7541_/X VGND VGND VPWR VPWR _7549_/A
+ sky130_fd_sc_hd__o221a_1
X_4754_ _4803_/A _4915_/B VGND VGND VPWR VPWR _5647_/B sky130_fd_sc_hd__or2_4
XFILLER_146_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7473_ _7473_/A _7479_/C _7478_/D VGND VGND VPWR VPWR _7522_/A sky130_fd_sc_hd__or3_2
XFILLER_174_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4685_ _4823_/A _4685_/B _4685_/C VGND VGND VPWR VPWR _4806_/B sky130_fd_sc_hd__or3_4
X_9212_ _9212_/CLK _9212_/D _9797_/SET_B VGND VGND VPWR VPWR _9212_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6424_ _9348_/Q VGND VGND VPWR VPWR _6424_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6355_ _6351_/Y _5598_/B _6352_/Y _5532_/B _6354_/Y VGND VGND VPWR VPWR _6356_/C
+ sky130_fd_sc_hd__o221a_1
X_9143_ _9679_/CLK _9143_/D _9730_/SET_B VGND VGND VPWR VPWR _9143_/Q sky130_fd_sc_hd__dfrtp_1
X_5306_ _9567_/Q _5303_/A hold577/A _5303_/Y VGND VGND VPWR VPWR _5306_/X sky130_fd_sc_hd__a22o_1
X_9074_ _9705_/CLK _9074_/D VGND VGND VPWR VPWR _9074_/Q sky130_fd_sc_hd__dfxtp_1
X_6286_ _6270_/Y _4937_/X _6273_/X _6279_/X _6285_/X VGND VGND VPWR VPWR _6357_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8025_ _8037_/B _8032_/B VGND VGND VPWR VPWR _8026_/A sky130_fd_sc_hd__or2_1
XFILLER_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5237_ _5237_/A _6015_/B VGND VGND VPWR VPWR _5237_/Y sky130_fd_sc_hd__nor2_1
X_5168_ _6165_/A _5179_/B VGND VGND VPWR VPWR _5169_/A sky130_fd_sc_hd__or2_1
XFILLER_96_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5099_ _9004_/X _9702_/Q _5101_/S VGND VGND VPWR VPWR _5100_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8927_ _7319_/Y _9681_/Q _9001_/S VGND VGND VPWR VPWR _8927_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8858_ _8858_/A VGND VGND VPWR VPWR _8858_/X sky130_fd_sc_hd__clkbuf_1
X_7809_ _7999_/A _8005_/A _7809_/C _7809_/D VGND VGND VPWR VPWR _7810_/D sky130_fd_sc_hd__nand4bb_1
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8789_ _8789_/A VGND VGND VPWR VPWR _8790_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold7 hold7/A VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4470_ _9619_/Q _4470_/A1 _9828_/Q VGND VGND VPWR VPWR _9034_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold407 hold407/A VGND VGND VPWR VPWR hold408/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 hold418/A VGND VGND VPWR VPWR _4689_/C sky130_fd_sc_hd__buf_2
XFILLER_7_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold429 _5520_/X VGND VGND VPWR VPWR _9422_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_171_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6140_ _9577_/Q VGND VGND VPWR VPWR _6140_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6071_/A VGND VGND VPWR VPWR _6072_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5022_ _6017_/A VGND VGND VPWR VPWR _5023_/A sky130_fd_sc_hd__clkbuf_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9830_ _9830_/CLK _9830_/D _9537_/SET_B VGND VGND VPWR VPWR _9830_/Q sky130_fd_sc_hd__dfrtp_2
X_6973_ _6971_/Y _5103_/B _6972_/Y _6165_/A VGND VGND VPWR VPWR _6973_/X sky130_fd_sc_hd__o22a_1
XFILLER_80_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9761_ _9810_/CLK _9761_/D _7042_/B VGND VGND VPWR VPWR _9761_/Q sky130_fd_sc_hd__dfrtp_1
X_9692_ _9695_/CLK hold74/X _9689_/SET_B VGND VGND VPWR VPWR _9692_/Q sky130_fd_sc_hd__dfrtp_1
X_8712_ _8745_/C _8747_/D _8712_/C _8749_/A VGND VGND VPWR VPWR _8713_/C sky130_fd_sc_hd__or4_1
X_5924_ _5889_/A _8916_/X _8960_/X _9181_/Q VGND VGND VPWR VPWR _9181_/D sky130_fd_sc_hd__o22a_1
X_5855_ _9234_/Q _5849_/A hold136/X _5849_/Y VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__a22o_1
X_8643_ _8643_/A _8738_/A _8704_/C _8643_/D VGND VGND VPWR VPWR _8645_/B sky130_fd_sc_hd__or4_1
XFILLER_179_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4806_ _4922_/B _4806_/B VGND VGND VPWR VPWR _5971_/B sky130_fd_sc_hd__or2_4
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5786_ _5847_/A _5786_/B VGND VGND VPWR VPWR _5787_/A sky130_fd_sc_hd__or2_1
XFILLER_119_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8574_ _8570_/Y _8567_/Y _8560_/X _8506_/B VGND VGND VPWR VPWR _8710_/C sky130_fd_sc_hd__a31o_1
X_4737_ _9219_/Q VGND VGND VPWR VPWR _4737_/Y sky130_fd_sc_hd__clkinv_4
X_7525_ _7525_/A VGND VGND VPWR VPWR _7525_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_147_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4668_ _4969_/A VGND VGND VPWR VPWR _4669_/A sky130_fd_sc_hd__clkbuf_1
X_7456_ _4684_/Y _7500_/A _4814_/Y _7501_/A _7455_/X VGND VGND VPWR VPWR _7456_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6407_ _6402_/Y _5706_/B _6403_/Y _5805_/B _6406_/X VGND VGND VPWR VPWR _6407_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4599_ _4599_/A VGND VGND VPWR VPWR _4600_/A sky130_fd_sc_hd__buf_2
X_9126_ _8879_/A1 _9126_/D _6041_/X VGND VGND VPWR VPWR _9126_/Q sky130_fd_sc_hd__dfrtp_2
X_7387_ _6528_/Y _7137_/A _6614_/Y _7138_/A _7386_/X VGND VGND VPWR VPWR _7387_/X
+ sky130_fd_sc_hd__o221a_1
X_6338_ _6338_/A _6338_/B _6338_/C _6338_/D VGND VGND VPWR VPWR _6357_/C sky130_fd_sc_hd__and4_2
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6269_ _6180_/A _6268_/Y _9084_/Q _6180_/Y VGND VGND VPWR VPWR _9084_/D sky130_fd_sc_hd__o22a_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9057_ _9718_/CLK _9057_/D VGND VGND VPWR VPWR _9057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8008_ _8008_/A _8260_/A VGND VGND VPWR VPWR _8161_/B sky130_fd_sc_hd__or2_1
XFILLER_29_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5640_ _9342_/Q _5638_/A hold510/X _5638_/Y VGND VGND VPWR VPWR _5640_/X sky130_fd_sc_hd__a22o_1
X_5571_ _5571_/A VGND VGND VPWR VPWR _5572_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_191_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7310_ _6172_/Y _7167_/X _6159_/Y _7168_/X VGND VGND VPWR VPWR _7310_/X sky130_fd_sc_hd__o22a_1
XFILLER_129_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8290_ _8290_/A _8532_/B _8359_/B VGND VGND VPWR VPWR _8293_/A sky130_fd_sc_hd__or3_1
X_4522_ _6083_/A VGND VGND VPWR VPWR _5282_/A sky130_fd_sc_hd__buf_6
Xhold215 hold215/A VGND VGND VPWR VPWR hold216/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 hold204/A VGND VGND VPWR VPWR _9638_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold226 hold226/A VGND VGND VPWR VPWR _9114_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7241_ _6403_/Y _7161_/X _6433_/Y _7162_/X VGND VGND VPWR VPWR _7241_/X sky130_fd_sc_hd__o22a_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold259 hold259/A VGND VGND VPWR VPWR hold260/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 _5304_/X VGND VGND VPWR VPWR hold249/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold237 hold237/A VGND VGND VPWR VPWR hold238/A sky130_fd_sc_hd__dlygate4sd3_1
X_7172_ _7172_/A VGND VGND VPWR VPWR _7172_/X sky130_fd_sc_hd__buf_4
XFILLER_98_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _9789_/Q VGND VGND VPWR VPWR _6123_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6054_/A VGND VGND VPWR VPWR _6054_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5005_ _9744_/Q _4989_/A _9743_/Q _4989_/Y VGND VGND VPWR VPWR _9744_/D sky130_fd_sc_hd__a22o_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9813_ _9831_/CLK _9813_/D _9727_/SET_B VGND VGND VPWR VPWR _9813_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_66_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9744_ _4467_/A1 _9744_/D _5004_/X VGND VGND VPWR VPWR _9744_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _6956_/A _6956_/B _6956_/C _6956_/D VGND VGND VPWR VPWR _6976_/B sky130_fd_sc_hd__and4_1
XFILLER_14_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5907_ _9198_/Q _5904_/A hold696/A _5904_/Y VGND VGND VPWR VPWR _5907_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6887_ _9501_/Q VGND VGND VPWR VPWR _6887_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9675_ _9833_/CLK _9675_/D _9730_/SET_B VGND VGND VPWR VPWR _9675_/Q sky130_fd_sc_hd__dfstp_1
X_8626_ _8382_/C _8586_/B _8625_/Y _8372_/B _8422_/B VGND VGND VPWR VPWR _8720_/B
+ sky130_fd_sc_hd__a311o_1
X_5838_ _9095_/Q _9833_/Q _5669_/Y _5837_/X VGND VGND VPWR VPWR _9245_/D sky130_fd_sc_hd__a31o_1
X_8557_ _8557_/A _8557_/B VGND VGND VPWR VPWR _8745_/B sky130_fd_sc_hd__nor2_1
X_5769_ _9287_/Q _5741_/A _5766_/B _5723_/A VGND VGND VPWR VPWR _9287_/D sky130_fd_sc_hd__o22a_1
XFILLER_135_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7508_ _7508_/A VGND VGND VPWR VPWR _7508_/X sky130_fd_sc_hd__buf_6
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8488_ _7903_/X _8383_/B _8049_/X _8487_/X _8053_/X VGND VGND VPWR VPWR _8490_/C
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_107_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7439_ _4919_/Y _7487_/A _4864_/Y _7488_/A VGND VGND VPWR VPWR _7439_/X sky130_fd_sc_hd__o22a_1
XFILLER_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9109_ _4471_/A1 _9109_/D _6177_/A VGND VGND VPWR VPWR _9109_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput309 _9785_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_2
XFILLER_153_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6810_ _9559_/Q VGND VGND VPWR VPWR _6810_/Y sky130_fd_sc_hd__clkinv_2
X_7790_ _7790_/A VGND VGND VPWR VPWR _8702_/C sky130_fd_sc_hd__buf_4
XFILLER_90_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6741_ _9468_/Q VGND VGND VPWR VPWR _6741_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9460_ _9550_/CLK _9460_/D _9571_/SET_B VGND VGND VPWR VPWR _9460_/Q sky130_fd_sc_hd__dfrtp_1
X_6672_ _6670_/Y _5805_/B _6671_/Y _5818_/B VGND VGND VPWR VPWR _6672_/X sky130_fd_sc_hd__o22a_1
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9391_ _9391_/CLK _9391_/D _9689_/SET_B VGND VGND VPWR VPWR _9391_/Q sky130_fd_sc_hd__dfrtp_4
X_5623_ _9353_/Q _5622_/A _8959_/A1 _5622_/Y VGND VGND VPWR VPWR _9353_/D sky130_fd_sc_hd__a22o_1
X_8411_ _8672_/B _8411_/B VGND VGND VPWR VPWR _8687_/C sky130_fd_sc_hd__or2_1
X_8342_ _8489_/A _8342_/B VGND VGND VPWR VPWR _8343_/A sky130_fd_sc_hd__or2_1
X_5554_ _9400_/Q _5553_/A _6064_/B1 _5553_/Y VGND VGND VPWR VPWR _9400_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8273_ _8273_/A _8718_/B _8700_/B _8615_/B VGND VGND VPWR VPWR _8279_/A sky130_fd_sc_hd__or4_1
X_4505_ _9829_/Q _4485_/A _8969_/A1 _4485_/Y VGND VGND VPWR VPWR _9829_/D sky130_fd_sc_hd__a22o_1
X_5485_ _9447_/Q _5484_/A hold516/X _5484_/Y VGND VGND VPWR VPWR _5485_/X sky130_fd_sc_hd__a22o_1
X_7224_ _8821_/A _7173_/X _8841_/A _7174_/X VGND VGND VPWR VPWR _7224_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7155_ _7155_/A VGND VGND VPWR VPWR _7155_/X sky130_fd_sc_hd__buf_4
XFILLER_100_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6106_ _6106_/A VGND VGND VPWR VPWR _6106_/Y sky130_fd_sc_hd__clkinv_4
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _7092_/A _7117_/B VGND VGND VPWR VPWR _7156_/A sky130_fd_sc_hd__or2_4
XFILLER_132_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6037_ _6071_/A VGND VGND VPWR VPWR _6038_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_46_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7988_ _8182_/B VGND VGND VPWR VPWR _8420_/B sky130_fd_sc_hd__buf_6
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6939_ _9689_/Q VGND VGND VPWR VPWR _6939_/Y sky130_fd_sc_hd__inv_2
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9727_ _9729_/CLK _9727_/D _9727_/SET_B VGND VGND VPWR VPWR _9727_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_14_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9658_ _9830_/CLK _9658_/D _9537_/SET_B VGND VGND VPWR VPWR _9658_/Q sky130_fd_sc_hd__dfrtp_1
X_8609_ _8682_/A _8608_/Y _8394_/A VGND VGND VPWR VPWR _8683_/B sky130_fd_sc_hd__o21ai_1
XFILLER_10_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9589_ _9832_/CLK _9589_/D _9821_/SET_B VGND VGND VPWR VPWR _9589_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_157_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_csclk _8889_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_135_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold590 _5852_/X VGND VGND VPWR VPWR _9237_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_0_1_csclk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5270_ _9591_/Q _5265_/A _8964_/A1 _5265_/Y VGND VGND VPWR VPWR _9591_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8960_ _9097_/Q _8861_/X _9096_/Q VGND VGND VPWR VPWR _8960_/X sky130_fd_sc_hd__mux2_8
X_7911_ _8005_/A _8230_/A _7999_/A _8570_/A VGND VGND VPWR VPWR _7912_/A sky130_fd_sc_hd__or4_4
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8891_ _7532_/Y _9675_/Q _9020_/S VGND VGND VPWR VPWR _8891_/X sky130_fd_sc_hd__mux2_1
X_7842_ _8436_/D _8068_/A VGND VGND VPWR VPWR _8160_/A sky130_fd_sc_hd__or2_2
XFILLER_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7773_ _9110_/Q _7773_/A2 _9109_/Q _7773_/B2 _7772_/X VGND VGND VPWR VPWR _7773_/X
+ sky130_fd_sc_hd__a221o_1
X_4985_ _5017_/A VGND VGND VPWR VPWR _4986_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_168_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6724_ _9382_/Q VGND VGND VPWR VPWR _6724_/Y sky130_fd_sc_hd__clkinv_2
X_9512_ _9514_/CLK _9512_/D _9571_/SET_B VGND VGND VPWR VPWR _9512_/Q sky130_fd_sc_hd__dfrtp_1
X_9443_ _9791_/CLK _9443_/D _9817_/SET_B VGND VGND VPWR VPWR _9443_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6655_ _6655_/A VGND VGND VPWR VPWR _6655_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5606_ _9364_/Q _5600_/A hold136/X _5600_/Y VGND VGND VPWR VPWR _5606_/X sky130_fd_sc_hd__a22o_1
X_9374_ _9431_/CLK _9374_/D _9797_/SET_B VGND VGND VPWR VPWR _9374_/Q sky130_fd_sc_hd__dfstp_1
X_6586_ _9404_/Q VGND VGND VPWR VPWR _6586_/Y sky130_fd_sc_hd__clkinv_2
X_5537_ _9411_/Q _5534_/A hold577/A _5534_/Y VGND VGND VPWR VPWR _5537_/X sky130_fd_sc_hd__a22o_1
X_8325_ _8325_/A _8372_/B VGND VGND VPWR VPWR _8326_/B sky130_fd_sc_hd__or2_1
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8256_ _8353_/B VGND VGND VPWR VPWR _8256_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7207_ _6798_/Y _7180_/X _6769_/Y _7181_/X _7206_/X VGND VGND VPWR VPWR _7208_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5468_ _5468_/A VGND VGND VPWR VPWR _5468_/Y sky130_fd_sc_hd__inv_2
X_8187_ _8027_/Y _8586_/B _8186_/X VGND VGND VPWR VPWR _8189_/A sky130_fd_sc_hd__a21o_1
X_5399_ _5399_/A VGND VGND VPWR VPWR _5399_/Y sky130_fd_sc_hd__inv_2
X_7138_ _7138_/A VGND VGND VPWR VPWR _7138_/X sky130_fd_sc_hd__buf_4
XFILLER_59_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7069_ _9288_/Q _9287_/Q _7129_/B _7091_/C VGND VGND VPWR VPWR _7070_/A sky130_fd_sc_hd__or4_4
XFILLER_59_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR _6124_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ _9344_/Q VGND VGND VPWR VPWR _4770_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6440_ _9457_/Q VGND VGND VPWR VPWR _6440_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6371_ _9582_/Q VGND VGND VPWR VPWR _6371_/Y sky130_fd_sc_hd__clkinv_2
X_8110_ _8110_/A _8244_/A VGND VGND VPWR VPWR _8110_/Y sky130_fd_sc_hd__nand2_1
X_5322_ _5322_/A VGND VGND VPWR VPWR _5323_/A sky130_fd_sc_hd__clkbuf_2
X_9090_ _9751_/CLK _9090_/D _6082_/X VGND VGND VPWR VPWR _9090_/Q sky130_fd_sc_hd__dfstp_4
X_8041_ _8053_/A _8158_/A VGND VGND VPWR VPWR _8654_/A sky130_fd_sc_hd__nor2_1
X_5253_ _6008_/B1 _9601_/Q _5253_/S VGND VGND VPWR VPWR _5254_/A sky130_fd_sc_hd__mux2_1
X_5184_ _9649_/Q _5181_/A hold577/A _5181_/Y VGND VGND VPWR VPWR _5184_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8943_ _9663_/Q _8964_/A1 _8973_/S VGND VGND VPWR VPWR _8943_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8874_ _6575_/Y _9100_/Q _9019_/S VGND VGND VPWR VPWR _8874_/X sky130_fd_sc_hd__mux2_1
X_7825_ _7942_/C _7860_/A _8570_/A _8234_/A _7823_/X VGND VGND VPWR VPWR _7939_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4968_ _9752_/Q _9738_/Q _9092_/Q _6024_/B VGND VGND VPWR VPWR _9752_/D sky130_fd_sc_hd__o211a_1
X_7756_ _9131_/Q VGND VGND VPWR VPWR _7756_/Y sky130_fd_sc_hd__inv_2
X_6707_ _6707_/A VGND VGND VPWR VPWR _6707_/Y sky130_fd_sc_hd__inv_2
X_4899_ _9414_/Q VGND VGND VPWR VPWR _4899_/Y sky130_fd_sc_hd__inv_2
X_7687_ _6693_/Y _7515_/X _6776_/Y _7516_/X VGND VGND VPWR VPWR _7687_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9426_ _9574_/CLK _9426_/D _9571_/SET_B VGND VGND VPWR VPWR _9426_/Q sky130_fd_sc_hd__dfrtp_1
X_6638_ _8811_/A _5482_/B _6637_/Y _5313_/B VGND VGND VPWR VPWR _6638_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9357_ _9391_/CLK hold98/X _9563_/SET_B VGND VGND VPWR VPWR _9357_/Q sky130_fd_sc_hd__dfrtp_1
X_6569_ _6569_/A VGND VGND VPWR VPWR _6569_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_152_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8308_ _8552_/A _8312_/B VGND VGND VPWR VPWR _8641_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_16_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9420_/CLK sky130_fd_sc_hd__clkbuf_16
X_9288_ _9297_/CLK _9288_/D _9797_/SET_B VGND VGND VPWR VPWR _9288_/Q sky130_fd_sc_hd__dfstp_2
X_8239_ _8567_/A _8625_/B _8625_/C VGND VGND VPWR VPWR _8255_/B sky130_fd_sc_hd__or3_1
XFILLER_160_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater406 _9537_/SET_B VGND VGND VPWR VPWR _9563_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5940_ _9172_/Q _5937_/A hold696/X _5937_/Y VGND VGND VPWR VPWR _9172_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5871_ _9224_/Q _5868_/A hold577/A _5868_/Y VGND VGND VPWR VPWR _5871_/X sky130_fd_sc_hd__a22o_1
X_7610_ _6202_/Y _7502_/X _6200_/Y _7503_/X VGND VGND VPWR VPWR _7610_/X sky130_fd_sc_hd__o22a_1
XFILLER_61_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8590_ _8435_/Y _8596_/B _8443_/A _8596_/B _8589_/X VGND VGND VPWR VPWR _8590_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4822_ _9557_/Q VGND VGND VPWR VPWR _4822_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_193_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4753_ _9328_/Q VGND VGND VPWR VPWR _4753_/Y sky130_fd_sc_hd__clkinv_4
X_7541_ _6741_/Y _7509_/X _6798_/Y _7510_/X VGND VGND VPWR VPWR _7541_/X sky130_fd_sc_hd__o22a_1
X_7472_ _7479_/A _9293_/Q _7478_/C _9297_/Q VGND VGND VPWR VPWR _7521_/A sky130_fd_sc_hd__or4_4
X_6423_ _9436_/Q VGND VGND VPWR VPWR _6423_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4684_ _9167_/Q VGND VGND VPWR VPWR _4684_/Y sky130_fd_sc_hd__clkinv_4
X_9211_ _9212_/CLK _9211_/D _9797_/SET_B VGND VGND VPWR VPWR _9211_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6354_ _8860_/A _4700_/Y input57/X _6353_/Y VGND VGND VPWR VPWR _6354_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9142_ _9577_/CLK _9142_/D _9571_/SET_B VGND VGND VPWR VPWR _9142_/Q sky130_fd_sc_hd__dfrtp_1
X_5305_ _9568_/Q _5303_/A hold510/X _5303_/Y VGND VGND VPWR VPWR _5305_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9073_ _9718_/CLK _9073_/D VGND VGND VPWR VPWR _9073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6285_ _6280_/Y _4854_/X _6281_/Y _5133_/B _6284_/X VGND VGND VPWR VPWR _6285_/X
+ sky130_fd_sc_hd__o221a_2
X_8024_ _8567_/A _8132_/B _8139_/A VGND VGND VPWR VPWR _8037_/B sky130_fd_sc_hd__or3_2
XFILLER_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5236_ _5236_/A VGND VGND VPWR VPWR _5236_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5167_ _9660_/Q _5159_/A _8975_/A1 _5159_/Y VGND VGND VPWR VPWR _9660_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5098_ _5098_/A VGND VGND VPWR VPWR _9703_/D sky130_fd_sc_hd__clkbuf_1
X_8926_ _8925_/X _9185_/Q _9096_/Q VGND VGND VPWR VPWR _8926_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7808_ _8567_/A VGND VGND VPWR VPWR _8005_/A sky130_fd_sc_hd__inv_2
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8788_ _8788_/A VGND VGND VPWR VPWR _8788_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7739_ _9091_/Q _9094_/Q VGND VGND VPWR VPWR _7739_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9409_ _9695_/CLK hold86/X _9689_/SET_B VGND VGND VPWR VPWR _9409_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold8 hold8/A VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_74_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold408 hold408/A VGND VGND VPWR VPWR _9425_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_171_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold419 _4808_/B VGND VGND VPWR VPWR _4943_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _6081_/A VGND VGND VPWR VPWR _6017_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9760_ net399_3/A _9760_/D _4969_/A VGND VGND VPWR VPWR _9760_/Q sky130_fd_sc_hd__dfrtn_1
X_8711_ _8755_/A _8745_/D _8748_/B VGND VGND VPWR VPWR _8712_/C sky130_fd_sc_hd__or3_1
X_6972_ _6972_/A VGND VGND VPWR VPWR _6972_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9691_ _9695_/CLK hold80/X _9689_/SET_B VGND VGND VPWR VPWR _9691_/Q sky130_fd_sc_hd__dfrtp_1
X_5923_ _5889_/A _8918_/X _8960_/X _9182_/Q VGND VGND VPWR VPWR _9182_/D sky130_fd_sc_hd__o22a_1
X_5854_ _9235_/Q _5849_/A hold612/X _5849_/Y VGND VGND VPWR VPWR _5854_/X sky130_fd_sc_hd__a22o_1
X_8642_ _8642_/A _8642_/B VGND VGND VPWR VPWR _8704_/C sky130_fd_sc_hd__or2_1
X_8573_ _8649_/A _8573_/B _8776_/D _8656_/D VGND VGND VPWR VPWR _8577_/A sky130_fd_sc_hd__or4_1
X_4805_ _9156_/Q VGND VGND VPWR VPWR _4805_/Y sky130_fd_sc_hd__inv_2
X_7524_ _6951_/Y _7519_/X _6863_/Y _7520_/X _7523_/X VGND VGND VPWR VPWR _7531_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5785_ _5741_/Y _5779_/Y _5784_/Y _9281_/Q _5784_/A VGND VGND VPWR VPWR _9281_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_147_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4736_ _4726_/Y _5698_/B _4728_/Y _5805_/B _4735_/X VGND VGND VPWR VPWR _4812_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4667_ _9757_/Q _4657_/A _8992_/X _4657_/Y VGND VGND VPWR VPWR _9757_/D sky130_fd_sc_hd__a22o_2
X_7455_ _4868_/Y _7502_/A _4948_/Y _7503_/A VGND VGND VPWR VPWR _7455_/X sky130_fd_sc_hd__o22a_1
XFILLER_79_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7386_ _6587_/Y _7139_/A _6643_/Y _7140_/A VGND VGND VPWR VPWR _7386_/X sky130_fd_sc_hd__o22a_1
X_6406_ _6404_/Y _5818_/B _6405_/Y _5797_/B VGND VGND VPWR VPWR _6406_/X sky130_fd_sc_hd__o22a_2
XFILLER_162_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6337_ _6332_/Y _5805_/B _6333_/Y _5902_/B _6336_/X VGND VGND VPWR VPWR _6338_/D
+ sky130_fd_sc_hd__o221a_1
X_4598_ _5201_/A _4598_/B VGND VGND VPWR VPWR _4599_/A sky130_fd_sc_hd__or2_1
X_9125_ _8879_/A1 _9125_/D _6044_/X VGND VGND VPWR VPWR _9125_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_135_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6268_ _6268_/A _6268_/B _6268_/C _6268_/D VGND VGND VPWR VPWR _6268_/Y sky130_fd_sc_hd__nand4_4
X_9056_ _9718_/CLK _9056_/D VGND VGND VPWR VPWR _9056_/Q sky130_fd_sc_hd__dfxtp_1
X_8007_ _7789_/B _8144_/B _7789_/B _8144_/B VGND VGND VPWR VPWR _8008_/A sky130_fd_sc_hd__o2bb2a_1
X_6199_ _9568_/Q VGND VGND VPWR VPWR _6199_/Y sky130_fd_sc_hd__inv_2
X_5219_ _9625_/Q _5216_/Y _8962_/X _5216_/A VGND VGND VPWR VPWR _9625_/D sky130_fd_sc_hd__o22a_1
XFILLER_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8909_ _7694_/Y _9671_/Q _9020_/S VGND VGND VPWR VPWR _8909_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5570_ _5570_/A _5570_/B VGND VGND VPWR VPWR _5571_/A sky130_fd_sc_hd__or2_1
XFILLER_129_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ _9820_/Q _4513_/A _8975_/A1 _4513_/Y VGND VGND VPWR VPWR _9820_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold216 hold216/A VGND VGND VPWR VPWR _9492_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold205 _5606_/X VGND VGND VPWR VPWR hold206/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7240_ _6387_/Y _7155_/X _6423_/Y _7156_/X _7239_/X VGND VGND VPWR VPWR _7243_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold249 hold249/A VGND VGND VPWR VPWR hold250/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _5503_/X VGND VGND VPWR VPWR hold228/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold238 hold238/A VGND VGND VPWR VPWR _9311_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7171_ _7171_/A VGND VGND VPWR VPWR _7171_/X sky130_fd_sc_hd__buf_4
X_6122_ _9421_/Q VGND VGND VPWR VPWR _6122_/Y sky130_fd_sc_hd__clkinv_2
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6053_/A _6053_/B _6053_/C _6053_/D VGND VGND VPWR VPWR _6054_/A sky130_fd_sc_hd__or4_1
X_5004_ _5004_/A VGND VGND VPWR VPWR _5004_/X sky130_fd_sc_hd__clkbuf_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9812_ _9812_/CLK _9812_/D _7042_/B VGND VGND VPWR VPWR _9812_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9743_ _4467_/A1 _9743_/D _5007_/X VGND VGND VPWR VPWR _9743_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _6950_/Y _5979_/B _6951_/Y _5866_/B _6954_/X VGND VGND VPWR VPWR _6956_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5906_ _9199_/Q _5904_/A hold510/X _5904_/Y VGND VGND VPWR VPWR _9199_/D sky130_fd_sc_hd__a22o_1
X_9674_ _9833_/CLK _9674_/D _9730_/SET_B VGND VGND VPWR VPWR _9674_/Q sky130_fd_sc_hd__dfstp_1
X_8625_ _8625_/A _8625_/B _8625_/C VGND VGND VPWR VPWR _8625_/Y sky130_fd_sc_hd__nor3_1
X_6886_ _9467_/Q VGND VGND VPWR VPWR _6886_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5837_ _9098_/Q _5718_/A _5669_/Y _5782_/B _9245_/Q VGND VGND VPWR VPWR _5837_/X
+ sky130_fd_sc_hd__o221a_1
X_8556_ _8556_/A _8556_/B _8556_/C VGND VGND VPWR VPWR _8647_/B sky130_fd_sc_hd__or3_1
X_5768_ _5768_/A VGND VGND VPWR VPWR _9288_/D sky130_fd_sc_hd__inv_2
X_8487_ _8314_/A _7953_/A _8205_/A _8567_/C _8126_/A VGND VGND VPWR VPWR _8487_/X
+ sky130_fd_sc_hd__a311o_1
X_4719_ _9175_/Q VGND VGND VPWR VPWR _4719_/Y sky130_fd_sc_hd__clkinv_2
X_7507_ _7507_/A VGND VGND VPWR VPWR _7507_/X sky130_fd_sc_hd__buf_6
XFILLER_190_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5699_ _5699_/A VGND VGND VPWR VPWR _5700_/A sky130_fd_sc_hd__clkbuf_2
X_7438_ _7467_/A _7477_/A _9297_/Q VGND VGND VPWR VPWR _7488_/A sky130_fd_sc_hd__or3_2
XFILLER_162_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7369_ _6811_/Y _7151_/X _6742_/Y _7152_/X VGND VGND VPWR VPWR _7369_/X sky130_fd_sc_hd__o22a_1
X_9108_ _4471_/A1 _9108_/D _6177_/A VGND VGND VPWR VPWR _9108_/Q sky130_fd_sc_hd__dfrtp_4
X_9039_ _9607_/Q _8813_/A VGND VGND VPWR VPWR _9039_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_130_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6740_ _6735_/Y _5378_/B _6736_/Y _5359_/B _6739_/X VGND VGND VPWR VPWR _6747_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6671_ _9256_/Q VGND VGND VPWR VPWR _6671_/Y sky130_fd_sc_hd__inv_2
X_9390_ _9391_/CLK _9390_/D _9689_/SET_B VGND VGND VPWR VPWR _9390_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5622_ _5622_/A VGND VGND VPWR VPWR _5622_/Y sky130_fd_sc_hd__inv_2
X_8410_ _8410_/A _8619_/C _8717_/A _8620_/C VGND VGND VPWR VPWR _8414_/A sky130_fd_sc_hd__or4_1
X_8341_ _8341_/A _8341_/B VGND VGND VPWR VPWR _8342_/B sky130_fd_sc_hd__nor2_1
X_5553_ _5553_/A VGND VGND VPWR VPWR _5553_/Y sky130_fd_sc_hd__inv_2
X_4504_ _4504_/A VGND VGND VPWR VPWR _9830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8272_ _8272_/A _8302_/B VGND VGND VPWR VPWR _8615_/B sky130_fd_sc_hd__nor2_1
X_5484_ _5484_/A VGND VGND VPWR VPWR _5484_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_172_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7223_ _8789_/A _7071_/D _8807_/A _7166_/X _7222_/X VGND VGND VPWR VPWR _7230_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7154_ _6896_/Y _7149_/X _6970_/Y _7150_/X _7153_/X VGND VGND VPWR VPWR _7165_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6105_ _9473_/Q VGND VGND VPWR VPWR _6105_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_86_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7085_ _7092_/A _7100_/B VGND VGND VPWR VPWR _7181_/A sky130_fd_sc_hd__or2_2
XFILLER_132_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _9128_/Q _6026_/A _8946_/X _6026_/Y VGND VGND VPWR VPWR _9128_/D sky130_fd_sc_hd__a22o_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7987_ _7987_/A VGND VGND VPWR VPWR _8182_/B sky130_fd_sc_hd__clkbuf_8
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _6933_/Y _5047_/B _6934_/Y _6166_/A _6937_/X VGND VGND VPWR VPWR _6956_/A
+ sky130_fd_sc_hd__o221a_1
X_9726_ _9728_/CLK _9726_/D _9727_/SET_B VGND VGND VPWR VPWR _9726_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9657_ _9830_/CLK _9657_/D _9731_/SET_B VGND VGND VPWR VPWR _9657_/Q sky130_fd_sc_hd__dfrtp_1
X_6869_ _9675_/Q VGND VGND VPWR VPWR _6869_/Y sky130_fd_sc_hd__inv_2
X_8608_ _8608_/A _8608_/B VGND VGND VPWR VPWR _8608_/Y sky130_fd_sc_hd__nor2_1
X_9588_ _9832_/CLK _9588_/D _9797_/SET_B VGND VGND VPWR VPWR _9588_/Q sky130_fd_sc_hd__dfstp_1
X_8539_ _8539_/A _8437_/X VGND VGND VPWR VPWR _8543_/C sky130_fd_sc_hd__or2b_1
XFILLER_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold580 _5641_/X VGND VGND VPWR VPWR _9341_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold591 _9702_/Q VGND VGND VPWR VPWR hold592/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8890_ _9657_/Q hold696/A _8971_/S VGND VGND VPWR VPWR _8890_/X sky130_fd_sc_hd__mux2_1
X_7910_ _7957_/A _8288_/B VGND VGND VPWR VPWR _8776_/A sky130_fd_sc_hd__nor2_2
X_7841_ _7876_/A _8674_/A VGND VGND VPWR VPWR _8068_/A sky130_fd_sc_hd__or2_4
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7772_ _9108_/Q _7772_/B VGND VGND VPWR VPWR _7772_/X sky130_fd_sc_hd__and2_1
X_4984_ _9134_/Q _9090_/Q _4971_/A _4981_/Y _4983_/X VGND VGND VPWR VPWR _9750_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_51_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9511_ _9514_/CLK _9511_/D _9571_/SET_B VGND VGND VPWR VPWR _9511_/Q sky130_fd_sc_hd__dfstp_1
X_6723_ _9822_/Q VGND VGND VPWR VPWR _6723_/Y sky130_fd_sc_hd__inv_4
XFILLER_176_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6654_ _9823_/Q VGND VGND VPWR VPWR _8823_/A sky130_fd_sc_hd__clkinv_8
X_9442_ _9791_/CLK _9442_/D _9817_/SET_B VGND VGND VPWR VPWR _9442_/Q sky130_fd_sc_hd__dfrtp_1
X_5605_ _9365_/Q _5600_/A hold612/X _5600_/Y VGND VGND VPWR VPWR _5605_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9373_ _9600_/CLK _9373_/D _9821_/SET_B VGND VGND VPWR VPWR _9373_/Q sky130_fd_sc_hd__dfstp_1
X_6585_ _6580_/Y _4525_/B _6581_/Y _5282_/B _6584_/X VGND VGND VPWR VPWR _6598_/B
+ sky130_fd_sc_hd__o221a_1
X_5536_ _9412_/Q _5534_/A hold510/X _5534_/Y VGND VGND VPWR VPWR _5536_/X sky130_fd_sc_hd__a22o_1
X_8324_ _8667_/A _8324_/B _8324_/C VGND VGND VPWR VPWR _8372_/B sky130_fd_sc_hd__and3_1
X_8255_ _8255_/A _8255_/B VGND VGND VPWR VPWR _8353_/B sky130_fd_sc_hd__or2_1
XFILLER_145_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5467_ _5467_/A VGND VGND VPWR VPWR _5468_/A sky130_fd_sc_hd__clkbuf_2
X_7206_ _6681_/Y _7182_/X _6723_/Y _7183_/X VGND VGND VPWR VPWR _7206_/X sky130_fd_sc_hd__o22a_1
XFILLER_87_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8186_ _8027_/Y _8432_/B _8185_/X VGND VGND VPWR VPWR _8186_/X sky130_fd_sc_hd__a21o_1
X_5398_ _5398_/A VGND VGND VPWR VPWR _5399_/A sky130_fd_sc_hd__clkbuf_2
X_7137_ _7137_/A VGND VGND VPWR VPWR _7137_/X sky130_fd_sc_hd__buf_4
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7068_ _7068_/A _9289_/Q VGND VGND VPWR VPWR _7129_/B sky130_fd_sc_hd__or2_2
X_6019_ _6053_/C _6015_/B _6015_/Y VGND VGND VPWR VPWR _9132_/D sky130_fd_sc_hd__a21oi_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9709_ _9730_/CLK _9709_/D _9730_/SET_B VGND VGND VPWR VPWR _9709_/Q sky130_fd_sc_hd__dfstp_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6370_ _6365_/Y _4865_/X _6366_/Y _5513_/B _6369_/X VGND VGND VPWR VPWR _6383_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5321_ _5474_/A _5321_/B VGND VGND VPWR VPWR _5322_/A sky130_fd_sc_hd__or2_1
X_8040_ _8040_/A VGND VGND VPWR VPWR _8158_/A sky130_fd_sc_hd__buf_6
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5252_ _5252_/A VGND VGND VPWR VPWR _5252_/X sky130_fd_sc_hd__clkbuf_1
X_5183_ _9650_/Q _5181_/A hold510/X _5181_/Y VGND VGND VPWR VPWR _5183_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8942_ _9759_/Q _6176_/Y _8999_/S VGND VGND VPWR VPWR _8942_/X sky130_fd_sc_hd__mux2_1
X_8873_ _6575_/Y input2/X input1/X VGND VGND VPWR VPWR _8873_/X sky130_fd_sc_hd__mux2_4
X_7824_ _7942_/C _7860_/A _7823_/X VGND VGND VPWR VPWR _8570_/B sky130_fd_sc_hd__o21ai_2
XFILLER_36_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4967_ _7039_/A VGND VGND VPWR VPWR _6024_/B sky130_fd_sc_hd__inv_2
X_7755_ _9130_/Q _7754_/B _7754_/Y VGND VGND VPWR VPWR _7755_/X sky130_fd_sc_hd__o21a_1
X_4898_ _6142_/A _4898_/B VGND VGND VPWR VPWR _5133_/B sky130_fd_sc_hd__or2_4
X_6706_ _9765_/Q VGND VGND VPWR VPWR _6706_/Y sky130_fd_sc_hd__clkinv_4
X_7686_ _6669_/Y _7507_/X _6736_/Y _7508_/X _7685_/X VGND VGND VPWR VPWR _7693_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9425_ _9574_/CLK _9425_/D _9571_/SET_B VGND VGND VPWR VPWR _9425_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6637_ _9560_/Q VGND VGND VPWR VPWR _6637_/Y sky130_fd_sc_hd__clkinv_2
X_9356_ _9391_/CLK _9356_/D _9563_/SET_B VGND VGND VPWR VPWR _9356_/Q sky130_fd_sc_hd__dfrtp_1
X_6568_ _9151_/Q VGND VGND VPWR VPWR _7735_/A sky130_fd_sc_hd__inv_4
XFILLER_118_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5519_ _9423_/Q _5515_/A _6067_/B1 _5515_/Y VGND VGND VPWR VPWR _5519_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8307_ _8307_/A _8687_/B VGND VGND VPWR VPWR _8309_/A sky130_fd_sc_hd__or2_1
X_6499_ _9197_/Q VGND VGND VPWR VPWR _6499_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9287_ _9322_/CLK _9287_/D _9797_/SET_B VGND VGND VPWR VPWR _9287_/Q sky130_fd_sc_hd__dfstp_4
X_8238_ _8388_/A _8388_/B _8237_/X VGND VGND VPWR VPWR _8625_/C sky130_fd_sc_hd__o21ai_2
XFILLER_133_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8169_ _8169_/A _8682_/B VGND VGND VPWR VPWR _8718_/A sky130_fd_sc_hd__nor2_1
XFILLER_120_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater407 _9571_/SET_B VGND VGND VPWR VPWR _9537_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_77_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5870_ _9225_/Q _5868_/A hold510/X _5868_/Y VGND VGND VPWR VPWR _9225_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4821_ _4813_/Y _4585_/B _4814_/Y _5263_/B _4820_/X VGND VGND VPWR VPWR _4852_/A
+ sky130_fd_sc_hd__o221a_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7540_ _6806_/Y _7497_/X _7537_/X _7539_/X VGND VGND VPWR VPWR _7550_/C sky130_fd_sc_hd__o211a_1
X_4752_ _4752_/A _5771_/B VGND VGND VPWR VPWR _4752_/X sky130_fd_sc_hd__or2_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4683_ _4913_/A _4764_/B VGND VGND VPWR VPWR _5581_/B sky130_fd_sc_hd__or2_4
X_7471_ _7471_/A _7479_/C _7471_/C VGND VGND VPWR VPWR _7520_/A sky130_fd_sc_hd__or3_2
X_9210_ _9212_/CLK _9210_/D _9797_/SET_B VGND VGND VPWR VPWR _9210_/Q sky130_fd_sc_hd__dfrtp_1
X_6422_ _9504_/Q VGND VGND VPWR VPWR _6422_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9141_ _9574_/CLK _9141_/D _9571_/SET_B VGND VGND VPWR VPWR _9141_/Q sky130_fd_sc_hd__dfrtp_1
X_6353_ _6353_/A VGND VGND VPWR VPWR _6353_/Y sky130_fd_sc_hd__inv_6
XFILLER_127_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5304_ _9569_/Q _5303_/A hold516/A _5303_/Y VGND VGND VPWR VPWR _5304_/X sky130_fd_sc_hd__a22o_1
X_9072_ _9718_/CLK _9072_/D VGND VGND VPWR VPWR _9072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6284_ _8864_/X _6282_/Y _6283_/Y _4863_/X VGND VGND VPWR VPWR _6284_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_130_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8023_ _8053_/A VGND VGND VPWR VPWR _8586_/A sky130_fd_sc_hd__clkinv_4
X_5235_ _6017_/A VGND VGND VPWR VPWR _5236_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5166_ _9661_/Q _5159_/A _8969_/A1 _5159_/Y VGND VGND VPWR VPWR _9661_/D sky130_fd_sc_hd__a22o_1
X_5097_ _9005_/X _9703_/Q _5101_/S VGND VGND VPWR VPWR _5098_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8925_ _7297_/Y _9680_/Q _9001_/S VGND VGND VPWR VPWR _8925_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8856_ _9833_/Q _6282_/Y _8975_/A1 _6282_/A _4473_/A VGND VGND VPWR VPWR _8856_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7807_ _7942_/C VGND VGND VPWR VPWR _7999_/A sky130_fd_sc_hd__inv_2
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5999_ _5999_/A VGND VGND VPWR VPWR _5999_/X sky130_fd_sc_hd__clkbuf_4
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8787_ _8787_/A VGND VGND VPWR VPWR _8788_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_169_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7738_ _7738_/A VGND VGND VPWR VPWR _7738_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9408_ _9695_/CLK _9408_/D _9689_/SET_B VGND VGND VPWR VPWR _9408_/Q sky130_fd_sc_hd__dfrtp_1
X_7669_ _6929_/Y _7515_/X _6864_/Y _7516_/X VGND VGND VPWR VPWR _7669_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9339_ _9643_/CLK _9339_/D _9689_/SET_B VGND VGND VPWR VPWR _9339_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput290 _8858_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_2
XFILLER_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold409 _5514_/X VGND VGND VPWR VPWR hold410/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5020_/A VGND VGND VPWR VPWR _9741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8710_ _8710_/A _8710_/B _8710_/C _8710_/D VGND VGND VPWR VPWR _8741_/D sky130_fd_sc_hd__or4_2
XFILLER_93_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6971_ _9697_/Q VGND VGND VPWR VPWR _6971_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_65_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9690_ _9694_/CLK _9690_/D _9689_/SET_B VGND VGND VPWR VPWR _9690_/Q sky130_fd_sc_hd__dfrtp_1
X_5922_ _5889_/A _8920_/X _8960_/X _9183_/Q VGND VGND VPWR VPWR _9183_/D sky130_fd_sc_hd__o22a_1
X_5853_ _9236_/Q _5849_/A hold53/X _5849_/Y VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_15_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9318_/CLK sky130_fd_sc_hd__clkbuf_16
X_8641_ _8641_/A _8641_/B _8641_/C _8641_/D VGND VGND VPWR VPWR _8738_/A sky130_fd_sc_hd__or4_4
XFILLER_61_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8572_ _8514_/Y _8570_/Y _8560_/X _8501_/C VGND VGND VPWR VPWR _8656_/D sky130_fd_sc_hd__a31o_1
X_4804_ _4804_/A VGND VGND VPWR VPWR _6353_/A sky130_fd_sc_hd__buf_12
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5784_ _5784_/A VGND VGND VPWR VPWR _5784_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7523_ _6910_/Y _7521_/X _6856_/Y _7522_/X VGND VGND VPWR VPWR _7523_/X sky130_fd_sc_hd__o22a_1
X_4735_ _7336_/A _5658_/B _4733_/Y _5818_/B VGND VGND VPWR VPWR _4735_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7454_ _7477_/A _7476_/B _7471_/C VGND VGND VPWR VPWR _7503_/A sky130_fd_sc_hd__or3_2
X_4666_ _4666_/A VGND VGND VPWR VPWR _4666_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4597_ _4643_/A _4898_/B VGND VGND VPWR VPWR _4598_/B sky130_fd_sc_hd__or2_4
X_7385_ _7385_/A _7385_/B _7385_/C VGND VGND VPWR VPWR _7385_/Y sky130_fd_sc_hd__nand3_2
X_6405_ _9272_/Q VGND VGND VPWR VPWR _6405_/Y sky130_fd_sc_hd__inv_2
X_6336_ _6334_/Y _4865_/X _6335_/Y _5935_/B VGND VGND VPWR VPWR _6336_/X sky130_fd_sc_hd__o22a_1
X_9124_ _9751_/CLK _9124_/D _6047_/X VGND VGND VPWR VPWR _9124_/Q sky130_fd_sc_hd__dfrtp_4
X_9055_ _9718_/CLK _9055_/D VGND VGND VPWR VPWR _9055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6267_ _6267_/A _6267_/B _6267_/C _6267_/D VGND VGND VPWR VPWR _6268_/D sky130_fd_sc_hd__and4_2
X_8006_ _8006_/A _8006_/B _8006_/C VGND VGND VPWR VPWR _8144_/B sky130_fd_sc_hd__or3_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6198_ _6194_/Y _5609_/B _6195_/Y _5482_/B _6197_/Y VGND VGND VPWR VPWR _6205_/C
+ sky130_fd_sc_hd__o221a_1
X_5218_ _9626_/Q _5216_/Y _8973_/X _5216_/A VGND VGND VPWR VPWR _9626_/D sky130_fd_sc_hd__o22a_1
XFILLER_69_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5149_ _9671_/Q _5146_/A _8965_/A1 _5146_/Y VGND VGND VPWR VPWR _9671_/D sky130_fd_sc_hd__a22o_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8908_ _8907_/X _9214_/Q _9096_/Q VGND VGND VPWR VPWR _8908_/X sky130_fd_sc_hd__mux2_1
X_8839_ _8839_/A VGND VGND VPWR VPWR _8840_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_40_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4520_ _9821_/Q _4513_/A _8969_/A1 _4513_/Y VGND VGND VPWR VPWR _9821_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold206 hold206/A VGND VGND VPWR VPWR hold207/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold217 hold217/A VGND VGND VPWR VPWR hold217/X sky130_fd_sc_hd__buf_12
Xhold239 _5580_/X VGND VGND VPWR VPWR hold240/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold228/A VGND VGND VPWR VPWR hold229/A sky130_fd_sc_hd__dlygate4sd3_1
X_7170_ _6951_/Y _7071_/D _6824_/Y _7166_/X _7169_/X VGND VGND VPWR VPWR _7186_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ _9447_/Q VGND VGND VPWR VPWR _6121_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_112_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6052_/A VGND VGND VPWR VPWR _6052_/X sky130_fd_sc_hd__clkbuf_1
X_5003_ _5017_/A VGND VGND VPWR VPWR _5004_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9811_ _9817_/CLK _9811_/D _7042_/B VGND VGND VPWR VPWR _9811_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6954_ _6952_/Y _5036_/B _6953_/Y _5946_/B VGND VGND VPWR VPWR _6954_/X sky130_fd_sc_hd__o22a_1
X_9742_ _9751_/CLK _9742_/D _5010_/X VGND VGND VPWR VPWR _9742_/Q sky130_fd_sc_hd__dfrtp_1
X_5905_ _9200_/Q _5904_/A hold516/X _5904_/Y VGND VGND VPWR VPWR _9200_/D sky130_fd_sc_hd__a22o_1
X_9673_ _9673_/CLK _9673_/D _9797_/SET_B VGND VGND VPWR VPWR _9673_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8624_ _8624_/A _8624_/B VGND VGND VPWR VPWR _8688_/B sky130_fd_sc_hd__or2_1
X_6885_ _9545_/Q VGND VGND VPWR VPWR _6885_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5836_ _9246_/Q _5828_/A _8975_/A1 _5828_/Y VGND VGND VPWR VPWR _9246_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8555_ _8555_/A VGND VGND VPWR VPWR _8555_/X sky130_fd_sc_hd__clkbuf_1
X_5767_ _9097_/Q _7128_/A _7129_/A _5765_/A _5741_/Y VGND VGND VPWR VPWR _5768_/A
+ sky130_fd_sc_hd__a32o_1
X_8486_ _8486_/A _8486_/B VGND VGND VPWR VPWR _8490_/B sky130_fd_sc_hd__or2_1
X_7506_ _6950_/Y _7497_/X _7499_/X _7505_/X VGND VGND VPWR VPWR _7532_/C sky130_fd_sc_hd__o211a_1
X_5698_ _5698_/A _5698_/B VGND VGND VPWR VPWR _5699_/A sky130_fd_sc_hd__or2_1
X_4718_ _4718_/A VGND VGND VPWR VPWR _6196_/A sky130_fd_sc_hd__buf_8
XFILLER_162_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4649_ _7042_/B VGND VGND VPWR VPWR _6083_/B sky130_fd_sc_hd__inv_2
X_7437_ _7479_/A _9293_/Q _7476_/B _7471_/C VGND VGND VPWR VPWR _7487_/A sky130_fd_sc_hd__or4_4
XFILLER_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7368_ _6713_/Y _7144_/X _6803_/Y _7145_/X _7367_/X VGND VGND VPWR VPWR _7375_/A
+ sky130_fd_sc_hd__o221a_1
X_9107_ _9705_/CLK _9107_/D _6177_/A VGND VGND VPWR VPWR _9107_/Q sky130_fd_sc_hd__dfrtp_1
X_6319_ _9251_/Q VGND VGND VPWR VPWR _6319_/Y sky130_fd_sc_hd__clkinv_2
X_7299_ _6170_/Y _7137_/X _6164_/Y _7138_/X _7298_/X VGND VGND VPWR VPWR _7299_/X
+ sky130_fd_sc_hd__o221a_1
X_9038_ _9606_/Q _8811_/A VGND VGND VPWR VPWR _9038_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_89_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6670_ _9262_/Q VGND VGND VPWR VPWR _6670_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5621_ _5621_/A VGND VGND VPWR VPWR _5622_/A sky130_fd_sc_hd__clkbuf_2
X_8340_ _8340_/A VGND VGND VPWR VPWR _8642_/A sky130_fd_sc_hd__inv_2
X_5552_ _5552_/A VGND VGND VPWR VPWR _5552_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4503_ hold136/X _9830_/Q _6049_/S VGND VGND VPWR VPWR _4504_/A sky130_fd_sc_hd__mux2_1
X_8271_ _8277_/A _8274_/B VGND VGND VPWR VPWR _8700_/B sky130_fd_sc_hd__nor2_1
X_5483_ _5483_/A VGND VGND VPWR VPWR _5484_/A sky130_fd_sc_hd__buf_2
XFILLER_132_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7222_ _8805_/A _7167_/X _7731_/A _7168_/X VGND VGND VPWR VPWR _7222_/X sky130_fd_sc_hd__o22a_1
X_7153_ _6885_/Y _7151_/X _6863_/Y _7152_/X VGND VGND VPWR VPWR _7153_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6104_ _9543_/Q VGND VGND VPWR VPWR _6104_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7084_ _7113_/A _7129_/B _7084_/C VGND VGND VPWR VPWR _7161_/A sky130_fd_sc_hd__or3_4
XFILLER_112_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6035_ _6035_/A VGND VGND VPWR VPWR _6035_/X sky130_fd_sc_hd__clkbuf_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7986_ _8421_/D _8421_/B _8120_/C VGND VGND VPWR VPWR _7987_/A sky130_fd_sc_hd__or3_1
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9725_ _9729_/CLK _9725_/D _9727_/SET_B VGND VGND VPWR VPWR _9725_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6937_ _6935_/Y _5551_/B _6936_/Y _6112_/B VGND VGND VPWR VPWR _6937_/X sky130_fd_sc_hd__o22a_1
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9656_ _9830_/CLK _9656_/D _9731_/SET_B VGND VGND VPWR VPWR _9656_/Q sky130_fd_sc_hd__dfrtp_1
X_6868_ _9670_/Q VGND VGND VPWR VPWR _6868_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8607_ _8607_/A _8682_/B VGND VGND VPWR VPWR _8762_/B sky130_fd_sc_hd__nor2_1
X_9587_ _9827_/CLK _9587_/D _9797_/SET_B VGND VGND VPWR VPWR _9587_/Q sky130_fd_sc_hd__dfrtp_1
X_5819_ _5819_/A VGND VGND VPWR VPWR _5820_/A sky130_fd_sc_hd__clkbuf_2
X_8538_ _8538_/A _8538_/B VGND VGND VPWR VPWR _8737_/C sky130_fd_sc_hd__nor2_1
X_6799_ _9792_/Q VGND VGND VPWR VPWR _6799_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8469_ _8469_/A _8643_/D VGND VGND VPWR VPWR _8470_/B sky130_fd_sc_hd__or2_1
XFILLER_163_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold570 _5243_/X VGND VGND VPWR VPWR _9609_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_150_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold581 _5938_/X VGND VGND VPWR VPWR _9174_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold592 hold592/A VGND VGND VPWR VPWR hold592/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput190 wb_dat_i[3] VGND VGND VPWR VPWR _9006_/A1 sky130_fd_sc_hd__clkbuf_1
X_7840_ _8421_/C _7996_/B _8421_/B VGND VGND VPWR VPWR _8674_/A sky130_fd_sc_hd__or3_4
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7771_ _9110_/Q _7771_/A2 _9109_/Q _7771_/B2 _7770_/X VGND VGND VPWR VPWR _7771_/X
+ sky130_fd_sc_hd__a221o_1
X_4983_ _6053_/A _6053_/B _6053_/C _9750_/Q VGND VGND VPWR VPWR _4983_/X sky130_fd_sc_hd__o31a_1
X_9510_ _9514_/CLK _9510_/D _9571_/SET_B VGND VGND VPWR VPWR _9510_/Q sky130_fd_sc_hd__dfstp_1
X_6722_ _6722_/A _6722_/B _6722_/C _6722_/D VGND VGND VPWR VPWR _6816_/B sky130_fd_sc_hd__and4_1
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6653_ _9565_/Q VGND VGND VPWR VPWR _8829_/A sky130_fd_sc_hd__inv_8
X_9441_ _9798_/CLK _9441_/D _9817_/SET_B VGND VGND VPWR VPWR _9441_/Q sky130_fd_sc_hd__dfstp_1
X_5604_ _9366_/Q _5600_/A hold53/X _5600_/Y VGND VGND VPWR VPWR _5604_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9372_ _9431_/CLK _9372_/D _9821_/SET_B VGND VGND VPWR VPWR _9372_/Q sky130_fd_sc_hd__dfrtp_1
X_6584_ _6582_/Y _5123_/B _6583_/Y _4915_/X VGND VGND VPWR VPWR _6584_/X sky130_fd_sc_hd__o22a_1
X_5535_ _9413_/Q _5534_/A hold516/X _5534_/Y VGND VGND VPWR VPWR _5535_/X sky130_fd_sc_hd__a22o_1
X_8323_ _8720_/A _8323_/B VGND VGND VPWR VPWR _8325_/A sky130_fd_sc_hd__or2_1
XFILLER_145_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8254_ _8383_/B _8302_/B _8354_/D VGND VGND VPWR VPWR _8266_/B sky130_fd_sc_hd__o21ai_1
X_5466_ _5474_/A _5466_/B VGND VGND VPWR VPWR _5467_/A sky130_fd_sc_hd__or2_1
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7205_ _6794_/Y _5756_/X _6704_/Y _7071_/A _7204_/X VGND VGND VPWR VPWR _7208_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8185_ _8185_/A _8404_/A _8617_/A _8669_/B VGND VGND VPWR VPWR _8185_/X sky130_fd_sc_hd__or4_1
X_5397_ _5474_/A _5397_/B VGND VGND VPWR VPWR _5398_/A sky130_fd_sc_hd__or2_1
XFILLER_98_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7136_ _7136_/A VGND VGND VPWR VPWR _7136_/X sky130_fd_sc_hd__buf_4
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7067_ _7067_/A VGND VGND VPWR VPWR _7071_/C sky130_fd_sc_hd__buf_4
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6018_ _6018_/A VGND VGND VPWR VPWR _6018_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7969_ _7887_/A _8229_/A _7968_/Y VGND VGND VPWR VPWR _7970_/B sky130_fd_sc_hd__o21ba_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9708_ _4471_/A1 _9708_/D _6177_/A VGND VGND VPWR VPWR _9708_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9639_ _9643_/CLK _9639_/D _9689_/SET_B VGND VGND VPWR VPWR _9639_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5320_ _9557_/Q _5315_/A _6008_/B1 _5315_/Y VGND VGND VPWR VPWR _9557_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5251_ _6067_/B1 _9602_/Q _5251_/S VGND VGND VPWR VPWR _5252_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5182_ _9651_/Q _5181_/A hold516/X _5181_/Y VGND VGND VPWR VPWR _5182_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8941_ _7755_/X _9129_/Q _9093_/Q VGND VGND VPWR VPWR _8941_/X sky130_fd_sc_hd__mux2_1
X_8872_ _9635_/Q input91/X _8877_/S VGND VGND VPWR VPWR _8872_/X sky130_fd_sc_hd__mux2_1
X_7823_ _7999_/A _7823_/B VGND VGND VPWR VPWR _7823_/X sky130_fd_sc_hd__or2_1
XFILLER_169_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7754_ _9130_/Q _7754_/B VGND VGND VPWR VPWR _7754_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6705_ _9203_/Q VGND VGND VPWR VPWR _6705_/Y sky130_fd_sc_hd__inv_2
X_4966_ _4966_/A VGND VGND VPWR VPWR _7039_/A sky130_fd_sc_hd__buf_2
XFILLER_149_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7685_ _6726_/Y _7509_/X _6731_/Y _7510_/X VGND VGND VPWR VPWR _7685_/X sky130_fd_sc_hd__o22a_1
X_4897_ _9674_/Q VGND VGND VPWR VPWR _4897_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9424_ _9574_/CLK _9424_/D _9571_/SET_B VGND VGND VPWR VPWR _9424_/Q sky130_fd_sc_hd__dfstp_1
X_6636_ _9443_/Q VGND VGND VPWR VPWR _8811_/A sky130_fd_sc_hd__inv_8
XFILLER_192_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9355_ _9391_/CLK _9355_/D _9689_/SET_B VGND VGND VPWR VPWR _9355_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_164_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6567_ _6562_/Y _6353_/A _7731_/A _5902_/B _6566_/X VGND VGND VPWR VPWR _6567_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5518_ _9424_/Q _5515_/A hold217/X _5515_/Y VGND VGND VPWR VPWR _9424_/D sky130_fd_sc_hd__a22o_1
X_8306_ _8366_/A _8306_/B VGND VGND VPWR VPWR _8687_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6498_ _9231_/Q VGND VGND VPWR VPWR _6498_/Y sky130_fd_sc_hd__inv_2
X_9286_ _9729_/CLK _9286_/D _9727_/SET_B VGND VGND VPWR VPWR _9286_/Q sky130_fd_sc_hd__dfrtp_1
X_8237_ _7942_/C _8236_/Y _7876_/A _8000_/Y VGND VGND VPWR VPWR _8237_/X sky130_fd_sc_hd__a2bb2o_1
X_5449_ _9471_/Q _5445_/X hold577/A _5446_/Y VGND VGND VPWR VPWR _5449_/X sky130_fd_sc_hd__a22o_1
XFILLER_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8168_ _8396_/A _8168_/B _8613_/A _8725_/B VGND VGND VPWR VPWR _8172_/A sky130_fd_sc_hd__or4_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7119_ _4763_/Y _7167_/A _4688_/Y _7168_/A VGND VGND VPWR VPWR _7119_/X sky130_fd_sc_hd__o22a_1
X_8099_ _8563_/B VGND VGND VPWR VPWR _8102_/A sky130_fd_sc_hd__inv_2
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater408 _9727_/SET_B VGND VGND VPWR VPWR _9571_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_93_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4820_ _4817_/Y _5144_/B _4819_/Y _4634_/B VGND VGND VPWR VPWR _4820_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4922_/B _4801_/B VGND VGND VPWR VPWR _5771_/B sky130_fd_sc_hd__or2_4
XFILLER_147_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4682_ _4685_/B _4685_/C _4682_/C VGND VGND VPWR VPWR _4732_/B sky130_fd_sc_hd__or3_4
X_7470_ _7471_/A _7478_/C _9297_/Q VGND VGND VPWR VPWR _7519_/A sky130_fd_sc_hd__or3_2
XFILLER_186_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6421_ _9514_/Q VGND VGND VPWR VPWR _6421_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9140_ _9577_/CLK _9140_/D _9571_/SET_B VGND VGND VPWR VPWR _9140_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6352_ _9411_/Q VGND VGND VPWR VPWR _6352_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5303_ _5303_/A VGND VGND VPWR VPWR _5303_/Y sky130_fd_sc_hd__inv_2
X_9071_ _9718_/CLK _9071_/D VGND VGND VPWR VPWR _9071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6283_ _6283_/A VGND VGND VPWR VPWR _6283_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_142_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5234_ _9612_/Q _5226_/Y _8966_/X _5226_/A VGND VGND VPWR VPWR _5234_/X sky130_fd_sc_hd__o22a_1
X_8022_ _8190_/B VGND VGND VPWR VPWR _8594_/A sky130_fd_sc_hd__buf_2
XFILLER_88_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5165_ _9662_/Q _5159_/A _8965_/A1 _5159_/Y VGND VGND VPWR VPWR _9662_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5096_ _5096_/A VGND VGND VPWR VPWR _9704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8924_ _8923_/X _9184_/Q _9096_/Q VGND VGND VPWR VPWR _8924_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8855_ _8855_/A _8855_/B VGND VGND VPWR VPWR _9102_/D sky130_fd_sc_hd__nor2_1
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7806_ _7806_/A _7806_/B _7806_/C _7806_/D VGND VGND VPWR VPWR _7810_/C sky130_fd_sc_hd__nand4_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _6083_/A _5998_/B VGND VGND VPWR VPWR _5998_/X sky130_fd_sc_hd__or2_1
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8786_ _8786_/A VGND VGND VPWR VPWR _8786_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4949_ _4949_/A _4953_/B VGND VGND VPWR VPWR _5329_/B sky130_fd_sc_hd__or2_4
X_7737_ _7737_/A VGND VGND VPWR VPWR _7738_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7668_ _6966_/Y _7507_/X _6855_/Y _7508_/X _7667_/X VGND VGND VPWR VPWR _7675_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9407_ _9695_/CLK _9407_/D _9689_/SET_B VGND VGND VPWR VPWR _9407_/Q sky130_fd_sc_hd__dfstp_1
X_6619_ _9547_/Q VGND VGND VPWR VPWR _8819_/A sky130_fd_sc_hd__inv_8
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7599_ _6319_/Y _7521_/X _6275_/Y _7522_/X VGND VGND VPWR VPWR _7599_/X sky130_fd_sc_hd__o22a_1
XFILLER_125_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9338_ _9695_/CLK _9338_/D _9689_/SET_B VGND VGND VPWR VPWR _9338_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9269_ _9431_/CLK _9269_/D _9817_/SET_B VGND VGND VPWR VPWR _9269_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput280 _9026_/Z VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_2
Xoutput291 _7048_/Y VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_2
XFILLER_59_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6970_ _9274_/Q VGND VGND VPWR VPWR _6970_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5921_ _5889_/A _8922_/X _8960_/X _9184_/Q VGND VGND VPWR VPWR _9184_/D sky130_fd_sc_hd__o22a_1
XFILLER_80_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5852_ _9237_/Q _5849_/A hold696/A _5849_/Y VGND VGND VPWR VPWR _5852_/X sky130_fd_sc_hd__a22o_1
X_8640_ _8737_/D _8701_/C _8769_/A _8699_/D VGND VGND VPWR VPWR _8643_/A sky130_fd_sc_hd__or4_2
XFILLER_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8571_ _8565_/Y _8570_/Y _8560_/X _8497_/B VGND VGND VPWR VPWR _8776_/D sky130_fd_sc_hd__a31o_1
X_4803_ _4803_/A _4920_/A VGND VGND VPWR VPWR _4804_/A sky130_fd_sc_hd__or2_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5783_ _7028_/A _5669_/Y _5741_/Y _5782_/X VGND VGND VPWR VPWR _5784_/A sky130_fd_sc_hd__a31o_1
XFILLER_34_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4734_ _4941_/A _4801_/B VGND VGND VPWR VPWR _5818_/B sky130_fd_sc_hd__or2_4
XFILLER_21_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7522_ _7522_/A VGND VGND VPWR VPWR _7522_/X sky130_fd_sc_hd__buf_6
XFILLER_159_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7453_ _7460_/A _7478_/C _7478_/D VGND VGND VPWR VPWR _7502_/A sky130_fd_sc_hd__or3_2
X_4665_ _4969_/A VGND VGND VPWR VPWR _4666_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_174_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4596_ _4689_/A _4750_/D _4750_/A _4708_/B VGND VGND VPWR VPWR _4869_/A sky130_fd_sc_hd__or4_4
X_7384_ _7384_/A _7384_/B _7384_/C _7384_/D VGND VGND VPWR VPWR _7385_/C sky130_fd_sc_hd__and4_1
X_6404_ _9258_/Q VGND VGND VPWR VPWR _6404_/Y sky130_fd_sc_hd__clkinv_2
X_9123_ _9830_/CLK _9123_/D _9537_/SET_B VGND VGND VPWR VPWR _9123_/Q sky130_fd_sc_hd__dfrtp_2
X_6335_ _9172_/Q VGND VGND VPWR VPWR _6335_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_130_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9054_ _9718_/CLK _9054_/D VGND VGND VPWR VPWR _9054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8005_ _8005_/A _8132_/B VGND VGND VPWR VPWR _8011_/A sky130_fd_sc_hd__or2_2
XFILLER_103_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6266_ _6261_/Y _4865_/X _6262_/Y _5133_/B _6265_/X VGND VGND VPWR VPWR _6267_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6197_ input69/X _8973_/S input50/X _8975_/S VGND VGND VPWR VPWR _6197_/Y sky130_fd_sc_hd__a22oi_4
X_5217_ _9627_/Q _5216_/Y _8944_/X _5216_/A VGND VGND VPWR VPWR _9627_/D sky130_fd_sc_hd__o22a_1
XFILLER_69_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5148_ _9672_/Q _5146_/A _8964_/A1 _5146_/Y VGND VGND VPWR VPWR _9672_/D sky130_fd_sc_hd__a22o_1
X_5079_ _7765_/A _7766_/A _8852_/A VGND VGND VPWR VPWR _5085_/A sky130_fd_sc_hd__a21oi_1
XFILLER_178_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8907_ _7676_/Y _9670_/Q _9020_/S VGND VGND VPWR VPWR _8907_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8838_ _8838_/A VGND VGND VPWR VPWR _8838_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8769_ _8769_/A _8769_/B _8769_/C _8769_/D VGND VGND VPWR VPWR _8770_/A sky130_fd_sc_hd__or4_1
XFILLER_12_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold207 hold207/A VGND VGND VPWR VPWR _9364_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold229 hold229/A VGND VGND VPWR VPWR _9432_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_144_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold218 _5386_/X VGND VGND VPWR VPWR hold219/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6120_ _6114_/Y _5263_/B _6115_/Y _4611_/B _6119_/X VGND VGND VPWR VPWR _6127_/C
+ sky130_fd_sc_hd__o221a_4
XFILLER_140_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6071_/A VGND VGND VPWR VPWR _6052_/A sky130_fd_sc_hd__clkbuf_1
X_5002_ hold36/A _4989_/A _9744_/Q _4989_/Y VGND VGND VPWR VPWR _9745_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9810_ _9810_/CLK _9810_/D _7042_/B VGND VGND VPWR VPWR _9810_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9741_ _8879_/A1 _9741_/D _5018_/X VGND VGND VPWR VPWR _9741_/Q sky130_fd_sc_hd__dfrtp_1
X_6953_ _9163_/Q VGND VGND VPWR VPWR _6953_/Y sky130_fd_sc_hd__clkinv_4
X_6884_ _9493_/Q VGND VGND VPWR VPWR _6884_/Y sky130_fd_sc_hd__clkinv_4
X_5904_ _5904_/A VGND VGND VPWR VPWR _5904_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9672_ _9832_/CLK _9672_/D _9797_/SET_B VGND VGND VPWR VPWR _9672_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8623_ _8045_/A _8321_/C _8322_/B VGND VGND VPWR VPWR _8624_/B sky130_fd_sc_hd__o21ai_1
X_5835_ _9247_/Q _5828_/A _8969_/A1 _5828_/Y VGND VGND VPWR VPWR _9247_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8554_ _8645_/A _8554_/B _8645_/C _8554_/D VGND VGND VPWR VPWR _8555_/A sky130_fd_sc_hd__or4_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5766_ _9288_/Q _5766_/B VGND VGND VPWR VPWR _7129_/A sky130_fd_sc_hd__or2_2
X_8485_ _7941_/B _8666_/B _7935_/X VGND VGND VPWR VPWR _8486_/B sky130_fd_sc_hd__o21ai_1
X_7505_ _6830_/Y _7500_/X _6891_/Y _7501_/X _7504_/X VGND VGND VPWR VPWR _7505_/X
+ sky130_fd_sc_hd__o221a_1
X_5697_ _9311_/Q _5689_/A hold601/A _5689_/Y VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__a22o_1
X_4717_ _4803_/A _4925_/B VGND VGND VPWR VPWR _4718_/A sky130_fd_sc_hd__or2_1
X_4648_ _4648_/A VGND VGND VPWR VPWR _4648_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7436_ _9296_/Q _7436_/B VGND VGND VPWR VPWR _7476_/B sky130_fd_sc_hd__or2_2
XFILLER_162_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9106_ _4471_/A1 _9106_/D _6177_/A VGND VGND VPWR VPWR _9106_/Q sky130_fd_sc_hd__dfrtp_1
X_7367_ _6763_/Y _7067_/A _6774_/Y _7146_/X VGND VGND VPWR VPWR _7367_/X sky130_fd_sc_hd__o22a_1
X_4579_ _5250_/A _4579_/B VGND VGND VPWR VPWR _4582_/S sky130_fd_sc_hd__or2_1
X_6318_ _9385_/Q VGND VGND VPWR VPWR _6318_/Y sky130_fd_sc_hd__inv_2
X_7298_ _6144_/Y _7139_/X _6105_/Y _7140_/X VGND VGND VPWR VPWR _7298_/X sky130_fd_sc_hd__o22a_1
XFILLER_89_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9037_ _9605_/Q _8809_/A VGND VGND VPWR VPWR _9037_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6249_ _9154_/Q VGND VGND VPWR VPWR _6249_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_14_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9576_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold90 hold90/A VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_29_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9416_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5620_ _5698_/A _5620_/B VGND VGND VPWR VPWR _5621_/A sky130_fd_sc_hd__or2_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5551_ _5698_/A _5551_/B VGND VGND VPWR VPWR _5551_/X sky130_fd_sc_hd__or2_1
X_4502_ _5250_/A _4502_/B VGND VGND VPWR VPWR _6049_/S sky130_fd_sc_hd__or2_2
X_8270_ _8272_/A _8306_/B VGND VGND VPWR VPWR _8718_/B sky130_fd_sc_hd__nor2_2
X_7221_ _7221_/A _7221_/B _7221_/C _7221_/D VGND VGND VPWR VPWR _7231_/B sky130_fd_sc_hd__and4_1
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5482_ _5570_/A _5482_/B VGND VGND VPWR VPWR _5483_/A sky130_fd_sc_hd__or2_1
XFILLER_144_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7152_ _7152_/A VGND VGND VPWR VPWR _7152_/X sky130_fd_sc_hd__buf_6
X_6103_ _9491_/Q VGND VGND VPWR VPWR _6103_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7083_ _7157_/A _7155_/A _7146_/A _7171_/A VGND VGND VPWR VPWR _7094_/B sky130_fd_sc_hd__and4_1
XFILLER_100_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6034_ _6071_/A VGND VGND VPWR VPWR _6035_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_100_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7985_ _8421_/C _8236_/A VGND VGND VPWR VPWR _8120_/C sky130_fd_sc_hd__or2_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6936_ _9433_/Q VGND VGND VPWR VPWR _6936_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9724_ _9751_/CLK _9724_/D _5056_/X VGND VGND VPWR VPWR _9724_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9655_ _9736_/CLK _9655_/D _9731_/SET_B VGND VGND VPWR VPWR _9655_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6867_ _6862_/Y _4844_/X _6863_/Y _5301_/B _6866_/X VGND VGND VPWR VPWR _6909_/A
+ sky130_fd_sc_hd__o221a_1
X_8606_ _8678_/A _8678_/B _8678_/C _8605_/X VGND VGND VPWR VPWR _8606_/X sky130_fd_sc_hd__or4b_1
X_9586_ _9600_/CLK _9586_/D _9821_/SET_B VGND VGND VPWR VPWR _9586_/Q sky130_fd_sc_hd__dfrtp_1
X_6798_ _9442_/Q VGND VGND VPWR VPWR _6798_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_22_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5818_ _5990_/A _5818_/B VGND VGND VPWR VPWR _5819_/A sky130_fd_sc_hd__or2_1
X_8537_ _8383_/A _8540_/A _7904_/D _7924_/X VGND VGND VPWR VPWR _8538_/B sky130_fd_sc_hd__o22a_1
X_5749_ _9289_/Q VGND VGND VPWR VPWR _7081_/B sky130_fd_sc_hd__inv_2
XFILLER_182_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8468_ _8518_/A _8581_/A VGND VGND VPWR VPWR _8643_/D sky130_fd_sc_hd__or2_2
XFILLER_190_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8399_ _8399_/A _8700_/B VGND VGND VPWR VPWR _8615_/C sky130_fd_sc_hd__or2_1
X_7419_ _7419_/A _7419_/B _7419_/C _7419_/D VGND VGND VPWR VPWR _7429_/B sky130_fd_sc_hd__and4_1
XFILLER_190_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold560 _5789_/X VGND VGND VPWR VPWR _9280_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold571 _5172_/X VGND VGND VPWR VPWR _9658_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold593 hold593/A VGND VGND VPWR VPWR hold593/X sky130_fd_sc_hd__buf_12
XFILLER_150_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold582 _5039_/X VGND VGND VPWR VPWR _9737_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput180 wb_dat_i[23] VGND VGND VPWR VPWR _7782_/B sky130_fd_sc_hd__clkbuf_1
Xinput191 wb_dat_i[4] VGND VGND VPWR VPWR _9007_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7770_ _9108_/Q _7770_/B VGND VGND VPWR VPWR _7770_/X sky130_fd_sc_hd__and2_1
X_4982_ _9090_/Q VGND VGND VPWR VPWR _6053_/B sky130_fd_sc_hd__clkinv_4
XFILLER_189_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6721_ _6721_/A _6721_/B _6721_/C _6721_/D VGND VGND VPWR VPWR _6722_/D sky130_fd_sc_hd__and4_1
XFILLER_189_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6652_ _9807_/Q VGND VGND VPWR VPWR _6652_/Y sky130_fd_sc_hd__inv_2
X_9440_ _9686_/CLK _9440_/D _9817_/SET_B VGND VGND VPWR VPWR _9440_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5603_ _9367_/Q _5600_/A hold696/A _5600_/Y VGND VGND VPWR VPWR _5603_/X sky130_fd_sc_hd__a22o_1
X_9371_ _9431_/CLK _9371_/D _9821_/SET_B VGND VGND VPWR VPWR _9371_/Q sky130_fd_sc_hd__dfrtp_1
X_8322_ _8317_/X _8322_/B _8322_/C VGND VGND VPWR VPWR _8323_/B sky130_fd_sc_hd__nand3b_1
X_6583_ _6583_/A VGND VGND VPWR VPWR _6583_/Y sky130_fd_sc_hd__inv_2
X_5534_ _5534_/A VGND VGND VPWR VPWR _5534_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5465_ _9458_/Q _5456_/X hold601/X _5457_/Y VGND VGND VPWR VPWR _5465_/X sky130_fd_sc_hd__a22o_1
X_8253_ _8383_/B _8306_/B VGND VGND VPWR VPWR _8354_/D sky130_fd_sc_hd__or2_2
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7204_ _7204_/A _7380_/B VGND VGND VPWR VPWR _7204_/X sky130_fd_sc_hd__or2_1
X_8184_ _8205_/A _8593_/A VGND VGND VPWR VPWR _8669_/B sky130_fd_sc_hd__nor2_1
X_5396_ _9505_/Q _5391_/A _6008_/B1 _5391_/Y VGND VGND VPWR VPWR _5396_/X sky130_fd_sc_hd__a22o_1
X_7135_ _7135_/A VGND VGND VPWR VPWR _7135_/X sky130_fd_sc_hd__buf_4
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7066_ _7121_/B _7084_/C VGND VGND VPWR VPWR _7067_/A sky130_fd_sc_hd__or2_4
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6017_ _6017_/A VGND VGND VPWR VPWR _6018_/A sky130_fd_sc_hd__clkbuf_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7968_ _7968_/A _7968_/B VGND VGND VPWR VPWR _7968_/Y sky130_fd_sc_hd__nand2_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9707_ _4471_/A1 _9707_/D _6177_/A VGND VGND VPWR VPWR _9707_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6919_ _6914_/Y _5858_/B _6915_/Y _5609_/B _6918_/X VGND VGND VPWR VPWR _6932_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7899_ _8557_/B _8304_/B VGND VGND VPWR VPWR _8709_/A sky130_fd_sc_hd__nor2_1
XFILLER_42_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9638_ _9643_/CLK _9638_/D _9689_/SET_B VGND VGND VPWR VPWR _9638_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9569_ _9569_/CLK _9569_/D _9563_/SET_B VGND VGND VPWR VPWR _9569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold390 hold390/A VGND VGND VPWR VPWR hold391/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5250_ _5250_/A _5250_/B VGND VGND VPWR VPWR _5251_/S sky130_fd_sc_hd__or2_1
XFILLER_114_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5181_ _5181_/A VGND VGND VPWR VPWR _5181_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8940_ _7739_/Y _5237_/A _9092_/Q VGND VGND VPWR VPWR _9100_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8871_ _9634_/Q input89/X _8877_/S VGND VGND VPWR VPWR _8871_/X sky130_fd_sc_hd__mux2_1
X_7822_ _7823_/B VGND VGND VPWR VPWR _7860_/A sky130_fd_sc_hd__inv_2
XFILLER_36_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4965_ _6053_/A _6053_/D _6053_/C VGND VGND VPWR VPWR _4966_/A sky130_fd_sc_hd__or3_1
X_7753_ _7753_/A VGND VGND VPWR VPWR _7754_/B sky130_fd_sc_hd__inv_2
X_6704_ _9137_/Q VGND VGND VPWR VPWR _6704_/Y sky130_fd_sc_hd__inv_2
X_9423_ _9574_/CLK _9423_/D _9571_/SET_B VGND VGND VPWR VPWR _9423_/Q sky130_fd_sc_hd__dfrtp_1
X_7684_ _6762_/Y _7497_/X _7681_/X _7683_/X VGND VGND VPWR VPWR _7694_/C sky130_fd_sc_hd__o211a_1
X_4896_ _9768_/Q VGND VGND VPWR VPWR _4896_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6635_ _9534_/Q VGND VGND VPWR VPWR _6635_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9354_ _9391_/CLK _9354_/D _9689_/SET_B VGND VGND VPWR VPWR _9354_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6566_ _6564_/Y _5103_/B _6565_/Y _6083_/C VGND VGND VPWR VPWR _6566_/X sky130_fd_sc_hd__o22a_2
XFILLER_164_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5517_ _9425_/Q _5515_/A _6065_/B1 _5515_/Y VGND VGND VPWR VPWR _5517_/X sky130_fd_sc_hd__a22o_1
X_9285_ _9729_/CLK _9285_/D _9727_/SET_B VGND VGND VPWR VPWR _9285_/Q sky130_fd_sc_hd__dfrtp_1
X_8305_ _8305_/A _8411_/B VGND VGND VPWR VPWR _8307_/A sky130_fd_sc_hd__or2_1
X_8236_ _8236_/A _8236_/B VGND VGND VPWR VPWR _8236_/Y sky130_fd_sc_hd__nor2_1
XFILLER_133_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6497_ _6492_/Y _5570_/B _6493_/Y _5036_/B _6496_/X VGND VGND VPWR VPWR _6504_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_172_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5448_ _9472_/Q _5446_/A hold510/X _5446_/Y VGND VGND VPWR VPWR _5448_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5379_ _5379_/A VGND VGND VPWR VPWR _5380_/A sky130_fd_sc_hd__clkbuf_4
X_8167_ _8179_/A _8169_/A VGND VGND VPWR VPWR _8725_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8098_ _8098_/A _8578_/A VGND VGND VPWR VPWR _8103_/A sky130_fd_sc_hd__nand2_1
XFILLER_120_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7118_ _9288_/Q _9287_/Q _7118_/C _7129_/C VGND VGND VPWR VPWR _7167_/A sky130_fd_sc_hd__or4_4
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7049_ _9668_/Q _7049_/B VGND VGND VPWR VPWR _7050_/A sky130_fd_sc_hd__and2b_1
XFILLER_47_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater409 _7042_/B VGND VGND VPWR VPWR _9727_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_93_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _4750_/A _4750_/B _4750_/C _4750_/D VGND VGND VPWR VPWR _4922_/B sky130_fd_sc_hd__or4_4
XFILLER_159_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4681_ _9375_/Q VGND VGND VPWR VPWR _4681_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_146_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6420_ _6415_/Y _4585_/B _6416_/Y _4929_/X _6419_/X VGND VGND VPWR VPWR _6439_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_174_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6351_ _9367_/Q VGND VGND VPWR VPWR _6351_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_161_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5302_ _5302_/A VGND VGND VPWR VPWR _5303_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_127_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9070_ _9705_/CLK _9070_/D VGND VGND VPWR VPWR _9070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6282_ _6282_/A VGND VGND VPWR VPWR _6282_/Y sky130_fd_sc_hd__inv_6
X_5233_ _9613_/Q _5226_/Y _8945_/X hold666/X VGND VGND VPWR VPWR _9613_/D sky130_fd_sc_hd__o22a_1
X_8021_ _8035_/B _8032_/B VGND VGND VPWR VPWR _8190_/B sky130_fd_sc_hd__or2_1
Xclkbuf_opt_3_0_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR clkbuf_leaf_8_csclk/A
+ sky130_fd_sc_hd__clkbuf_16
X_5164_ _9663_/Q _5159_/A _8964_/A1 _5159_/Y VGND VGND VPWR VPWR _9663_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5095_ _9006_/X _9704_/Q _5101_/S VGND VGND VPWR VPWR _5096_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8923_ _7275_/Y _9679_/Q _9001_/S VGND VGND VPWR VPWR _8923_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8854_ _8854_/A _8855_/B VGND VGND VPWR VPWR _9103_/D sky130_fd_sc_hd__nor2_1
X_7805_ _7805_/A _7805_/B VGND VGND VPWR VPWR _7810_/B sky130_fd_sc_hd__nand2_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8785_ _8785_/A VGND VGND VPWR VPWR _8786_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5997_ _9143_/Q _5992_/A _8975_/A1 _5992_/Y VGND VGND VPWR VPWR _9143_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4948_ _9544_/Q VGND VGND VPWR VPWR _4948_/Y sky130_fd_sc_hd__inv_4
X_7736_ _7736_/A VGND VGND VPWR VPWR _7736_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4879_ _9820_/Q VGND VGND VPWR VPWR _4879_/Y sky130_fd_sc_hd__inv_4
X_7667_ _6898_/Y _7509_/X _6903_/Y _7510_/X VGND VGND VPWR VPWR _7667_/X sky130_fd_sc_hd__o22a_1
X_9406_ _9695_/CLK _9406_/D _9689_/SET_B VGND VGND VPWR VPWR _9406_/Q sky130_fd_sc_hd__dfstp_1
X_6618_ _9430_/Q VGND VGND VPWR VPWR _6618_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7598_ _6329_/Y _7513_/X _6305_/Y _7514_/X _7597_/X VGND VGND VPWR VPWR _7603_/B
+ sky130_fd_sc_hd__o221a_1
X_9337_ _9421_/CLK _9337_/D _9537_/SET_B VGND VGND VPWR VPWR _9337_/Q sky130_fd_sc_hd__dfstp_1
X_6549_ _6547_/Y _5990_/B _6548_/Y _5112_/B VGND VGND VPWR VPWR _6549_/X sky130_fd_sc_hd__o22a_1
XFILLER_145_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9268_ _9431_/CLK _9268_/D _9817_/SET_B VGND VGND VPWR VPWR _9268_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput270 _9051_/Z VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_2
X_8219_ _8745_/A _8219_/B VGND VGND VPWR VPWR _8219_/X sky130_fd_sc_hd__or2_1
X_9199_ _9225_/CLK _9199_/D _9731_/SET_B VGND VGND VPWR VPWR _9199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput281 _9027_/Z VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_2
Xoutput292 _7048_/A VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_2
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5920_ _5889_/X _8924_/X _8960_/X _9185_/Q VGND VGND VPWR VPWR _9185_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5851_ _9238_/Q _5849_/A hold510/X _5849_/Y VGND VGND VPWR VPWR _5851_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4802_ _4802_/A VGND VGND VPWR VPWR _4802_/Y sky130_fd_sc_hd__clkinv_4
X_8570_ _8570_/A _8570_/B VGND VGND VPWR VPWR _8570_/Y sky130_fd_sc_hd__nor2_4
XFILLER_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5782_ _9098_/Q _5782_/B _5816_/A VGND VGND VPWR VPWR _5782_/X sky130_fd_sc_hd__and3_1
XFILLER_21_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4733_ _9254_/Q VGND VGND VPWR VPWR _4733_/Y sky130_fd_sc_hd__inv_2
X_7521_ _7521_/A VGND VGND VPWR VPWR _7521_/X sky130_fd_sc_hd__buf_6
XFILLER_119_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7452_ _7478_/C _7477_/A _7471_/C VGND VGND VPWR VPWR _7501_/A sky130_fd_sc_hd__or3_2
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6403_ _9264_/Q VGND VGND VPWR VPWR _6403_/Y sky130_fd_sc_hd__clkinv_2
X_4664_ _9758_/Q _4657_/A _8996_/X _4657_/Y VGND VGND VPWR VPWR _9758_/D sky130_fd_sc_hd__a22o_1
XFILLER_162_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4595_ _9790_/Q _4587_/A _6008_/B1 _4587_/Y VGND VGND VPWR VPWR _9790_/D sky130_fd_sc_hd__a22o_1
X_7383_ _6731_/Y _7180_/X _6732_/Y _7181_/X _7382_/X VGND VGND VPWR VPWR _7384_/D
+ sky130_fd_sc_hd__o221a_2
X_6334_ _9140_/Q VGND VGND VPWR VPWR _6334_/Y sky130_fd_sc_hd__clkinv_2
X_9122_ _9751_/CLK _9122_/D _6052_/X VGND VGND VPWR VPWR _9122_/Q sky130_fd_sc_hd__dfrtp_4
X_9053_ _9632_/Q _8841_/A VGND VGND VPWR VPWR _9053_/Z sky130_fd_sc_hd__ebufn_1
X_6265_ _6263_/Y _5068_/B _6264_/Y _4883_/X VGND VGND VPWR VPWR _6265_/X sky130_fd_sc_hd__o22a_1
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8004_ _8230_/A _8140_/B _8006_/B VGND VGND VPWR VPWR _8132_/B sky130_fd_sc_hd__a21bo_2
XFILLER_142_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5216_ _5216_/A VGND VGND VPWR VPWR _5216_/Y sky130_fd_sc_hd__inv_2
X_6196_ _6196_/A VGND VGND VPWR VPWR _8973_/S sky130_fd_sc_hd__inv_6
XFILLER_130_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5147_ _9673_/Q _5146_/A _8959_/A1 _5146_/Y VGND VGND VPWR VPWR _9673_/D sky130_fd_sc_hd__a22o_1
X_5078_ _9709_/Q _5070_/A _8975_/A1 _5070_/Y VGND VGND VPWR VPWR _9709_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8906_ _8905_/X hold706/X _9096_/Q VGND VGND VPWR VPWR _8906_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8837_ _8837_/A VGND VGND VPWR VPWR _8838_/A sky130_fd_sc_hd__clkbuf_1
X_8768_ _8118_/A _8288_/B _8285_/A _8356_/X _8546_/C VGND VGND VPWR VPWR _8769_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_44_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7719_ _6362_/Y _7500_/A _6443_/Y _7501_/A _7718_/X VGND VGND VPWR VPWR _7719_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8699_ _8699_/A _8699_/B _8699_/C _8699_/D VGND VGND VPWR VPWR _8738_/C sky130_fd_sc_hd__or4_4
XFILLER_193_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold208 _5855_/X VGND VGND VPWR VPWR hold209/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold219 hold219/A VGND VGND VPWR VPWR hold220/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6050_/A VGND VGND VPWR VPWR _9123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5001_/A VGND VGND VPWR VPWR _5001_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6952_ _9731_/Q VGND VGND VPWR VPWR _6952_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9740_ _9751_/CLK _9740_/D _5023_/X VGND VGND VPWR VPWR _9740_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5903_ _5903_/A VGND VGND VPWR VPWR _5904_/A sky130_fd_sc_hd__clkbuf_4
X_9671_ _9833_/CLK _9671_/D _9797_/SET_B VGND VGND VPWR VPWR _9671_/Q sky130_fd_sc_hd__dfrtp_2
X_6883_ _6874_/Y _5351_/B _6877_/X _6882_/X VGND VGND VPWR VPWR _6909_/C sky130_fd_sc_hd__o211a_1
X_5834_ _9248_/Q _5828_/A _8965_/A1 _5828_/Y VGND VGND VPWR VPWR _9248_/D sky130_fd_sc_hd__a22o_1
X_8622_ _8622_/A _8717_/C _8687_/D _8758_/A VGND VGND VPWR VPWR _8628_/A sky130_fd_sc_hd__or4_4
XFILLER_22_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8553_ _8324_/C _8608_/B _8629_/A _8715_/A VGND VGND VPWR VPWR _8554_/D sky130_fd_sc_hd__a211o_1
X_5765_ _5765_/A _9287_/Q VGND VGND VPWR VPWR _7128_/A sky130_fd_sc_hd__or2_2
X_8484_ _7935_/A _8540_/A _8065_/A _8053_/B VGND VGND VPWR VPWR _8486_/A sky130_fd_sc_hd__o22ai_2
X_5696_ _9312_/Q _5689_/A _6067_/B1 _5689_/Y VGND VGND VPWR VPWR _9312_/D sky130_fd_sc_hd__a22o_1
X_7504_ _6819_/Y _7502_/X _6885_/Y _7503_/X VGND VGND VPWR VPWR _7504_/X sky130_fd_sc_hd__o22a_1
X_4716_ _8847_/A VGND VGND VPWR VPWR _4716_/Y sky130_fd_sc_hd__inv_2
X_4647_ _6008_/B1 _9761_/Q _4647_/S VGND VGND VPWR VPWR _4648_/A sky130_fd_sc_hd__mux2_1
X_7435_ _7473_/A _7479_/C _9297_/Q VGND VGND VPWR VPWR _7486_/A sky130_fd_sc_hd__or3_4
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7366_ _6761_/Y _7135_/X _6736_/Y _7136_/X _7365_/X VGND VGND VPWR VPWR _7385_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9105_ _4471_/A1 _9105_/D _6177_/A VGND VGND VPWR VPWR _9105_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6317_ _6312_/Y _6196_/A _6313_/Y _5068_/B _6316_/X VGND VGND VPWR VPWR _6338_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4578_ _6142_/A _4827_/A VGND VGND VPWR VPWR _4579_/B sky130_fd_sc_hd__or2_4
X_7297_ _7297_/A _7297_/B _7297_/C VGND VGND VPWR VPWR _7297_/Y sky130_fd_sc_hd__nand3_4
XFILLER_115_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9036_ _9604_/Q _8807_/A VGND VGND VPWR VPWR _9036_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6248_ _6243_/Y _5902_/B _6244_/Y _6282_/A _6247_/X VGND VGND VPWR VPWR _6267_/A
+ sky130_fd_sc_hd__o221a_1
X_6179_ _6179_/A VGND VGND VPWR VPWR _6180_/A sky130_fd_sc_hd__buf_2
XFILLER_130_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold91 hold91/A VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5550_ _9401_/Q _5545_/A _6008_/B1 _5545_/Y VGND VGND VPWR VPWR _9401_/D sky130_fd_sc_hd__a22o_1
X_4501_ _6142_/A _4953_/A VGND VGND VPWR VPWR _4502_/B sky130_fd_sc_hd__or2_4
XFILLER_8_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5481_ _9448_/Q _5475_/X _6008_/B1 _5476_/Y VGND VGND VPWR VPWR _5481_/X sky130_fd_sc_hd__a22o_1
X_7220_ _8793_/A _7160_/X _6548_/Y _7071_/B _7219_/X VGND VGND VPWR VPWR _7221_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA_0 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7151_ _7151_/A VGND VGND VPWR VPWR _7151_/X sky130_fd_sc_hd__buf_6
X_6102_ _6102_/A _6102_/B VGND VGND VPWR VPWR _6102_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7082_ _7091_/C _7100_/B VGND VGND VPWR VPWR _7171_/A sky130_fd_sc_hd__or2_2
XFILLER_140_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6033_ _9129_/Q _6026_/A _8947_/X _6026_/Y VGND VGND VPWR VPWR _9129_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7984_ _8118_/A _8229_/B _9110_/Q VGND VGND VPWR VPWR _8556_/B sky130_fd_sc_hd__o21ai_1
XFILLER_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9723_ _9723_/CLK _9723_/D _6177_/A VGND VGND VPWR VPWR _9723_/Q sky130_fd_sc_hd__dfrtp_1
X_6935_ _9397_/Q VGND VGND VPWR VPWR _6935_/Y sky130_fd_sc_hd__inv_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9654_ _9731_/CLK _9654_/D _9731_/SET_B VGND VGND VPWR VPWR _9654_/Q sky130_fd_sc_hd__dfrtp_1
X_6866_ _6864_/Y _5123_/B _6865_/Y _4611_/B VGND VGND VPWR VPWR _6866_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8605_ _8605_/A _8755_/D _8755_/B _8678_/D VGND VGND VPWR VPWR _8605_/X sky130_fd_sc_hd__or4_1
X_9585_ _9600_/CLK _9585_/D _9821_/SET_B VGND VGND VPWR VPWR _9585_/Q sky130_fd_sc_hd__dfstp_1
X_6797_ _6797_/A VGND VGND VPWR VPWR _6797_/Y sky130_fd_sc_hd__clkinv_2
X_5817_ hold703/X _9098_/Q _5816_/Y _9259_/Q _5784_/A VGND VGND VPWR VPWR _9259_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8536_ _8557_/B _8229_/A _8702_/A _8538_/A _8383_/B VGND VGND VPWR VPWR _8636_/A
+ sky130_fd_sc_hd__a311oi_1
X_5748_ _9290_/Q VGND VGND VPWR VPWR _7068_/A sky130_fd_sc_hd__inv_2
X_8467_ _8730_/A _8673_/A _8467_/C VGND VGND VPWR VPWR _8469_/A sky130_fd_sc_hd__or3_1
XFILLER_108_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5679_ _5675_/B _5673_/X _5675_/A _5677_/X _5678_/Y VGND VGND VPWR VPWR _9322_/D
+ sky130_fd_sc_hd__o311a_1
X_8398_ _8398_/A _8398_/B _8613_/C _8719_/A VGND VGND VPWR VPWR _8402_/A sky130_fd_sc_hd__or4_1
X_7418_ _6400_/Y _7160_/A _6476_/Y _7064_/A _7417_/X VGND VGND VPWR VPWR _7419_/D
+ sky130_fd_sc_hd__o221a_1
Xhold572 _5171_/X VGND VGND VPWR VPWR _9659_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold561 _5525_/X VGND VGND VPWR VPWR _9420_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold550 _5343_/X VGND VGND VPWR VPWR _9543_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7349_ _6857_/Y _7095_/B _6959_/Y _7157_/X VGND VGND VPWR VPWR _7349_/X sky130_fd_sc_hd__o22a_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold594 hold594/A VGND VGND VPWR VPWR hold594/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold583 _5173_/X VGND VGND VPWR VPWR _9657_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9019_ _8971_/S _6353_/Y _9019_/S VGND VGND VPWR VPWR _9019_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput181 wb_dat_i[24] VGND VGND VPWR VPWR _7769_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput170 wb_dat_i[14] VGND VGND VPWR VPWR _7781_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput192 wb_dat_i[5] VGND VGND VPWR VPWR _9008_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4981_ _9133_/Q _6053_/C VGND VGND VPWR VPWR _4981_/Y sky130_fd_sc_hd__nor2_1
X_6720_ _6716_/Y _5047_/B _6717_/Y _5532_/B _6719_/X VGND VGND VPWR VPWR _6721_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6651_ _6646_/Y _5359_/B _8835_/A _5417_/B _6650_/X VGND VGND VPWR VPWR _6658_/C
+ sky130_fd_sc_hd__o221a_1
X_5602_ _9368_/Q _5600_/A hold510/X _5600_/Y VGND VGND VPWR VPWR _5602_/X sky130_fd_sc_hd__a22o_1
X_9370_ _9600_/CLK _9370_/D _9821_/SET_B VGND VGND VPWR VPWR _9370_/Q sky130_fd_sc_hd__dfrtp_1
X_6582_ _9686_/Q VGND VGND VPWR VPWR _6582_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5533_ _5533_/A VGND VGND VPWR VPWR _5534_/A sky130_fd_sc_hd__clkbuf_4
X_8321_ _8321_/A _8420_/B _8321_/C VGND VGND VPWR VPWR _8322_/C sky130_fd_sc_hd__or3_1
XFILLER_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5464_ _9459_/Q _5457_/A hold593/X _5457_/Y VGND VGND VPWR VPWR _9459_/D sky130_fd_sc_hd__a22o_1
X_8252_ _8252_/A VGND VGND VPWR VPWR _8302_/B sky130_fd_sc_hd__buf_4
XFILLER_172_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7203_ _6806_/Y _7171_/X _6755_/Y _7172_/X _7202_/X VGND VGND VPWR VPWR _7208_/B
+ sky130_fd_sc_hd__o221a_1
X_8183_ _8243_/B _8592_/A VGND VGND VPWR VPWR _8617_/A sky130_fd_sc_hd__nor2_1
X_5395_ _9506_/Q _5391_/A _6067_/B1 _5391_/Y VGND VGND VPWR VPWR _9506_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7134_ _7134_/A VGND VGND VPWR VPWR _7134_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7065_ _7128_/A _7118_/C VGND VGND VPWR VPWR _7121_/B sky130_fd_sc_hd__or2_1
XFILLER_59_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6016_ _9133_/Q _6015_/Y _6011_/X VGND VGND VPWR VPWR _9133_/D sky130_fd_sc_hd__o21ba_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7967_ _8367_/A _7967_/B VGND VGND VPWR VPWR _7968_/B sky130_fd_sc_hd__and2_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9706_ _4471_/A1 _9706_/D _6177_/A VGND VGND VPWR VPWR _9706_/Q sky130_fd_sc_hd__dfrtp_1
X_7898_ _8563_/B _8304_/B VGND VGND VPWR VPWR _8505_/A sky130_fd_sc_hd__nor2_1
X_6918_ _6916_/Y _5589_/B _6917_/Y _6083_/C VGND VGND VPWR VPWR _6918_/X sky130_fd_sc_hd__o22a_2
X_9637_ _9695_/CLK _9637_/D _9689_/SET_B VGND VGND VPWR VPWR _9637_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_13_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9522_/CLK sky130_fd_sc_hd__clkbuf_16
X_6849_ _9485_/Q VGND VGND VPWR VPWR _6849_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_168_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9568_ _9569_/CLK _9568_/D _9563_/SET_B VGND VGND VPWR VPWR _9568_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9499_ _9569_/CLK _9499_/D _9563_/SET_B VGND VGND VPWR VPWR _9499_/Q sky130_fd_sc_hd__dfrtp_1
X_8519_ _8519_/A _8763_/C VGND VGND VPWR VPWR _8520_/B sky130_fd_sc_hd__or2_1
XFILLER_6_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_28_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9491_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold380 _5244_/X VGND VGND VPWR VPWR hold381/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold391 hold391/A VGND VGND VPWR VPWR _5553_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5180_ _5180_/A VGND VGND VPWR VPWR _5181_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8870_ _9633_/Q input81/X _8875_/S VGND VGND VPWR VPWR _8870_/X sky130_fd_sc_hd__mux2_1
X_7821_ _8625_/A _7904_/D _7827_/B VGND VGND VPWR VPWR _7823_/B sky130_fd_sc_hd__or3_1
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4964_ _9132_/Q VGND VGND VPWR VPWR _6053_/C sky130_fd_sc_hd__clkinv_2
X_7752_ _9129_/Q _7751_/B _7753_/A VGND VGND VPWR VPWR _7752_/X sky130_fd_sc_hd__o21a_1
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6703_ _6698_/Y _5068_/B _6699_/Y _5513_/B _6702_/X VGND VGND VPWR VPWR _6721_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9422_ _9574_/CLK _9422_/D _9571_/SET_B VGND VGND VPWR VPWR _9422_/Q sky130_fd_sc_hd__dfrtp_1
X_7683_ _6774_/Y _7500_/X _6756_/Y _7501_/X _7682_/X VGND VGND VPWR VPWR _7683_/X
+ sky130_fd_sc_hd__o221a_1
X_4895_ _4887_/Y _5359_/B _4889_/Y _4890_/X _4894_/X VGND VGND VPWR VPWR _4918_/A
+ sky130_fd_sc_hd__o221a_1
X_6634_ _9521_/Q VGND VGND VPWR VPWR _8817_/A sky130_fd_sc_hd__inv_8
XFILLER_192_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9353_ _9678_/CLK _9353_/D _9730_/SET_B VGND VGND VPWR VPWR _9353_/Q sky130_fd_sc_hd__dfrtp_1
X_6565_ _9089_/Q VGND VGND VPWR VPWR _6565_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_180_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5516_ _9426_/Q _5515_/A _6064_/B1 _5515_/Y VGND VGND VPWR VPWR _9426_/D sky130_fd_sc_hd__a22o_1
X_6496_ _6494_/Y _5068_/B _6495_/Y _5103_/B VGND VGND VPWR VPWR _6496_/X sky130_fd_sc_hd__o22a_1
X_9284_ _9831_/CLK _9284_/D _9727_/SET_B VGND VGND VPWR VPWR _9284_/Q sky130_fd_sc_hd__dfstp_1
X_8304_ _8383_/A _8304_/B VGND VGND VPWR VPWR _8411_/B sky130_fd_sc_hd__nor2_1
X_8235_ _8246_/A VGND VGND VPWR VPWR _8388_/B sky130_fd_sc_hd__inv_2
X_5447_ _9473_/Q _5446_/A hold516/X _5446_/Y VGND VGND VPWR VPWR _5447_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5378_ _5378_/A _5378_/B VGND VGND VPWR VPWR _5379_/A sky130_fd_sc_hd__or2_1
X_8166_ _8255_/A _8443_/A VGND VGND VPWR VPWR _8613_/A sky130_fd_sc_hd__nor2_1
X_8097_ _8429_/A _8209_/A VGND VGND VPWR VPWR _8578_/A sky130_fd_sc_hd__or2_1
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7117_ _7127_/A _7117_/B VGND VGND VPWR VPWR _7166_/A sky130_fd_sc_hd__or2_2
XFILLER_86_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7048_ _7048_/A VGND VGND VPWR VPWR _7048_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8999_ _5030_/S _6053_/B _8999_/S VGND VGND VPWR VPWR _8999_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4680_ _7034_/C VGND VGND VPWR VPWR _8999_/S sky130_fd_sc_hd__clkinv_4
XFILLER_174_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6350_ _6345_/Y _5112_/B _6346_/Y _5979_/B _6349_/X VGND VGND VPWR VPWR _6356_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_161_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5301_ _5378_/A _5301_/B VGND VGND VPWR VPWR _5302_/A sky130_fd_sc_hd__or2_1
XFILLER_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6281_ _9679_/Q VGND VGND VPWR VPWR _6281_/Y sky130_fd_sc_hd__inv_2
X_8020_ _8570_/A _8034_/A VGND VGND VPWR VPWR _8032_/B sky130_fd_sc_hd__or2_4
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5232_ _9614_/Q _5226_/Y _8965_/X _5226_/A VGND VGND VPWR VPWR _5232_/X sky130_fd_sc_hd__o22a_1
XFILLER_124_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5163_ _9664_/Q _5159_/A _8959_/A1 _5159_/Y VGND VGND VPWR VPWR _9664_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5094_ _5094_/A VGND VGND VPWR VPWR _9705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8922_ _8921_/X _9183_/Q _9096_/Q VGND VGND VPWR VPWR _8922_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8853_ _8853_/A _8855_/B VGND VGND VPWR VPWR _9104_/D sky130_fd_sc_hd__nor2_1
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7804_ _8570_/A VGND VGND VPWR VPWR _8234_/A sky130_fd_sc_hd__inv_2
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8784_ _8771_/Y _8765_/Y _8773_/X _8783_/X VGND VGND VPWR VPWR _8784_/X sky130_fd_sc_hd__a31o_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5996_ _9144_/Q _5992_/A _8969_/A1 _5992_/Y VGND VGND VPWR VPWR _9144_/D sky130_fd_sc_hd__a22o_1
X_7735_ _7735_/A VGND VGND VPWR VPWR _7736_/A sky130_fd_sc_hd__clkbuf_1
X_4947_ _4947_/A _4953_/B VGND VGND VPWR VPWR _5389_/B sky130_fd_sc_hd__or2_4
XFILLER_149_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7666_ _6960_/Y _7497_/X _7663_/X _7665_/X VGND VGND VPWR VPWR _7676_/C sky130_fd_sc_hd__o211a_1
X_4878_ _4933_/A _4939_/A VGND VGND VPWR VPWR _5340_/B sky130_fd_sc_hd__or2_4
XFILLER_165_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6617_ _6617_/A _6617_/B _6617_/C VGND VGND VPWR VPWR _6659_/B sky130_fd_sc_hd__and3_1
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9405_ _9728_/CLK _9405_/D _9727_/SET_B VGND VGND VPWR VPWR _9405_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9336_ _9695_/CLK _9336_/D _9537_/SET_B VGND VGND VPWR VPWR _9336_/Q sky130_fd_sc_hd__dfstp_1
X_7597_ _6308_/Y _7515_/X _6345_/Y _7516_/X VGND VGND VPWR VPWR _7597_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6548_ _9691_/Q VGND VGND VPWR VPWR _6548_/Y sky130_fd_sc_hd__inv_2
X_9267_ _9736_/CLK _9267_/D _9731_/SET_B VGND VGND VPWR VPWR _9267_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6479_ _6465_/Y _4715_/X _6468_/X _6474_/X _6478_/X VGND VGND VPWR VPWR _6505_/C
+ sky130_fd_sc_hd__o2111a_1
Xoutput271 _9052_/Z VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_2
Xoutput260 _9042_/Z VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_2
X_8218_ _8762_/A _8602_/A _8218_/C VGND VGND VPWR VPWR _8219_/B sky130_fd_sc_hd__or3_1
X_9198_ _9225_/CLK _9198_/D _9731_/SET_B VGND VGND VPWR VPWR _9198_/Q sky130_fd_sc_hd__dfrtp_1
X_8149_ _8260_/A _8241_/B _8260_/C VGND VGND VPWR VPWR _8264_/C sky130_fd_sc_hd__or3_4
Xoutput282 _9028_/Z VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_1
XFILLER_99_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput293 _9771_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_2
XFILLER_181_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5850_ _9239_/Q _5849_/A hold516/X _5849_/Y VGND VGND VPWR VPWR _5850_/X sky130_fd_sc_hd__a22o_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4801_ _4933_/B _4801_/B VGND VGND VPWR VPWR _5786_/B sky130_fd_sc_hd__or2_4
XFILLER_21_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5781_ _9322_/Q _9321_/Q _9320_/Q VGND VGND VPWR VPWR _5816_/A sky130_fd_sc_hd__or3_1
X_4732_ _4953_/A _4732_/B VGND VGND VPWR VPWR _5658_/B sky130_fd_sc_hd__or2_4
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7520_ _7520_/A VGND VGND VPWR VPWR _7520_/X sky130_fd_sc_hd__buf_6
X_7451_ _7479_/A _9293_/Q _7476_/B _9297_/Q VGND VGND VPWR VPWR _7500_/A sky130_fd_sc_hd__or4_2
X_4663_ _4663_/A VGND VGND VPWR VPWR _4663_/X sky130_fd_sc_hd__clkbuf_1
X_6402_ _9302_/Q VGND VGND VPWR VPWR _6402_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4594_ _9791_/Q _4587_/A _6067_/B1 _4587_/Y VGND VGND VPWR VPWR _9791_/D sky130_fd_sc_hd__a22o_1
X_7382_ _6683_/Y _7182_/X _6793_/Y _7183_/X VGND VGND VPWR VPWR _7382_/X sky130_fd_sc_hd__o22a_1
X_6333_ _9198_/Q VGND VGND VPWR VPWR _6333_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9121_ _9832_/CLK _9121_/D _9821_/SET_B VGND VGND VPWR VPWR _9121_/Q sky130_fd_sc_hd__dfrtp_1
X_9052_ _9052_/A _8839_/A VGND VGND VPWR VPWR _9052_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6264_ _6264_/A VGND VGND VPWR VPWR _6264_/Y sky130_fd_sc_hd__clkinv_4
X_8003_ _8019_/A _8034_/B VGND VGND VPWR VPWR _8137_/B sky130_fd_sc_hd__or2_4
X_5215_ _6353_/A _6196_/A _5250_/A _8998_/X VGND VGND VPWR VPWR _5216_/A sky130_fd_sc_hd__a211o_4
XFILLER_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6195_ _9446_/Q VGND VGND VPWR VPWR _6195_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5146_ _5146_/A VGND VGND VPWR VPWR _5146_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5077_ _9710_/Q _5070_/A _8969_/A1 _5070_/Y VGND VGND VPWR VPWR _9710_/D sky130_fd_sc_hd__a22o_1
XFILLER_111_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8905_ _7658_/Y _9669_/Q _9020_/S VGND VGND VPWR VPWR _8905_/X sky130_fd_sc_hd__mux2_1
X_8836_ _8836_/A VGND VGND VPWR VPWR _8836_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5979_ _6083_/A _5979_/B VGND VGND VPWR VPWR _5980_/A sky130_fd_sc_hd__or2_1
X_8767_ _8744_/Y _8775_/A _8754_/Y _8781_/A _8766_/Y VGND VGND VPWR VPWR _8767_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7718_ _6361_/Y _7502_/A _6378_/Y _7503_/A VGND VGND VPWR VPWR _7718_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8698_ _7873_/B _7901_/Y _8560_/A _8409_/B VGND VGND VPWR VPWR _8699_/B sky130_fd_sc_hd__a31o_1
XFILLER_193_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7649_ _4870_/Y _7509_/X _4940_/Y _7510_/X VGND VGND VPWR VPWR _7649_/X sky130_fd_sc_hd__o22a_1
XFILLER_153_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9319_ _9319_/CLK _9319_/D _9797_/SET_B VGND VGND VPWR VPWR _9319_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold209 hold209/A VGND VGND VPWR VPWR hold210/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5000_ _5017_/A VGND VGND VPWR VPWR _5001_/A sky130_fd_sc_hd__clkbuf_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6951_ _9220_/Q VGND VGND VPWR VPWR _6951_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5902_ _6083_/A _5902_/B VGND VGND VPWR VPWR _5903_/A sky130_fd_sc_hd__or2_1
XFILLER_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9670_ _9833_/CLK _9670_/D _9797_/SET_B VGND VGND VPWR VPWR _9670_/Q sky130_fd_sc_hd__dfrtp_2
X_6882_ _6878_/Y _4890_/X _6879_/Y _5321_/B _6881_/X VGND VGND VPWR VPWR _6882_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_179_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5833_ _9249_/Q _5828_/A _8964_/A1 _5828_/Y VGND VGND VPWR VPWR _9249_/D sky130_fd_sc_hd__a22o_1
X_8621_ _8750_/B _8621_/B _8621_/C VGND VGND VPWR VPWR _8758_/A sky130_fd_sc_hd__or3_1
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8552_ _8552_/A _8702_/B _8702_/C VGND VGND VPWR VPWR _8645_/C sky130_fd_sc_hd__nor3_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5764_ _5723_/A _7113_/A _7081_/B _5719_/A _5763_/X VGND VGND VPWR VPWR _9289_/D
+ sky130_fd_sc_hd__o311a_1
X_7503_ _7503_/A VGND VGND VPWR VPWR _7503_/X sky130_fd_sc_hd__clkbuf_8
X_5695_ _9313_/Q _5689_/A hold217/X _5689_/Y VGND VGND VPWR VPWR _9313_/D sky130_fd_sc_hd__a22o_1
X_8483_ _8483_/A _8483_/B VGND VGND VPWR VPWR _8491_/A sky130_fd_sc_hd__nand2_1
X_4715_ _4818_/B _4865_/B VGND VGND VPWR VPWR _4715_/X sky130_fd_sc_hd__or2_4
XFILLER_135_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4646_ _4646_/A VGND VGND VPWR VPWR _9762_/D sky130_fd_sc_hd__clkbuf_1
X_7434_ _7441_/A _7436_/B VGND VGND VPWR VPWR _7479_/C sky130_fd_sc_hd__or2_2
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7365_ _6676_/Y _7137_/X _6787_/Y _7138_/X _7364_/X VGND VGND VPWR VPWR _7365_/X
+ sky130_fd_sc_hd__o221a_1
X_4577_ _4577_/A VGND VGND VPWR VPWR _9800_/D sky130_fd_sc_hd__clkbuf_1
Xhold710 hold710/A VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__clkbuf_2
X_9104_ _4471_/A1 _9104_/D _6177_/A VGND VGND VPWR VPWR _9104_/Q sky130_fd_sc_hd__dfrtp_1
X_6316_ _7270_/A _5636_/B _6315_/Y _5866_/B VGND VGND VPWR VPWR _6316_/X sky130_fd_sc_hd__o22a_1
XFILLER_115_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7296_ _7296_/A _7296_/B _7296_/C _7296_/D VGND VGND VPWR VPWR _7297_/C sky130_fd_sc_hd__and4_1
X_9035_ _9603_/Q _8805_/A VGND VGND VPWR VPWR _9035_/Z sky130_fd_sc_hd__ebufn_1
X_6247_ _6245_/Y _4598_/B _6246_/Y _5036_/B VGND VGND VPWR VPWR _6247_/X sky130_fd_sc_hd__o22a_1
XFILLER_39_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6178_ _7005_/B _6178_/B VGND VGND VPWR VPWR _6179_/A sky130_fd_sc_hd__or2_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5129_ _9684_/Q _5125_/A _6067_/B1 _5125_/Y VGND VGND VPWR VPWR _5129_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8819_ _8819_/A VGND VGND VPWR VPWR _8820_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9799_ _9800_/CLK _9799_/D _9821_/SET_B VGND VGND VPWR VPWR _9799_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_187_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold81 hold81/A VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4500_ _4750_/A _4750_/B _4689_/A _4642_/B VGND VGND VPWR VPWR _4953_/A sky130_fd_sc_hd__or4_4
X_5480_ _9449_/Q _5476_/A _6067_/B1 _5476_/Y VGND VGND VPWR VPWR _9449_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_1 _6613_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7150_ _7150_/A VGND VGND VPWR VPWR _7150_/X sky130_fd_sc_hd__buf_6
X_6101_ _6096_/Y _5866_/B _6097_/Y _5687_/B _6100_/X VGND VGND VPWR VPWR _6102_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7081_ _9290_/Q _7081_/B _9288_/Q _9287_/Q VGND VGND VPWR VPWR _7100_/B sky130_fd_sc_hd__or4_1
XFILLER_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6032_ _6032_/A VGND VGND VPWR VPWR _6032_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7983_ _7983_/A VGND VGND VPWR VPWR _7983_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6934_ _6934_/A VGND VGND VPWR VPWR _6934_/Y sky130_fd_sc_hd__clkinv_4
X_9722_ _9723_/CLK _9722_/D _6177_/A VGND VGND VPWR VPWR _9722_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9653_ _9731_/CLK _9653_/D _9731_/SET_B VGND VGND VPWR VPWR _9653_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8604_ _8604_/A _8714_/C _8715_/A VGND VGND VPWR VPWR _8678_/D sky130_fd_sc_hd__or3_1
X_6865_ _9775_/Q VGND VGND VPWR VPWR _6865_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6796_ _6791_/Y _5329_/B _6792_/Y _5263_/B _6795_/X VGND VGND VPWR VPWR _6814_/A
+ sky130_fd_sc_hd__o221a_1
X_9584_ _9600_/CLK _9584_/D _9821_/SET_B VGND VGND VPWR VPWR _9584_/Q sky130_fd_sc_hd__dfrtp_1
X_5816_ _5816_/A VGND VGND VPWR VPWR _5816_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8535_ _8656_/A _8535_/B _8535_/C VGND VGND VPWR VPWR _8699_/C sky130_fd_sc_hd__or3_1
X_5747_ _5765_/A _5766_/B VGND VGND VPWR VPWR _7113_/A sky130_fd_sc_hd__or2_2
XFILLER_41_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8466_ _8209_/A _8443_/B _8465_/X VGND VGND VPWR VPWR _8467_/C sky130_fd_sc_hd__o21bai_1
X_5678_ _5675_/B _5673_/X _5675_/A VGND VGND VPWR VPWR _5678_/Y sky130_fd_sc_hd__o21ai_1
X_7417_ _6404_/Y _7161_/A _6443_/Y _7162_/A VGND VGND VPWR VPWR _7417_/X sky130_fd_sc_hd__o22a_1
XFILLER_135_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8397_ _8725_/B _8541_/B VGND VGND VPWR VPWR _8719_/A sky130_fd_sc_hd__or2_1
X_4629_ _9770_/Q _4625_/A hold217/X _4625_/Y VGND VGND VPWR VPWR _9770_/D sky130_fd_sc_hd__a22o_1
Xhold562 _5193_/X VGND VGND VPWR VPWR _9643_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold551 _5562_/X VGND VGND VPWR VPWR _9395_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold540 _5613_/X VGND VGND VPWR VPWR _9360_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7348_ _6897_/Y _7149_/X _6966_/Y _7150_/X _7347_/X VGND VGND VPWR VPWR _7353_/B
+ sky130_fd_sc_hd__o221a_1
Xhold595 hold595/A VGND VGND VPWR VPWR hold595/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold573 _5640_/X VGND VGND VPWR VPWR _9342_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold584 _5639_/X VGND VGND VPWR VPWR _9343_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7279_ _6263_/Y _7071_/C _6255_/Y _7146_/X VGND VGND VPWR VPWR _7279_/X sky130_fd_sc_hd__o22a_1
XFILLER_103_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9018_ _8975_/S _6353_/Y _9019_/S VGND VGND VPWR VPWR _9018_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput171 wb_dat_i[15] VGND VGND VPWR VPWR _7783_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput160 wb_adr_i[6] VGND VGND VPWR VPWR _7942_/C sky130_fd_sc_hd__buf_4
Xinput182 wb_dat_i[25] VGND VGND VPWR VPWR _7771_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput193 wb_dat_i[6] VGND VGND VPWR VPWR _9009_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4980_ _4980_/A VGND VGND VPWR VPWR _4980_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6650_ _6648_/Y _5144_/B _6649_/Y _4892_/X VGND VGND VPWR VPWR _6650_/X sky130_fd_sc_hd__o22a_1
X_5601_ _9369_/Q _5600_/A hold516/X _5600_/Y VGND VGND VPWR VPWR _5601_/X sky130_fd_sc_hd__a22o_1
X_6581_ _9581_/Q VGND VGND VPWR VPWR _6581_/Y sky130_fd_sc_hd__clkinv_2
X_8320_ _8387_/A _8625_/C _8387_/B VGND VGND VPWR VPWR _8321_/A sky130_fd_sc_hd__or3b_1
X_5532_ _5570_/A _5532_/B VGND VGND VPWR VPWR _5533_/A sky130_fd_sc_hd__or2_1
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5463_ _9460_/Q _5456_/X hold136/X _5457_/Y VGND VGND VPWR VPWR _5463_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9516_/CLK sky130_fd_sc_hd__clkbuf_16
X_8251_ _8702_/A _8268_/C VGND VGND VPWR VPWR _8252_/A sky130_fd_sc_hd__or2_1
XFILLER_172_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7202_ _6725_/Y _7173_/X _6717_/Y _7174_/X VGND VGND VPWR VPWR _7202_/X sky130_fd_sc_hd__o22a_1
X_8182_ _8592_/A _8182_/B VGND VGND VPWR VPWR _8404_/A sky130_fd_sc_hd__nor2_1
X_5394_ _9507_/Q _5391_/A hold217/X _5391_/Y VGND VGND VPWR VPWR _9507_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7133_ _7133_/A _7133_/B _7133_/C VGND VGND VPWR VPWR _7134_/A sky130_fd_sc_hd__and3_1
XFILLER_101_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7064_ _7064_/A VGND VGND VPWR VPWR _7071_/B sky130_fd_sc_hd__buf_6
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6015_ _6053_/C _6015_/B VGND VGND VPWR VPWR _6015_/Y sky130_fd_sc_hd__nor2_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9705_ _9705_/CLK _9705_/D _6177_/A VGND VGND VPWR VPWR _9705_/Q sky130_fd_sc_hd__dfrtp_1
X_7966_ _8657_/A _7966_/B VGND VGND VPWR VPWR _7967_/B sky130_fd_sc_hd__nor2_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7897_ _7897_/A VGND VGND VPWR VPWR _8304_/B sky130_fd_sc_hd__clkbuf_2
X_6917_ _9087_/Q VGND VGND VPWR VPWR _6917_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9636_ _9643_/CLK _9636_/D _9689_/SET_B VGND VGND VPWR VPWR _9636_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6848_ _6848_/A VGND VGND VPWR VPWR _6848_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9567_ _9569_/CLK _9567_/D _9563_/SET_B VGND VGND VPWR VPWR _9567_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6779_ _9330_/Q VGND VGND VPWR VPWR _6779_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_168_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8518_ _8518_/A _8518_/B VGND VGND VPWR VPWR _8763_/C sky130_fd_sc_hd__or2_2
XFILLER_10_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9498_ _9569_/CLK _9498_/D _9563_/SET_B VGND VGND VPWR VPWR _9498_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8449_ _8449_/A VGND VGND VPWR VPWR _8649_/B sky130_fd_sc_hd__inv_2
Xhold381 hold381/A VGND VGND VPWR VPWR hold382/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold370 hold370/A VGND VGND VPWR VPWR hold371/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold392 _5551_/X VGND VGND VPWR VPWR _5552_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7820_ _8005_/A VGND VGND VPWR VPWR _8625_/A sky130_fd_sc_hd__buf_2
X_4963_ _9133_/Q VGND VGND VPWR VPWR _6053_/D sky130_fd_sc_hd__inv_2
X_7751_ _9129_/Q _7751_/B VGND VGND VPWR VPWR _7753_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7682_ _6810_/Y _7502_/X _6811_/Y _7503_/X VGND VGND VPWR VPWR _7682_/X sky130_fd_sc_hd__o22a_1
X_6702_ _6700_/Y _4854_/X _6701_/Y _4611_/B VGND VGND VPWR VPWR _6702_/X sky130_fd_sc_hd__o22a_2
X_9421_ _9421_/CLK _9421_/D _9537_/SET_B VGND VGND VPWR VPWR _9421_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4894_ _4891_/Y _4892_/X _4893_/Y _4579_/B VGND VGND VPWR VPWR _4894_/X sky130_fd_sc_hd__o22a_2
X_6633_ _6618_/Y _5505_/B _6621_/X _6627_/X _6632_/X VGND VGND VPWR VPWR _6659_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_192_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9352_ _9678_/CLK _9352_/D _9730_/SET_B VGND VGND VPWR VPWR _9352_/Q sky130_fd_sc_hd__dfrtp_1
X_6564_ _9699_/Q VGND VGND VPWR VPWR _6564_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_192_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5515_ _5515_/A VGND VGND VPWR VPWR _5515_/Y sky130_fd_sc_hd__inv_2
X_9283_ _9831_/CLK _9283_/D _9727_/SET_B VGND VGND VPWR VPWR _9283_/Q sky130_fd_sc_hd__dfrtp_1
X_8303_ _8303_/A _8620_/B VGND VGND VPWR VPWR _8305_/A sky130_fd_sc_hd__or2_1
X_6495_ _9700_/Q VGND VGND VPWR VPWR _6495_/Y sky130_fd_sc_hd__clkinv_2
X_8234_ _8234_/A _8234_/B _8236_/A VGND VGND VPWR VPWR _8246_/A sky130_fd_sc_hd__or3_4
XFILLER_172_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5446_ _5446_/A VGND VGND VPWR VPWR _5446_/Y sky130_fd_sc_hd__inv_2
X_5377_ _9518_/Q _5369_/A hold601/X _5369_/Y VGND VGND VPWR VPWR _5377_/X sky130_fd_sc_hd__a22o_1
XFILLER_160_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8165_ _8155_/Y _8156_/Y _8156_/Y _8432_/B _8164_/X VGND VGND VPWR VPWR _8168_/B
+ sky130_fd_sc_hd__a221o_1
X_8096_ _8096_/A _8750_/C VGND VGND VPWR VPWR _8098_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7116_ _7116_/A _7116_/B _7116_/C _7116_/D VGND VGND VPWR VPWR _7133_/B sky130_fd_sc_hd__and4_1
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7047_ _7047_/A VGND VGND VPWR VPWR _7048_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_47_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8998_ _8973_/S _6353_/Y _9019_/S VGND VGND VPWR VPWR _8998_/X sky130_fd_sc_hd__mux2_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7949_ _7957_/A _8281_/B VGND VGND VPWR VPWR _7949_/X sky130_fd_sc_hd__or2_2
XFILLER_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9619_ _9830_/CLK _9619_/D _9537_/SET_B VGND VGND VPWR VPWR _9619_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5300_ _9570_/Q _5291_/X hold601/A _5292_/Y VGND VGND VPWR VPWR _5300_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6280_ _6280_/A VGND VGND VPWR VPWR _6280_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_142_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5231_ _9615_/Q _5226_/Y _8964_/X _5226_/A VGND VGND VPWR VPWR _5231_/X sky130_fd_sc_hd__o22a_1
XFILLER_115_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5162_ _9665_/Q _5159_/A hold696/X _5159_/Y VGND VGND VPWR VPWR _9665_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5093_ _9007_/X _9705_/Q _5101_/S VGND VGND VPWR VPWR _5094_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_12_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9391_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8921_ _7253_/Y _9678_/Q _9001_/S VGND VGND VPWR VPWR _8921_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8852_ _8852_/A _8855_/B VGND VGND VPWR VPWR _9105_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_27_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9734_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7803_ _7803_/A _7803_/B _7803_/C _7803_/D VGND VGND VPWR VPWR _8006_/A sky130_fd_sc_hd__nand4_1
X_8783_ _8774_/Y _8775_/Y _8777_/X _8782_/X VGND VGND VPWR VPWR _8783_/X sky130_fd_sc_hd__a31o_1
XFILLER_37_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7734_ _7734_/A VGND VGND VPWR VPWR _7734_/X sky130_fd_sc_hd__clkbuf_1
X_5995_ _9145_/Q _5992_/A _8965_/A1 _5992_/Y VGND VGND VPWR VPWR _9145_/D sky130_fd_sc_hd__a22o_1
XFILLER_12_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4946_ _9505_/Q VGND VGND VPWR VPWR _4946_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4877_ _9536_/Q VGND VGND VPWR VPWR _4877_/Y sky130_fd_sc_hd__clkinv_4
X_7665_ _6953_/Y _7500_/X _6836_/Y _7501_/X _7664_/X VGND VGND VPWR VPWR _7665_/X
+ sky130_fd_sc_hd__o221a_1
X_7596_ _6339_/Y _7507_/X _6287_/Y _7508_/X _7595_/X VGND VGND VPWR VPWR _7603_/A
+ sky130_fd_sc_hd__o221a_1
X_6616_ _8787_/A _5036_/B _6612_/Y _5818_/B _6615_/X VGND VGND VPWR VPWR _6617_/C
+ sky130_fd_sc_hd__o221a_1
X_9404_ _9579_/CLK _9404_/D _9727_/SET_B VGND VGND VPWR VPWR _9404_/Q sky130_fd_sc_hd__dfrtp_1
X_9335_ _9569_/CLK _9335_/D _9563_/SET_B VGND VGND VPWR VPWR _9335_/Q sky130_fd_sc_hd__dfrtp_1
X_6547_ _9146_/Q VGND VGND VPWR VPWR _6547_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9266_ _9736_/CLK _9266_/D _9731_/SET_B VGND VGND VPWR VPWR _9266_/Q sky130_fd_sc_hd__dfrtp_1
X_6478_ _6475_/Y _4854_/X _6476_/Y _5123_/B _6477_/Y VGND VGND VPWR VPWR _6478_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput261 _9043_/Z VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput250 _9033_/Z VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_1
X_8217_ _8563_/A _8557_/A _8216_/Y VGND VGND VPWR VPWR _8218_/C sky130_fd_sc_hd__o21bai_1
X_9197_ _9416_/CLK _9197_/D _9731_/SET_B VGND VGND VPWR VPWR _9197_/Q sky130_fd_sc_hd__dfrtp_1
X_5429_ _5429_/A VGND VGND VPWR VPWR _5430_/A sky130_fd_sc_hd__clkbuf_2
Xoutput272 _9053_/Z VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_2
X_8148_ _8241_/C VGND VGND VPWR VPWR _8260_/C sky130_fd_sc_hd__inv_2
Xoutput294 _9772_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_2
Xoutput283 _8879_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8079_ _8563_/A _8594_/A VGND VGND VPWR VPWR _8458_/A sky130_fd_sc_hd__or2_1
XFILLER_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_151_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4800_ _9273_/Q VGND VGND VPWR VPWR _4800_/Y sky130_fd_sc_hd__inv_4
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _9322_/Q _9321_/Q _5780_/C _9319_/Q VGND VGND VPWR VPWR _5782_/B sky130_fd_sc_hd__or4_2
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _9323_/Q VGND VGND VPWR VPWR _7336_/A sky130_fd_sc_hd__clkinv_2
X_7450_ _4838_/Y _7498_/A _4763_/Y _5727_/A VGND VGND VPWR VPWR _7450_/X sky130_fd_sc_hd__o22a_1
X_4662_ _4969_/A VGND VGND VPWR VPWR _4663_/A sky130_fd_sc_hd__clkbuf_1
X_6401_ _6399_/Y _5786_/B _6400_/Y _5839_/B VGND VGND VPWR VPWR _6401_/X sky130_fd_sc_hd__o22a_1
X_7381_ _6743_/Y _5756_/A _6716_/Y _7061_/A _7380_/X VGND VGND VPWR VPWR _7384_/C
+ sky130_fd_sc_hd__o221a_1
X_9120_ _9832_/CLK _9120_/D _9821_/SET_B VGND VGND VPWR VPWR _9120_/Q sky130_fd_sc_hd__dfrtp_1
X_4593_ _9792_/Q _4587_/A hold217/A _4587_/Y VGND VGND VPWR VPWR _9792_/D sky130_fd_sc_hd__a22o_1
X_6332_ _9265_/Q VGND VGND VPWR VPWR _6332_/Y sky130_fd_sc_hd__inv_2
X_9051_ _9051_/A _8837_/A VGND VGND VPWR VPWR _9051_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6263_ _9715_/Q VGND VGND VPWR VPWR _6263_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_103_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8002_ _8570_/A _8000_/Y _8234_/A _8234_/B VGND VGND VPWR VPWR _8034_/B sky130_fd_sc_hd__o22a_1
XFILLER_115_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5214_ _9094_/Q _6015_/B _9628_/Q VGND VGND VPWR VPWR _9628_/D sky130_fd_sc_hd__a21o_1
X_6194_ _9360_/Q VGND VGND VPWR VPWR _6194_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_111_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5145_ _5145_/A VGND VGND VPWR VPWR _5146_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5076_ _9711_/Q _5070_/A _8965_/A1 _5070_/Y VGND VGND VPWR VPWR _9711_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8904_ _8903_/X _9212_/Q _9096_/Q VGND VGND VPWR VPWR _8904_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8835_ _8835_/A VGND VGND VPWR VPWR _8836_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_44_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8766_ _8771_/A _8773_/C _8765_/Y VGND VGND VPWR VPWR _8766_/Y sky130_fd_sc_hd__o21ai_1
X_5978_ _9156_/Q _5973_/A _8975_/A1 _5973_/Y VGND VGND VPWR VPWR _5978_/X sky130_fd_sc_hd__a22o_1
X_8697_ _8697_/A VGND VGND VPWR VPWR _8697_/Y sky130_fd_sc_hd__clkinv_2
X_7717_ _6422_/Y _7498_/A _6392_/Y _5727_/A VGND VGND VPWR VPWR _7717_/X sky130_fd_sc_hd__o22a_1
X_4929_ _6117_/A _6142_/B VGND VGND VPWR VPWR _4929_/X sky130_fd_sc_hd__or2_4
XFILLER_138_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7648_ _4786_/Y _7497_/X _7645_/X _7647_/X VGND VGND VPWR VPWR _7658_/C sky130_fd_sc_hd__o211a_1
XFILLER_193_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7579_ _6429_/Y _7515_/X _6470_/Y _7516_/X VGND VGND VPWR VPWR _7579_/X sky130_fd_sc_hd__o22a_1
X_9318_ _9318_/CLK _9318_/D _9537_/SET_B VGND VGND VPWR VPWR _9318_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9249_ _9420_/CLK _9249_/D _9537_/SET_B VGND VGND VPWR VPWR _9249_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6950_ _9149_/Q VGND VGND VPWR VPWR _6950_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5901_ _9201_/Q _5896_/A _6008_/B1 _5896_/Y VGND VGND VPWR VPWR _5901_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6881_ _9829_/Q _6282_/Y _6880_/Y _6117_/X VGND VGND VPWR VPWR _6881_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5832_ _9250_/Q _5828_/A hold53/X _5828_/Y VGND VGND VPWR VPWR _5832_/X sky130_fd_sc_hd__a22o_1
X_8620_ _8620_/A _8620_/B _8620_/C VGND VGND VPWR VPWR _8687_/D sky130_fd_sc_hd__or3_1
X_8551_ _8551_/A _8735_/A _8642_/B _8704_/B VGND VGND VPWR VPWR _8554_/B sky130_fd_sc_hd__or4_1
XFILLER_61_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5763_ _9288_/Q _9287_/Q _9097_/Q _9289_/Q VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__a31o_1
X_4714_ _9201_/Q VGND VGND VPWR VPWR _4714_/Y sky130_fd_sc_hd__clkinv_2
X_7502_ _7502_/A VGND VGND VPWR VPWR _7502_/X sky130_fd_sc_hd__clkbuf_8
X_5694_ _9314_/Q _5689_/A _8964_/A1 _5689_/Y VGND VGND VPWR VPWR _9314_/D sky130_fd_sc_hd__a22o_1
X_8482_ _7903_/X _8272_/A _8586_/A _8156_/Y VGND VGND VPWR VPWR _8707_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4645_ _6067_/B1 _9762_/Q _4645_/S VGND VGND VPWR VPWR _4646_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7433_ _9296_/Q VGND VGND VPWR VPWR _7441_/A sky130_fd_sc_hd__inv_2
Xhold700 _7017_/Y VGND VGND VPWR VPWR _9106_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7364_ _6754_/Y _7139_/X _6726_/Y _7140_/X VGND VGND VPWR VPWR _7364_/X sky130_fd_sc_hd__o22a_1
X_4576_ _6008_/B1 _9800_/Q _4576_/S VGND VGND VPWR VPWR _4577_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9103_ _4471_/A1 _9103_/D _6177_/A VGND VGND VPWR VPWR _9103_/Q sky130_fd_sc_hd__dfrtp_1
X_6315_ _9224_/Q VGND VGND VPWR VPWR _6315_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_1_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9034_ _9034_/A _8803_/A VGND VGND VPWR VPWR _9034_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_143_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7295_ _6195_/Y _7180_/X _6194_/Y _7181_/X _7294_/X VGND VGND VPWR VPWR _7296_/D
+ sky130_fd_sc_hd__o221a_1
X_6246_ _9736_/Q VGND VGND VPWR VPWR _6246_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_39_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6177_ _6177_/A VGND VGND VPWR VPWR _7005_/B sky130_fd_sc_hd__inv_2
XFILLER_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5128_ _9685_/Q hold685/X hold217/X _5125_/Y VGND VGND VPWR VPWR _9685_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5059_ _6011_/B VGND VGND VPWR VPWR _6015_/B sky130_fd_sc_hd__clkinv_2
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8818_ _8818_/A VGND VGND VPWR VPWR _8818_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9798_ _9798_/CLK _9798_/D _9821_/SET_B VGND VGND VPWR VPWR _9798_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_52_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8749_ _8749_/A _8749_/B _8749_/C VGND VGND VPWR VPWR _8775_/A sky130_fd_sc_hd__or3_2
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold82 hold82/A VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold60 hold60/A VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold93 hold93/A VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_90_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_2 _7550_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6100_ _6098_/Y _5647_/B _6099_/Y _5532_/B VGND VGND VPWR VPWR _6100_/X sky130_fd_sc_hd__o22a_1
XFILLER_125_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7080_ _7106_/B _7084_/C VGND VGND VPWR VPWR _7146_/A sky130_fd_sc_hd__or2_2
XFILLER_79_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6031_ _6071_/A VGND VGND VPWR VPWR _6032_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7982_ _8678_/A _7982_/B VGND VGND VPWR VPWR _7983_/A sky130_fd_sc_hd__or2_1
XFILLER_66_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9721_ _9723_/CLK _9721_/D _6177_/A VGND VGND VPWR VPWR _9721_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6933_ _9726_/Q VGND VGND VPWR VPWR _6933_/Y sky130_fd_sc_hd__inv_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9652_ _9731_/CLK _9652_/D _9731_/SET_B VGND VGND VPWR VPWR _9652_/Q sky130_fd_sc_hd__dfrtp_1
X_6864_ _9684_/Q VGND VGND VPWR VPWR _6864_/Y sky130_fd_sc_hd__inv_2
X_8603_ _8666_/B _8674_/B VGND VGND VPWR VPWR _8755_/B sky130_fd_sc_hd__nor2_1
X_5815_ _9260_/Q _5807_/A _8975_/A1 _5807_/Y VGND VGND VPWR VPWR _9260_/D sky130_fd_sc_hd__a22o_1
X_6795_ _6793_/Y _5274_/B _6794_/Y _5417_/B VGND VGND VPWR VPWR _6795_/X sky130_fd_sc_hd__o22a_1
X_9583_ _9600_/CLK _9583_/D _9821_/SET_B VGND VGND VPWR VPWR _9583_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8534_ _8534_/A VGND VGND VPWR VPWR _8656_/A sky130_fd_sc_hd__inv_2
X_5746_ _9287_/Q VGND VGND VPWR VPWR _5766_/B sky130_fd_sc_hd__inv_2
XFILLER_41_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8465_ _8750_/A _8750_/B _8464_/X VGND VGND VPWR VPWR _8465_/X sky130_fd_sc_hd__or3b_1
X_5677_ _5685_/A _5677_/B VGND VGND VPWR VPWR _5677_/X sky130_fd_sc_hd__or2_1
XFILLER_175_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4628_ _9771_/Q _4625_/A _6065_/B1 _4625_/Y VGND VGND VPWR VPWR _9771_/D sky130_fd_sc_hd__a22o_1
X_7416_ _6424_/Y _7155_/A _6454_/Y _7156_/A _7415_/X VGND VGND VPWR VPWR _7419_/C
+ sky130_fd_sc_hd__o221a_1
Xhold530 _5115_/X VGND VGND VPWR VPWR _9695_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_8396_ _8396_/A _8637_/B VGND VGND VPWR VPWR _8613_/C sky130_fd_sc_hd__or2_1
Xhold552 _5563_/X VGND VGND VPWR VPWR _9394_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold563 _8958_/X VGND VGND VPWR VPWR hold563/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_150_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold541 _6001_/X VGND VGND VPWR VPWR _9142_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4559_ _6008_/B1 _9803_/Q _4559_/S VGND VGND VPWR VPWR _4560_/A sky130_fd_sc_hd__mux2_1
X_7347_ _6874_/Y _7151_/X _6876_/Y _7152_/X VGND VGND VPWR VPWR _7347_/X sky130_fd_sc_hd__o22a_1
Xhold596 _5502_/X VGND VGND VPWR VPWR _9433_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold574 _5851_/X VGND VGND VPWR VPWR _9238_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold585 _5524_/X VGND VGND VPWR VPWR _9421_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7278_ _6191_/Y _7135_/X _6226_/Y _7136_/X _7277_/X VGND VGND VPWR VPWR _7297_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6229_ _6224_/Y _6353_/A _6225_/Y _5866_/B _6228_/X VGND VGND VPWR VPWR _6242_/B
+ sky130_fd_sc_hd__o221a_1
X_9017_ _8784_/X _8770_/X _9017_/S VGND VGND VPWR VPWR _9017_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput172 wb_dat_i[16] VGND VGND VPWR VPWR _7768_/B sky130_fd_sc_hd__clkbuf_1
Xinput150 wb_adr_i[26] VGND VGND VPWR VPWR input150/X sky130_fd_sc_hd__clkbuf_1
Xinput161 wb_adr_i[7] VGND VGND VPWR VPWR _8570_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput183 wb_dat_i[26] VGND VGND VPWR VPWR _7773_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput194 wb_dat_i[7] VGND VGND VPWR VPWR _9010_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5600_ _5600_/A VGND VGND VPWR VPWR _5600_/Y sky130_fd_sc_hd__inv_2
X_6580_ _9818_/Q VGND VGND VPWR VPWR _6580_/Y sky130_fd_sc_hd__inv_2
X_5531_ _9414_/Q _5523_/A _8975_/A1 _5523_/Y VGND VGND VPWR VPWR _9414_/D sky130_fd_sc_hd__a22o_1
X_8250_ _8347_/B _8306_/B VGND VGND VPWR VPWR _8637_/C sky130_fd_sc_hd__nor2_2
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5462_ _9461_/Q _5456_/X _8964_/A1 _5457_/Y VGND VGND VPWR VPWR _5462_/X sky130_fd_sc_hd__a22o_1
X_7201_ _6718_/Y _7071_/D _6768_/Y _7166_/X _7200_/X VGND VGND VPWR VPWR _7208_/A
+ sky130_fd_sc_hd__o221a_1
X_8181_ _8181_/A _8616_/A _8403_/A _8772_/A VGND VGND VPWR VPWR _8185_/A sky130_fd_sc_hd__or4_1
X_5393_ _9508_/Q _5391_/A _6065_/B1 _5391_/Y VGND VGND VPWR VPWR _9508_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7132_ _7132_/A _7132_/B _7132_/C _7132_/D VGND VGND VPWR VPWR _7133_/C sky130_fd_sc_hd__and4_1
XFILLER_113_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7063_ _7091_/C _7117_/B VGND VGND VPWR VPWR _7064_/A sky130_fd_sc_hd__or2_2
XFILLER_59_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6014_ _6014_/A VGND VGND VPWR VPWR _6014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9704_ _4471_/A1 _9704_/D _6177_/A VGND VGND VPWR VPWR _9704_/Q sky130_fd_sc_hd__dfrtp_1
X_7965_ _8229_/A _8312_/B _7964_/Y VGND VGND VPWR VPWR _7966_/B sky130_fd_sc_hd__o21ai_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7896_ _8489_/A _8302_/A VGND VGND VPWR VPWR _7897_/A sky130_fd_sc_hd__or2_1
X_6916_ _9371_/Q VGND VGND VPWR VPWR _6916_/Y sky130_fd_sc_hd__inv_2
X_9635_ _9643_/CLK _9635_/D _9563_/SET_B VGND VGND VPWR VPWR _9635_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6847_ _6842_/Y _4634_/B _6843_/Y _4525_/B _6846_/X VGND VGND VPWR VPWR _6860_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9566_ _9569_/CLK hold56/X _9563_/SET_B VGND VGND VPWR VPWR _9566_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6778_ _6773_/Y _5133_/B _6774_/Y _5946_/B _6777_/X VGND VGND VPWR VPWR _6790_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8517_ _8745_/C _8659_/A _8517_/C VGND VGND VPWR VPWR _8519_/A sky130_fd_sc_hd__or3_1
XFILLER_10_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5729_ _9295_/Q _7471_/A _5723_/A _9296_/Q VGND VGND VPWR VPWR _5729_/X sky130_fd_sc_hd__o31a_1
XFILLER_50_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9497_ _9569_/CLK _9497_/D _9563_/SET_B VGND VGND VPWR VPWR _9497_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8448_ _8171_/B _8443_/B _8444_/X _8447_/Y VGND VGND VPWR VPWR _8448_/X sky130_fd_sc_hd__o211a_1
X_8379_ _8678_/A _8692_/B _8379_/C VGND VGND VPWR VPWR _8380_/A sky130_fd_sc_hd__or3_1
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold371 hold371/A VGND VGND VPWR VPWR _4642_/B sky130_fd_sc_hd__buf_2
Xhold360 _6117_/A VGND VGND VPWR VPWR hold361/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold382 hold382/A VGND VGND VPWR VPWR _9608_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_117_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold393 _9720_/Q VGND VGND VPWR VPWR hold394/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4962_ _9134_/Q VGND VGND VPWR VPWR _6053_/A sky130_fd_sc_hd__inv_2
X_7750_ _7750_/A VGND VGND VPWR VPWR _7751_/B sky130_fd_sc_hd__inv_2
X_7681_ _6743_/Y _7498_/X _6663_/Y _5727_/A VGND VGND VPWR VPWR _7681_/X sky130_fd_sc_hd__o22a_1
X_6701_ _9776_/Q VGND VGND VPWR VPWR _6701_/Y sky130_fd_sc_hd__clkinv_2
X_4893_ _9798_/Q VGND VGND VPWR VPWR _4893_/Y sky130_fd_sc_hd__inv_2
X_9420_ _9420_/CLK _9420_/D _9537_/SET_B VGND VGND VPWR VPWR _9420_/Q sky130_fd_sc_hd__dfrtp_1
X_6632_ _6628_/Y _5255_/B _8827_/A _5263_/B _6631_/X VGND VGND VPWR VPWR _6632_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6563_ _9196_/Q VGND VGND VPWR VPWR _7731_/A sky130_fd_sc_hd__inv_4
X_9351_ _9678_/CLK _9351_/D _9730_/SET_B VGND VGND VPWR VPWR _9351_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5514_ _5514_/A VGND VGND VPWR VPWR _5514_/X sky130_fd_sc_hd__clkbuf_2
X_6494_ _9713_/Q VGND VGND VPWR VPWR _6494_/Y sky130_fd_sc_hd__inv_2
X_9282_ _9831_/CLK _9282_/D _9727_/SET_B VGND VGND VPWR VPWR _9282_/Q sky130_fd_sc_hd__dfrtp_1
X_8302_ _8302_/A _8302_/B VGND VGND VPWR VPWR _8620_/B sky130_fd_sc_hd__nor2_1
X_8233_ _8236_/A _8234_/B _8234_/A VGND VGND VPWR VPWR _8388_/A sky130_fd_sc_hd__o21a_1
X_5445_ _5445_/A VGND VGND VPWR VPWR _5445_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8164_ _8436_/C _7876_/A _8435_/A _8159_/X _8163_/X VGND VGND VPWR VPWR _8164_/X
+ sky130_fd_sc_hd__a41o_1
X_5376_ _9519_/Q _5369_/A hold593/X _5369_/Y VGND VGND VPWR VPWR _9519_/D sky130_fd_sc_hd__a22o_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7115_ _4755_/Y _7160_/A _4790_/Y _7064_/A _7114_/X VGND VGND VPWR VPWR _7116_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_160_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8095_ _8666_/B _8209_/A VGND VGND VPWR VPWR _8750_/C sky130_fd_sc_hd__nor2_2
XFILLER_101_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7046_ _9628_/Q _7046_/B VGND VGND VPWR VPWR _7047_/A sky130_fd_sc_hd__or2_1
XFILLER_103_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8997_ _9758_/Q _6268_/Y _8999_/S VGND VGND VPWR VPWR _8997_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7948_ _8042_/B _8281_/B _7916_/X _7946_/X _8345_/A VGND VGND VPWR VPWR _7948_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9618_ _9830_/CLK _9618_/D _9537_/SET_B VGND VGND VPWR VPWR _9618_/Q sky130_fd_sc_hd__dfrtp_1
X_7879_ _7957_/A VGND VGND VPWR VPWR _8557_/B sky130_fd_sc_hd__buf_6
XFILLER_23_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9549_ _9550_/CLK _9549_/D _9537_/SET_B VGND VGND VPWR VPWR _9549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold190 hold190/A VGND VGND VPWR VPWR hold191/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_8_csclk clkbuf_leaf_8_csclk/A VGND VGND VPWR VPWR _9514_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5230_ _9616_/Q _5226_/Y _8939_/X _5226_/A VGND VGND VPWR VPWR _5230_/X sky130_fd_sc_hd__o22a_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5161_ _9666_/Q _5159_/A hold510/X _5159_/Y VGND VGND VPWR VPWR _9666_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5092_ _5092_/A VGND VGND VPWR VPWR _9706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8920_ _8919_/X _9182_/Q _9096_/Q VGND VGND VPWR VPWR _8920_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8851_ _8851_/A VGND VGND VPWR VPWR _8851_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7802_ _8436_/A _8436_/B _7802_/C VGND VGND VPWR VPWR _7827_/B sky130_fd_sc_hd__or3_2
X_8782_ _8754_/B _8779_/Y _8731_/A _8780_/Y _8781_/Y VGND VGND VPWR VPWR _8782_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5994_ _9146_/Q _5992_/A _8964_/A1 _5992_/Y VGND VGND VPWR VPWR _9146_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7733_ _7733_/A VGND VGND VPWR VPWR _7734_/A sky130_fd_sc_hd__clkbuf_1
X_4945_ _4936_/Y _4937_/X _4938_/Y _5406_/B _4944_/X VGND VGND VPWR VPWR _4956_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4876_ _4868_/Y _4869_/X _4870_/Y _5466_/B _4875_/X VGND VGND VPWR VPWR _4886_/C
+ sky130_fd_sc_hd__o221a_1
X_7664_ _6905_/Y _7502_/X _6874_/Y _7503_/X VGND VGND VPWR VPWR _7664_/X sky130_fd_sc_hd__o22a_1
X_7595_ _6270_/Y _7509_/X _6300_/Y _7510_/X VGND VGND VPWR VPWR _7595_/X sky130_fd_sc_hd__o22a_1
X_6615_ _6613_/Y _5647_/B _6614_/Y _5551_/B VGND VGND VPWR VPWR _6615_/X sky130_fd_sc_hd__o22a_1
X_9403_ _9729_/CLK _9403_/D _9727_/SET_B VGND VGND VPWR VPWR _9403_/Q sky130_fd_sc_hd__dfstp_1
X_9334_ _9569_/CLK _9334_/D _9563_/SET_B VGND VGND VPWR VPWR _9334_/Q sky130_fd_sc_hd__dfrtp_1
X_6546_ _9314_/Q VGND VGND VPWR VPWR _8801_/A sky130_fd_sc_hd__inv_4
XFILLER_192_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6477_ input56/X _6353_/Y _8859_/A _4700_/Y VGND VGND VPWR VPWR _6477_/Y sky130_fd_sc_hd__a22oi_4
X_9265_ _9736_/CLK _9265_/D _9731_/SET_B VGND VGND VPWR VPWR _9265_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput262 _9044_/Z VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_2
Xoutput251 _9034_/Z VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__buf_2
X_8216_ _8216_/A _8216_/B VGND VGND VPWR VPWR _8216_/Y sky130_fd_sc_hd__nand2_1
X_9196_ _9491_/CLK _9196_/D _9731_/SET_B VGND VGND VPWR VPWR _9196_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput240 _8788_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_2
X_5428_ _5474_/A _5428_/B VGND VGND VPWR VPWR _5429_/A sky130_fd_sc_hd__or2_1
Xoutput273 _8870_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_2
X_8147_ _7789_/B _8145_/Y _7874_/B _8145_/A VGND VGND VPWR VPWR _8241_/C sky130_fd_sc_hd__o22a_1
XFILLER_87_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput295 _9773_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_2
Xoutput284 _7042_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_2
X_5359_ _5474_/A _5359_/B VGND VGND VPWR VPWR _5360_/A sky130_fd_sc_hd__or2_1
XFILLER_58_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8078_ _8586_/A _8027_/Y _8077_/Y VGND VGND VPWR VPWR _8080_/A sky130_fd_sc_hd__a21oi_1
XFILLER_101_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7029_ _5718_/A _7022_/Y _7027_/Y _7030_/A VGND VGND VPWR VPWR _9097_/D sky130_fd_sc_hd__o22ai_1
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4951_/A _4801_/B VGND VGND VPWR VPWR _5805_/B sky130_fd_sc_hd__or2_4
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4661_ _9759_/Q _4657_/A _8997_/X _4657_/Y VGND VGND VPWR VPWR _9759_/D sky130_fd_sc_hd__a22o_1
XFILLER_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7380_ _7380_/A _7380_/B VGND VGND VPWR VPWR _7380_/X sky130_fd_sc_hd__or2_1
X_6400_ _9244_/Q VGND VGND VPWR VPWR _6400_/Y sky130_fd_sc_hd__inv_2
X_6331_ _6327_/Y _5647_/B _6328_/Y _5036_/B _6330_/X VGND VGND VPWR VPWR _6338_/C
+ sky130_fd_sc_hd__o221a_1
X_4592_ _9793_/Q _4587_/A _6065_/B1 _4587_/Y VGND VGND VPWR VPWR _9793_/D sky130_fd_sc_hd__a22o_1
XFILLER_155_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9050_ _9643_/Q _8835_/A VGND VGND VPWR VPWR _9050_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_142_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6262_ _9680_/Q VGND VGND VPWR VPWR _6262_/Y sky130_fd_sc_hd__inv_2
X_8001_ _7999_/A _8236_/B _8000_/Y VGND VGND VPWR VPWR _8019_/A sky130_fd_sc_hd__a21oi_1
XFILLER_170_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6193_ _6188_/Y _5112_/B _6189_/X _6192_/X VGND VGND VPWR VPWR _6205_/B sky130_fd_sc_hd__o211a_1
X_5213_ _5213_/A VGND VGND VPWR VPWR _5213_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5144_ _5282_/A _5144_/B VGND VGND VPWR VPWR _5145_/A sky130_fd_sc_hd__or2_1
XFILLER_29_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5075_ _9712_/Q _5070_/A _8964_/A1 _5070_/Y VGND VGND VPWR VPWR _9712_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8903_ _7640_/Y _9681_/Q _9020_/S VGND VGND VPWR VPWR _8903_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8834_ _8834_/A VGND VGND VPWR VPWR _8834_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8765_ _8765_/A _8765_/B _8765_/C VGND VGND VPWR VPWR _8765_/Y sky130_fd_sc_hd__nor3_4
X_5977_ _9157_/Q _5973_/A _8969_/A1 _5973_/Y VGND VGND VPWR VPWR _9157_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8696_ _8747_/A _8749_/B _8662_/Y _8679_/X _8695_/X VGND VGND VPWR VPWR _8697_/A
+ sky130_fd_sc_hd__o311a_1
X_4928_ _4928_/A VGND VGND VPWR VPWR _4928_/Y sky130_fd_sc_hd__inv_2
X_7716_ _6404_/Y _7491_/A _6447_/Y _7492_/A _7715_/X VGND VGND VPWR VPWR _7730_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_138_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7647_ _4796_/Y _7500_/X _4858_/Y _7501_/X _7646_/X VGND VGND VPWR VPWR _7647_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4859_ _4941_/A _4933_/A VGND VGND VPWR VPWR _5255_/B sky130_fd_sc_hd__or2_4
X_7578_ _6399_/Y _7507_/X _6421_/Y _7508_/X _7577_/X VGND VGND VPWR VPWR _7585_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_180_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9317_ _9522_/CLK _9317_/D _9537_/SET_B VGND VGND VPWR VPWR _9317_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6529_ _9243_/Q VGND VGND VPWR VPWR _6529_/Y sky130_fd_sc_hd__inv_2
X_9248_ _9392_/CLK _9248_/D _9689_/SET_B VGND VGND VPWR VPWR _9248_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9179_ _9679_/CLK _9179_/D _9730_/SET_B VGND VGND VPWR VPWR _9179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_11_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9569_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9731_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5900_ _9202_/Q _5896_/A _6067_/B1 _5896_/Y VGND VGND VPWR VPWR _5900_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6880_ _6880_/A VGND VGND VPWR VPWR _6880_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5831_ _9251_/Q _5828_/A hold577/A _5828_/Y VGND VGND VPWR VPWR _5831_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8550_ _8324_/C _7868_/Y _8436_/A _7802_/C _8373_/B VGND VGND VPWR VPWR _8704_/B
+ sky130_fd_sc_hd__a41o_1
X_5762_ _7068_/A _5759_/Y _5723_/A _7107_/B VGND VGND VPWR VPWR _9290_/D sky130_fd_sc_hd__o22ai_1
X_4713_ _4705_/Y _5839_/B _4707_/Y _5979_/B _4712_/X VGND VGND VPWR VPWR _4725_/C
+ sky130_fd_sc_hd__o221a_1
X_7501_ _7501_/A VGND VGND VPWR VPWR _7501_/X sky130_fd_sc_hd__buf_4
XFILLER_147_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8481_ _8560_/A _8105_/B _8102_/C _8103_/B VGND VGND VPWR VPWR _8659_/A sky130_fd_sc_hd__a31o_1
X_5693_ _9315_/Q _5689_/A _6064_/B1 _5689_/Y VGND VGND VPWR VPWR _9315_/D sky130_fd_sc_hd__a22o_1
X_4644_ _5250_/A _4644_/B VGND VGND VPWR VPWR _4647_/S sky130_fd_sc_hd__or2_2
X_7432_ _9294_/Q _7432_/B VGND VGND VPWR VPWR _7473_/A sky130_fd_sc_hd__or2_2
Xhold701 _7018_/Y VGND VGND VPWR VPWR _9108_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_146_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7363_ _7363_/A _7363_/B _7363_/C VGND VGND VPWR VPWR _7363_/Y sky130_fd_sc_hd__nand3_2
X_4575_ _6189_/A _4947_/A _5282_/A VGND VGND VPWR VPWR _4576_/S sky130_fd_sc_hd__or3_1
X_6314_ _9341_/Q VGND VGND VPWR VPWR _7270_/A sky130_fd_sc_hd__clkinv_2
X_9102_ _4471_/A1 _9102_/D _6177_/A VGND VGND VPWR VPWR _9107_/D sky130_fd_sc_hd__dfrtp_1
X_7294_ _6219_/Y _7182_/X _6220_/Y _7183_/X VGND VGND VPWR VPWR _7294_/X sky130_fd_sc_hd__o22a_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9033_ _9033_/A _8801_/A VGND VGND VPWR VPWR _9033_/Z sky130_fd_sc_hd__ebufn_2
X_6245_ _9788_/Q VGND VGND VPWR VPWR _6245_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6176_ _6102_/Y _6176_/B _6176_/C _6176_/D VGND VGND VPWR VPWR _6176_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_97_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5127_ _9686_/Q hold685/X _6065_/B1 _5125_/Y VGND VGND VPWR VPWR _9686_/D sky130_fd_sc_hd__a22o_1
X_5058_ _9090_/Q _9092_/Q _9093_/Q VGND VGND VPWR VPWR _6011_/B sky130_fd_sc_hd__or3_2
XFILLER_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8817_ _8817_/A VGND VGND VPWR VPWR _8818_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9797_ _9798_/CLK _9797_/D _9797_/SET_B VGND VGND VPWR VPWR _9797_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_52_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8748_ _8748_/A _8748_/B _8748_/C _8748_/D VGND VGND VPWR VPWR _8749_/C sky130_fd_sc_hd__or4_1
XFILLER_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8679_ _8663_/Y _8675_/Y _8677_/Y _8756_/C VGND VGND VPWR VPWR _8679_/X sky130_fd_sc_hd__a31o_1
XFILLER_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 hold50/A VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold72 hold72/A VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold94 hold94/A VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR net399_3/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 _5201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6030_ _9130_/Q _6026_/A _8941_/X _6026_/Y VGND VGND VPWR VPWR _9130_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7981_ _8693_/A _8604_/A _7981_/C VGND VGND VPWR VPWR _7982_/B sky130_fd_sc_hd__or3_1
XFILLER_94_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9720_ _9723_/CLK _9720_/D _6177_/A VGND VGND VPWR VPWR _9720_/Q sky130_fd_sc_hd__dfrtp_1
X_6932_ _6932_/A _6932_/B _6932_/C _6932_/D VGND VGND VPWR VPWR _6976_/A sky130_fd_sc_hd__and4_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6863_ _9563_/Q VGND VGND VPWR VPWR _6863_/Y sky130_fd_sc_hd__clkinv_8
X_9651_ _9651_/CLK _9651_/D _9563_/SET_B VGND VGND VPWR VPWR _9651_/Q sky130_fd_sc_hd__dfrtp_1
X_8602_ _8602_/A _8602_/B VGND VGND VPWR VPWR _8755_/D sky130_fd_sc_hd__or2_2
X_5814_ _9261_/Q _5807_/A _8969_/A1 _5807_/Y VGND VGND VPWR VPWR _9261_/D sky130_fd_sc_hd__a22o_1
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6794_ _9486_/Q VGND VGND VPWR VPWR _6794_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9582_ _9582_/CLK _9582_/D _7042_/B VGND VGND VPWR VPWR _9582_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8533_ _7901_/Y _8344_/Y _8709_/A _8411_/B VGND VGND VPWR VPWR _8641_/D sky130_fd_sc_hd__a211o_1
X_5745_ _9288_/Q VGND VGND VPWR VPWR _5765_/A sky130_fd_sc_hd__inv_2
X_8464_ _8596_/A _8443_/B _8461_/X _8463_/Y VGND VGND VPWR VPWR _8464_/X sky130_fd_sc_hd__o211a_1
X_5676_ _9096_/Q _7028_/C _9098_/Q VGND VGND VPWR VPWR _5677_/B sky130_fd_sc_hd__a21o_1
XFILLER_148_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7415_ _6448_/Y _7056_/A _6410_/Y _7157_/A VGND VGND VPWR VPWR _7415_/X sky130_fd_sc_hd__o22a_1
X_4627_ _9772_/Q _4625_/A _6064_/B1 _4625_/Y VGND VGND VPWR VPWR _9772_/D sky130_fd_sc_hd__a22o_1
Xhold520 _5409_/X VGND VGND VPWR VPWR _9499_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_8395_ _8205_/A _8158_/A _8385_/Y _8265_/X _8394_/X VGND VGND VPWR VPWR _8398_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_135_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold553 _5116_/X VGND VGND VPWR VPWR _9694_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold531 _5829_/X VGND VGND VPWR VPWR _9253_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold542 _5710_/X VGND VGND VPWR VPWR _9304_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_150_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7346_ _6914_/Y _7144_/X _6831_/Y _7145_/X _7345_/X VGND VGND VPWR VPWR _7353_/A
+ sky130_fd_sc_hd__o221a_1
X_4558_ _5250_/A _4558_/B VGND VGND VPWR VPWR _4559_/S sky130_fd_sc_hd__or2_2
Xhold575 _9706_/Q VGND VGND VPWR VPWR hold576/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _5242_/X VGND VGND VPWR VPWR _9610_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_173_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold597 _5071_/X VGND VGND VPWR VPWR _9716_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_7277_ _6209_/Y _7137_/X _6182_/Y _7138_/X _7276_/X VGND VGND VPWR VPWR _7277_/X
+ sky130_fd_sc_hd__o221a_1
Xhold586 _5160_/X VGND VGND VPWR VPWR _9667_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_4489_ _4823_/A _4685_/B _4823_/C VGND VGND VPWR VPWR _4803_/A sky130_fd_sc_hd__or3_4
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6228_ _6226_/Y _5378_/B _6227_/Y _5367_/B VGND VGND VPWR VPWR _6228_/X sky130_fd_sc_hd__o22a_1
X_9016_ _8767_/Y _8739_/X _9017_/S VGND VGND VPWR VPWR _9016_/X sky130_fd_sc_hd__mux2_1
X_6159_ _9200_/Q VGND VGND VPWR VPWR _6159_/Y sky130_fd_sc_hd__inv_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater392 _8959_/A1 VGND VGND VPWR VPWR _6064_/B1 sky130_fd_sc_hd__buf_12
XFILLER_60_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput151 wb_adr_i[27] VGND VGND VPWR VPWR _5960_/A sky130_fd_sc_hd__clkbuf_1
Xinput140 wb_adr_i[17] VGND VGND VPWR VPWR _7803_/A sky130_fd_sc_hd__clkbuf_1
Xinput162 wb_adr_i[8] VGND VGND VPWR VPWR _7809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput184 wb_dat_i[27] VGND VGND VPWR VPWR _7775_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput173 wb_dat_i[17] VGND VGND VPWR VPWR _7770_/B sky130_fd_sc_hd__clkbuf_1
Xinput195 wb_dat_i[8] VGND VGND VPWR VPWR _7769_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5530_ _9415_/Q _5523_/A _8969_/A1 _5523_/Y VGND VGND VPWR VPWR _9415_/D sky130_fd_sc_hd__a22o_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5461_ _9462_/Q _5456_/X hold53/X _5457_/Y VGND VGND VPWR VPWR _5461_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7200_ _6692_/Y _7167_/X _6786_/Y _7168_/X VGND VGND VPWR VPWR _7200_/X sky130_fd_sc_hd__o22a_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8180_ _8180_/A _8682_/B VGND VGND VPWR VPWR _8772_/A sky130_fd_sc_hd__nor2_1
X_5392_ _9509_/Q _5391_/A _6064_/B1 _5391_/Y VGND VGND VPWR VPWR _9509_/D sky130_fd_sc_hd__a22o_1
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7131_ _4950_/Y _7180_/A _4792_/Y _7181_/A _7130_/X VGND VGND VPWR VPWR _7132_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7062_ _7129_/A _7118_/C VGND VGND VPWR VPWR _7117_/B sky130_fd_sc_hd__or2_1
XFILLER_113_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6013_ _6017_/A VGND VGND VPWR VPWR _6014_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7964_ _8641_/A _7964_/B VGND VGND VPWR VPWR _7964_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9703_ _4471_/A1 _9703_/D _6177_/A VGND VGND VPWR VPWR _9703_/Q sky130_fd_sc_hd__dfrtp_1
X_6915_ _9355_/Q VGND VGND VPWR VPWR _6915_/Y sky130_fd_sc_hd__inv_2
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7895_ _8567_/A _7933_/B _7999_/A _8570_/A VGND VGND VPWR VPWR _8302_/A sky130_fd_sc_hd__or4_4
XFILLER_82_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9634_ _9643_/CLK _9634_/D _9563_/SET_B VGND VGND VPWR VPWR _9634_/Q sky130_fd_sc_hd__dfrtp_1
X_6846_ _6844_/Y _4892_/X _6845_/Y _4644_/B VGND VGND VPWR VPWR _6846_/X sky130_fd_sc_hd__o22a_1
XFILLER_50_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9565_ _9569_/CLK hold65/X _9563_/SET_B VGND VGND VPWR VPWR _9565_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6777_ _6775_/Y _4863_/X _6776_/Y _5123_/B VGND VGND VPWR VPWR _6777_/X sky130_fd_sc_hd__o22a_2
X_8516_ _8516_/A _8516_/B VGND VGND VPWR VPWR _8517_/C sky130_fd_sc_hd__or2_1
X_5728_ _9297_/Q _5719_/Y _5723_/Y _5723_/A _5727_/X VGND VGND VPWR VPWR _9297_/D
+ sky130_fd_sc_hd__o32a_1
X_9496_ _9569_/CLK hold62/X _9563_/SET_B VGND VGND VPWR VPWR _9496_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8447_ _8447_/A VGND VGND VPWR VPWR _8447_/Y sky130_fd_sc_hd__inv_2
X_5659_ _5659_/A VGND VGND VPWR VPWR _5659_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8378_ _8715_/A _8378_/B VGND VGND VPWR VPWR _8379_/C sky130_fd_sc_hd__or2_1
XFILLER_136_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold350 hold350/A VGND VGND VPWR VPWR hold350/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_89_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold361 hold361/A VGND VGND VPWR VPWR hold362/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7329_ _4733_/Y _7161_/X _4858_/Y _7162_/X VGND VGND VPWR VPWR _7329_/X sky130_fd_sc_hd__o22a_1
Xhold372 _5195_/X VGND VGND VPWR VPWR hold373/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold383 _9721_/Q VGND VGND VPWR VPWR hold384/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 hold394/A VGND VGND VPWR VPWR hold395/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4961_ _4961_/A VGND VGND VPWR VPWR _4961_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4892_ _6117_/A _4922_/B VGND VGND VPWR VPWR _4892_/X sky130_fd_sc_hd__or2_4
X_7680_ _6671_/Y _7491_/X _6803_/Y _7492_/X _7679_/X VGND VGND VPWR VPWR _7694_/B
+ sky130_fd_sc_hd__o221a_1
X_6700_ _6700_/A VGND VGND VPWR VPWR _6700_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6631_ _9111_/Q _6282_/Y _6630_/Y _4623_/B VGND VGND VPWR VPWR _6631_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9350_ _9678_/CLK _9350_/D _9730_/SET_B VGND VGND VPWR VPWR _9350_/Q sky130_fd_sc_hd__dfrtp_1
X_6562_ _6562_/A VGND VGND VPWR VPWR _6562_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8301_ _8301_/A _8409_/B VGND VGND VPWR VPWR _8303_/A sky130_fd_sc_hd__or2_1
XFILLER_145_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6493_ _9734_/Q VGND VGND VPWR VPWR _6493_/Y sky130_fd_sc_hd__inv_2
X_5513_ _5698_/A _5513_/B VGND VGND VPWR VPWR _5513_/X sky130_fd_sc_hd__or2_1
X_9281_ _9322_/CLK _9281_/D _9797_/SET_B VGND VGND VPWR VPWR _9281_/Q sky130_fd_sc_hd__dfrtp_1
X_8232_ _8387_/A VGND VGND VPWR VPWR _8625_/B sky130_fd_sc_hd__inv_2
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5444_ _5570_/A _5444_/B VGND VGND VPWR VPWR _5444_/X sky130_fd_sc_hd__or2_1
XFILLER_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8163_ _7925_/B _8608_/A _8588_/A _8162_/Y VGND VGND VPWR VPWR _8163_/X sky130_fd_sc_hd__o31a_1
X_5375_ _9520_/Q _5369_/A hold136/X _5369_/Y VGND VGND VPWR VPWR _5375_/X sky130_fd_sc_hd__a22o_1
X_7114_ _4728_/Y _7161_/A _4814_/Y _7162_/A VGND VGND VPWR VPWR _7114_/X sky130_fd_sc_hd__o22a_1
X_8094_ _8094_/A _8434_/A VGND VGND VPWR VPWR _8096_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7045_ _7045_/A VGND VGND VPWR VPWR _7045_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8996_ _9757_/Q _6357_/Y _8999_/S VGND VGND VPWR VPWR _8996_/X sky130_fd_sc_hd__mux2_1
X_7947_ _7953_/A _8274_/B VGND VGND VPWR VPWR _8345_/A sky130_fd_sc_hd__or2_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _8421_/D _8436_/B _8436_/C _8236_/A VGND VGND VPWR VPWR _7957_/A sky130_fd_sc_hd__or4_4
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9617_ _9736_/CLK _9617_/D _9731_/SET_B VGND VGND VPWR VPWR _9617_/Q sky130_fd_sc_hd__dfrtp_1
X_6829_ _6824_/Y _5559_/B _6825_/Y _4929_/X _6828_/X VGND VGND VPWR VPWR _6861_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9548_ _9576_/CLK _9548_/D _9537_/SET_B VGND VGND VPWR VPWR _9548_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9479_ _9483_/CLK _9479_/D _9727_/SET_B VGND VGND VPWR VPWR _9479_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold180 hold180/A VGND VGND VPWR VPWR hold181/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xhold191 hold191/A VGND VGND VPWR VPWR hold191/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5160_ _9667_/Q _5159_/A hold516/X _5159_/Y VGND VGND VPWR VPWR _5160_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5091_ _9008_/X _9706_/Q _5101_/S VGND VGND VPWR VPWR _5092_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8850_ _8850_/A _8850_/B VGND VGND VPWR VPWR _8850_/Y sky130_fd_sc_hd__nor2_2
X_7801_ _7875_/B VGND VGND VPWR VPWR _7802_/C sky130_fd_sc_hd__inv_2
X_8781_ _8781_/A VGND VGND VPWR VPWR _8781_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5993_ _9147_/Q _5992_/A _8959_/A1 _5992_/Y VGND VGND VPWR VPWR _9147_/D sky130_fd_sc_hd__a22o_1
X_7732_ _7732_/A VGND VGND VPWR VPWR _7732_/X sky130_fd_sc_hd__clkbuf_1
X_4944_ _4940_/Y _5505_/B _4942_/Y _5543_/B VGND VGND VPWR VPWR _4944_/X sky130_fd_sc_hd__o22a_1
X_7663_ _6887_/Y _7498_/X _6969_/Y _5727_/X VGND VGND VPWR VPWR _7663_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4875_ _4872_/Y _5378_/B _4874_/Y _4545_/B VGND VGND VPWR VPWR _4875_/X sky130_fd_sc_hd__o22a_1
X_9402_ _9728_/CLK _9402_/D _9727_/SET_B VGND VGND VPWR VPWR _9402_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7594_ _6346_/Y _7497_/X _7591_/X _7593_/X VGND VGND VPWR VPWR _7604_/C sky130_fd_sc_hd__o211a_1
X_6614_ _9399_/Q VGND VGND VPWR VPWR _6614_/Y sky130_fd_sc_hd__inv_2
X_9333_ _9569_/CLK _9333_/D _9563_/SET_B VGND VGND VPWR VPWR _9333_/Q sky130_fd_sc_hd__dfrtp_1
X_6545_ _9235_/Q VGND VGND VPWR VPWR _8791_/A sky130_fd_sc_hd__inv_4
XFILLER_137_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9264_ _9734_/CLK _9264_/D _9731_/SET_B VGND VGND VPWR VPWR _9264_/Q sky130_fd_sc_hd__dfrtp_1
X_8215_ _8418_/A _8215_/B VGND VGND VPWR VPWR _8216_/B sky130_fd_sc_hd__nor2_1
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6476_ _9687_/Q VGND VGND VPWR VPWR _6476_/Y sky130_fd_sc_hd__clkinv_4
Xoutput230 _8834_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_2
Xoutput252 _9035_/Z VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_2
X_9195_ _9491_/CLK _9195_/D _9731_/SET_B VGND VGND VPWR VPWR _9195_/Q sky130_fd_sc_hd__dfrtp_1
X_5427_ _9484_/Q _5419_/A _8975_/A1 _5419_/Y VGND VGND VPWR VPWR _9484_/D sky130_fd_sc_hd__a22o_1
Xoutput241 _7734_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_2
Xoutput263 _9045_/Z VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_2
Xoutput274 _8871_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_2
X_8146_ _7869_/A _8145_/A _8009_/A _8145_/Y VGND VGND VPWR VPWR _8241_/B sky130_fd_sc_hd__a22o_1
Xoutput285 _8878_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_2
X_5358_ _9531_/Q _5353_/A _6008_/B1 _5353_/Y VGND VGND VPWR VPWR _9531_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8077_ _8429_/A _8593_/A _8076_/X VGND VGND VPWR VPWR _8077_/Y sky130_fd_sc_hd__o21ai_1
Xoutput296 _9800_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_2
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7028_ _7028_/A _8861_/X _7028_/C VGND VGND VPWR VPWR _7030_/A sky130_fd_sc_hd__or3_1
X_5289_ _9578_/Q _5284_/A _6008_/B1 _5284_/Y VGND VGND VPWR VPWR _5289_/X sky130_fd_sc_hd__a22o_1
XFILLER_87_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8979_ hold404/X hold395/X _9629_/Q VGND VGND VPWR VPWR _8979_/X sky130_fd_sc_hd__mux2_4
XFILLER_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4660_ _4660_/A VGND VGND VPWR VPWR _4660_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6330_ input49/X _8975_/S _6329_/Y _5847_/B VGND VGND VPWR VPWR _6330_/X sky130_fd_sc_hd__o2bb2a_1
X_4591_ _9794_/Q _4587_/A _6064_/B1 _4587_/Y VGND VGND VPWR VPWR _9794_/D sky130_fd_sc_hd__a22o_1
XFILLER_155_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6261_ _9141_/Q VGND VGND VPWR VPWR _6261_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8000_ _8234_/B VGND VGND VPWR VPWR _8000_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_142_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6192_ _6190_/Y _5406_/B _6191_/Y _5340_/B VGND VGND VPWR VPWR _6192_/X sky130_fd_sc_hd__o22a_1
XFILLER_130_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5212_ _6017_/A VGND VGND VPWR VPWR _5213_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_69_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5143_ _9674_/Q _5135_/A _8975_/A1 _5135_/Y VGND VGND VPWR VPWR _9674_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5074_ _9713_/Q _5070_/A _8959_/A1 _5070_/Y VGND VGND VPWR VPWR _9713_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8902_ _8901_/X _9211_/Q _9096_/Q VGND VGND VPWR VPWR _8902_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8833_ _8833_/A VGND VGND VPWR VPWR _8834_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_92_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8764_ _8764_/A _8764_/B _8764_/C VGND VGND VPWR VPWR _8765_/B sky130_fd_sc_hd__or3_1
X_5976_ _9158_/Q _5973_/A _8965_/A1 _5973_/Y VGND VGND VPWR VPWR _9158_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8695_ _8680_/Y _8689_/Y _8691_/Y _8694_/X VGND VGND VPWR VPWR _8695_/X sky130_fd_sc_hd__a31o_1
X_4927_ _4919_/Y _5367_/B _4921_/Y _5428_/B _4926_/X VGND VGND VPWR VPWR _4956_/A
+ sky130_fd_sc_hd__o221a_1
X_7715_ _6495_/Y _7493_/A _6372_/Y _7494_/A VGND VGND VPWR VPWR _7715_/X sky130_fd_sc_hd__o22a_1
X_4858_ _9596_/Q VGND VGND VPWR VPWR _4858_/Y sky130_fd_sc_hd__clkinv_2
X_7646_ _4822_/Y _7502_/X _4952_/Y _7503_/X VGND VGND VPWR VPWR _7646_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9316_ _9318_/CLK _9316_/D _9571_/SET_B VGND VGND VPWR VPWR _9316_/Q sky130_fd_sc_hd__dfrtp_1
X_7577_ _6388_/Y _7509_/X _6359_/Y _7510_/X VGND VGND VPWR VPWR _7577_/X sky130_fd_sc_hd__o22a_1
X_4789_ _7125_/A _5636_/B _4782_/Y _5858_/B _4788_/X VGND VGND VPWR VPWR _4811_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6528_ _9285_/Q VGND VGND VPWR VPWR _6528_/Y sky130_fd_sc_hd__inv_2
X_6459_ _9462_/Q VGND VGND VPWR VPWR _6459_/Y sky130_fd_sc_hd__inv_2
X_9247_ _9392_/CLK _9247_/D _9537_/SET_B VGND VGND VPWR VPWR _9247_/Q sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_7_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9577_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9178_ _9679_/CLK _9178_/D _9730_/SET_B VGND VGND VPWR VPWR _9178_/Q sky130_fd_sc_hd__dfrtp_1
X_8129_ _8229_/B _8429_/A VGND VGND VPWR VPWR _8475_/B sky130_fd_sc_hd__nor2_1
XFILLER_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5830_ _9252_/Q _5828_/A hold510/X _5828_/Y VGND VGND VPWR VPWR _5830_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5761_ _9290_/Q _7081_/B _7113_/A VGND VGND VPWR VPWR _7107_/B sky130_fd_sc_hd__or3_1
X_8480_ _8557_/A _8563_/B VGND VGND VPWR VPWR _8745_/D sky130_fd_sc_hd__nor2_1
X_4712_ _4712_/A _5047_/B VGND VGND VPWR VPWR _4712_/X sky130_fd_sc_hd__or2_1
X_7500_ _7500_/A VGND VGND VPWR VPWR _7500_/X sky130_fd_sc_hd__buf_4
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5692_ _9316_/Q _5689_/A hold577/A _5689_/Y VGND VGND VPWR VPWR _5692_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7431_ _7479_/A _9293_/Q _7467_/A _7471_/C VGND VGND VPWR VPWR _7485_/A sky130_fd_sc_hd__or4_4
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4643_ _4643_/A _4915_/B VGND VGND VPWR VPWR _4644_/B sky130_fd_sc_hd__or2_4
Xhold702 _7019_/Y VGND VGND VPWR VPWR _9109_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_4574_ _4689_/A _4642_/B _4689_/C _4750_/B VGND VGND VPWR VPWR _4947_/A sky130_fd_sc_hd__or4_4
X_7362_ _7362_/A _7362_/B _7362_/C _7362_/D VGND VGND VPWR VPWR _7363_/C sky130_fd_sc_hd__and4_1
X_9101_ _4471_/A1 _9101_/D _6177_/A VGND VGND VPWR VPWR _9101_/Q sky130_fd_sc_hd__dfstp_1
X_6313_ _9714_/Q VGND VGND VPWR VPWR _6313_/Y sky130_fd_sc_hd__inv_2
X_7293_ _6231_/Y _5756_/X _6261_/Y _7071_/A _7292_/X VGND VGND VPWR VPWR _7296_/C
+ sky130_fd_sc_hd__o221a_1
X_9032_ _9032_/A _8799_/A VGND VGND VPWR VPWR _9032_/Z sky130_fd_sc_hd__ebufn_1
XFILLER_115_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6244_ _8865_/X VGND VGND VPWR VPWR _6244_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6175_ _6175_/A _6175_/B _6175_/C _6175_/D VGND VGND VPWR VPWR _6176_/D sky130_fd_sc_hd__and4_2
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5126_ _9687_/Q hold685/X _6064_/B1 _5125_/Y VGND VGND VPWR VPWR _9687_/D sky130_fd_sc_hd__a22o_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5057_ _9094_/Q VGND VGND VPWR VPWR _5057_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8816_ _8816_/A VGND VGND VPWR VPWR _8816_/X sky130_fd_sc_hd__clkbuf_1
X_9796_ _9798_/CLK _9796_/D _9797_/SET_B VGND VGND VPWR VPWR _9796_/Q sky130_fd_sc_hd__dfstp_1
X_5959_ _7816_/A _7816_/B VGND VGND VPWR VPWR _7874_/C sky130_fd_sc_hd__or2_1
X_8747_ _8747_/A _8747_/B _8747_/C _8747_/D VGND VGND VPWR VPWR _8748_/D sky130_fd_sc_hd__or4_1
XFILLER_52_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8678_ _8678_/A _8678_/B _8678_/C _8678_/D VGND VGND VPWR VPWR _8756_/C sky130_fd_sc_hd__or4_2
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7629_ _6154_/Y _7500_/X _6114_/Y _7501_/X _7628_/X VGND VGND VPWR VPWR _7629_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold40 hold40/A VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold73 hold73/A VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold84 hold84/A VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_4 _6083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7980_ _8629_/A _7980_/B VGND VGND VPWR VPWR _7981_/C sky130_fd_sc_hd__or2_1
X_6931_ _6926_/Y _5598_/B _6927_/Y _5927_/B _6930_/X VGND VGND VPWR VPWR _6932_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9650_ _9651_/CLK _9650_/D _9563_/SET_B VGND VGND VPWR VPWR _9650_/Q sky130_fd_sc_hd__dfrtp_1
X_6862_ _6862_/A VGND VGND VPWR VPWR _6862_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8601_ _8601_/A _8751_/A _8673_/B _8730_/B VGND VGND VPWR VPWR _8605_/A sky130_fd_sc_hd__or4_1
X_5813_ _9262_/Q _5807_/A _8965_/A1 _5807_/Y VGND VGND VPWR VPWR _9262_/D sky130_fd_sc_hd__a22o_1
XFILLER_62_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9581_ _9686_/CLK _9581_/D _7042_/B VGND VGND VPWR VPWR _9581_/Q sky130_fd_sc_hd__dfrtp_1
X_8532_ _8776_/A _8532_/B _8532_/C VGND VGND VPWR VPWR _8639_/D sky130_fd_sc_hd__or3_1
X_6793_ _9585_/Q VGND VGND VPWR VPWR _6793_/Y sky130_fd_sc_hd__clkinv_4
X_5744_ _9291_/Q VGND VGND VPWR VPWR _5753_/B sky130_fd_sc_hd__inv_2
XFILLER_157_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8463_ _8672_/C VGND VGND VPWR VPWR _8463_/Y sky130_fd_sc_hd__inv_2
X_5675_ _5675_/A _5675_/B _9320_/Q _9319_/Q VGND VGND VPWR VPWR _7028_/C sky130_fd_sc_hd__or4_2
XFILLER_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8394_ _8394_/A _8394_/B _8394_/C VGND VGND VPWR VPWR _8394_/X sky130_fd_sc_hd__and3_1
XFILLER_135_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4626_ _9773_/Q _4625_/A hold696/X _4625_/Y VGND VGND VPWR VPWR _9773_/D sky130_fd_sc_hd__a22o_1
X_7414_ _6430_/Y _7149_/A _6405_/Y _7150_/A _7413_/X VGND VGND VPWR VPWR _7419_/B
+ sky130_fd_sc_hd__o221a_1
Xhold510 hold510/A VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__buf_12
XFILLER_135_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7345_ _6971_/Y _7071_/C _6953_/Y _7146_/X VGND VGND VPWR VPWR _7345_/X sky130_fd_sc_hd__o22a_1
Xhold521 _5410_/X VGND VGND VPWR VPWR _9498_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold532 _5536_/X VGND VGND VPWR VPWR _9412_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold554 _5344_/X VGND VGND VPWR VPWR _9542_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold543 _5448_/X VGND VGND VPWR VPWR _9472_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_131_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4557_ _6142_/A _4951_/A VGND VGND VPWR VPWR _4558_/B sky130_fd_sc_hd__or2_4
Xhold565 _5194_/X VGND VGND VPWR VPWR _9642_/D sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold576 hold576/A VGND VGND VPWR VPWR hold576/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_143_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7276_ _6190_/Y _7139_/X _6256_/Y _7140_/X VGND VGND VPWR VPWR _7276_/X sky130_fd_sc_hd__o22a_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4488_ _4476_/Y _8985_/X hold470/X VGND VGND VPWR VPWR _4488_/X sky130_fd_sc_hd__a21bo_1
Xhold587 _4548_/X VGND VGND VPWR VPWR _9811_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6227_ _9524_/Q VGND VGND VPWR VPWR _6227_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9015_ _8734_/Y _8706_/X _9017_/S VGND VGND VPWR VPWR _9015_/X sky130_fd_sc_hd__mux2_1
Xhold598 _5485_/X VGND VGND VPWR VPWR _9447_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_6158_ _9155_/Q VGND VGND VPWR VPWR _6158_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9550_/CLK sky130_fd_sc_hd__clkbuf_16
X_5109_ _9697_/Q _5105_/A _8969_/A1 _5105_/Y VGND VGND VPWR VPWR _9697_/D sky130_fd_sc_hd__a22o_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _9086_/Q _6085_/A _8975_/A1 _6085_/Y VGND VGND VPWR VPWR _9086_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater393 hold53/X VGND VGND VPWR VPWR _8959_/A1 sky130_fd_sc_hd__buf_12
XFILLER_45_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_25_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9736_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9779_ _9819_/CLK _9779_/D _9821_/SET_B VGND VGND VPWR VPWR _9779_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_opt_2_1_wb_clk_i clkbuf_opt_2_1_wb_clk_i/A VGND VGND VPWR VPWR _9062_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput130 usr2_vcc_pwrgood VGND VGND VPWR VPWR _6707_/A sky130_fd_sc_hd__clkbuf_1
Xinput152 wb_adr_i[28] VGND VGND VPWR VPWR _5960_/B sky130_fd_sc_hd__clkbuf_1
Xinput141 wb_adr_i[18] VGND VGND VPWR VPWR _7803_/D sky130_fd_sc_hd__clkbuf_1
Xinput163 wb_adr_i[9] VGND VGND VPWR VPWR _7809_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_48_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput185 wb_dat_i[28] VGND VGND VPWR VPWR _7777_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput174 wb_dat_i[18] VGND VGND VPWR VPWR _7772_/B sky130_fd_sc_hd__clkbuf_1
Xinput196 wb_dat_i[9] VGND VGND VPWR VPWR _7771_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5460_ _9463_/Q _5456_/X hold577/A _5457_/Y VGND VGND VPWR VPWR _5460_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5391_ _5391_/A VGND VGND VPWR VPWR _5391_/Y sky130_fd_sc_hd__inv_2
X_7130_ _4836_/Y _7182_/A _4879_/Y _7183_/A VGND VGND VPWR VPWR _7130_/X sky130_fd_sc_hd__o22a_1
XFILLER_113_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7061_ _7061_/A VGND VGND VPWR VPWR _7071_/A sky130_fd_sc_hd__buf_4
XFILLER_140_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6012_ _9134_/Q _6011_/X _7039_/A _6015_/B VGND VGND VPWR VPWR _9134_/D sky130_fd_sc_hd__o22a_1
.ends

