magic
tech sky130A
magscale 1 2
timestamp 1681048878
<< obsli1 >>
rect 1104 2159 80868 107729
<< obsm1 >>
rect 1026 1504 81958 107840
<< metal2 >>
rect 5906 109390 5962 110190
rect 6458 109390 6514 110190
rect 7010 109390 7066 110190
rect 7562 109390 7618 110190
rect 8114 109390 8170 110190
rect 8666 109390 8722 110190
rect 9218 109390 9274 110190
rect 9770 109390 9826 110190
rect 10322 109390 10378 110190
rect 10874 109390 10930 110190
rect 11426 109390 11482 110190
rect 11978 109390 12034 110190
rect 12530 109390 12586 110190
rect 13082 109390 13138 110190
rect 13634 109390 13690 110190
rect 14186 109390 14242 110190
rect 14738 109390 14794 110190
rect 15290 109390 15346 110190
rect 15842 109390 15898 110190
rect 16394 109390 16450 110190
rect 16946 109390 17002 110190
rect 17498 109390 17554 110190
rect 18050 109390 18106 110190
rect 18602 109390 18658 110190
rect 19154 109390 19210 110190
rect 19706 109390 19762 110190
rect 20258 109390 20314 110190
rect 20810 109390 20866 110190
rect 21362 109390 21418 110190
rect 21914 109390 21970 110190
rect 22466 109390 22522 110190
rect 23018 109390 23074 110190
rect 23570 109390 23626 110190
rect 24122 109390 24178 110190
rect 24674 109390 24730 110190
rect 25226 109390 25282 110190
rect 25778 109390 25834 110190
rect 26330 109390 26386 110190
rect 26882 109390 26938 110190
rect 27434 109390 27490 110190
rect 27986 109390 28042 110190
rect 28538 109390 28594 110190
rect 29090 109390 29146 110190
rect 29642 109390 29698 110190
rect 30194 109390 30250 110190
rect 30746 109390 30802 110190
rect 31298 109390 31354 110190
rect 31850 109390 31906 110190
rect 32402 109390 32458 110190
rect 32954 109390 33010 110190
rect 33506 109390 33562 110190
rect 34058 109390 34114 110190
rect 34610 109390 34666 110190
rect 35162 109390 35218 110190
rect 35714 109390 35770 110190
rect 36266 109390 36322 110190
rect 36818 109390 36874 110190
rect 37370 109390 37426 110190
rect 37922 109390 37978 110190
rect 38474 109390 38530 110190
rect 39026 109390 39082 110190
rect 39578 109390 39634 110190
rect 40130 109390 40186 110190
rect 40682 109390 40738 110190
rect 41234 109390 41290 110190
rect 41786 109390 41842 110190
rect 42338 109390 42394 110190
rect 42890 109390 42946 110190
rect 43442 109390 43498 110190
rect 43994 109390 44050 110190
rect 44546 109390 44602 110190
rect 45098 109390 45154 110190
rect 45650 109390 45706 110190
rect 46202 109390 46258 110190
rect 46754 109390 46810 110190
rect 47306 109390 47362 110190
rect 47858 109390 47914 110190
rect 48410 109390 48466 110190
rect 48962 109390 49018 110190
rect 49514 109390 49570 110190
rect 50066 109390 50122 110190
rect 50618 109390 50674 110190
rect 51170 109390 51226 110190
rect 51722 109390 51778 110190
rect 52274 109390 52330 110190
rect 52826 109390 52882 110190
rect 53378 109390 53434 110190
rect 53930 109390 53986 110190
rect 54482 109390 54538 110190
rect 55034 109390 55090 110190
rect 55586 109390 55642 110190
rect 56138 109390 56194 110190
rect 56690 109390 56746 110190
rect 57242 109390 57298 110190
rect 57794 109390 57850 110190
rect 58346 109390 58402 110190
rect 58898 109390 58954 110190
rect 59450 109390 59506 110190
rect 60002 109390 60058 110190
rect 60554 109390 60610 110190
rect 61106 109390 61162 110190
rect 61658 109390 61714 110190
rect 62210 109390 62266 110190
rect 62762 109390 62818 110190
rect 63314 109390 63370 110190
rect 63866 109390 63922 110190
rect 64418 109390 64474 110190
rect 64970 109390 65026 110190
rect 65522 109390 65578 110190
rect 66074 109390 66130 110190
rect 66626 109390 66682 110190
rect 67178 109390 67234 110190
rect 67730 109390 67786 110190
rect 68282 109390 68338 110190
rect 68834 109390 68890 110190
rect 69386 109390 69442 110190
rect 69938 109390 69994 110190
rect 70490 109390 70546 110190
rect 71042 109390 71098 110190
rect 71594 109390 71650 110190
rect 72146 109390 72202 110190
rect 72698 109390 72754 110190
rect 73250 109390 73306 110190
rect 73802 109390 73858 110190
rect 74354 109390 74410 110190
rect 74906 109390 74962 110190
rect 75458 109390 75514 110190
rect 76010 109390 76066 110190
rect 2870 0 2926 800
rect 3698 0 3754 800
rect 4526 0 4582 800
rect 5354 0 5410 800
rect 6182 0 6238 800
rect 7010 0 7066 800
rect 7838 0 7894 800
rect 8666 0 8722 800
rect 9494 0 9550 800
rect 10322 0 10378 800
rect 11150 0 11206 800
rect 11978 0 12034 800
rect 12806 0 12862 800
rect 13634 0 13690 800
rect 14462 0 14518 800
rect 15290 0 15346 800
rect 16118 0 16174 800
rect 16946 0 17002 800
rect 17774 0 17830 800
rect 18602 0 18658 800
rect 19430 0 19486 800
rect 20258 0 20314 800
rect 21086 0 21142 800
rect 21914 0 21970 800
rect 22742 0 22798 800
rect 23570 0 23626 800
rect 24398 0 24454 800
rect 25226 0 25282 800
rect 26054 0 26110 800
rect 26882 0 26938 800
rect 27710 0 27766 800
rect 28538 0 28594 800
rect 29366 0 29422 800
rect 30194 0 30250 800
rect 31022 0 31078 800
rect 31850 0 31906 800
rect 32678 0 32734 800
rect 33506 0 33562 800
rect 34334 0 34390 800
rect 35162 0 35218 800
rect 35990 0 36046 800
rect 36818 0 36874 800
rect 37646 0 37702 800
rect 38474 0 38530 800
rect 39302 0 39358 800
rect 40130 0 40186 800
rect 40958 0 41014 800
rect 41786 0 41842 800
rect 42614 0 42670 800
rect 43442 0 43498 800
rect 44270 0 44326 800
rect 45098 0 45154 800
rect 45926 0 45982 800
rect 46754 0 46810 800
rect 47582 0 47638 800
rect 48410 0 48466 800
rect 49238 0 49294 800
rect 50066 0 50122 800
rect 50894 0 50950 800
rect 51722 0 51778 800
rect 52550 0 52606 800
rect 53378 0 53434 800
rect 54206 0 54262 800
rect 55034 0 55090 800
rect 55862 0 55918 800
rect 56690 0 56746 800
rect 57518 0 57574 800
rect 58346 0 58402 800
rect 59174 0 59230 800
rect 60002 0 60058 800
rect 60830 0 60886 800
rect 61658 0 61714 800
rect 62486 0 62542 800
rect 63314 0 63370 800
rect 64142 0 64198 800
rect 64970 0 65026 800
rect 65798 0 65854 800
rect 66626 0 66682 800
rect 67454 0 67510 800
rect 68282 0 68338 800
rect 69110 0 69166 800
rect 69938 0 69994 800
rect 70766 0 70822 800
rect 71594 0 71650 800
rect 72422 0 72478 800
rect 73250 0 73306 800
rect 74078 0 74134 800
rect 74906 0 74962 800
rect 75734 0 75790 800
rect 76562 0 76618 800
rect 77390 0 77446 800
rect 78218 0 78274 800
rect 79046 0 79102 800
<< obsm2 >>
rect 1030 109334 5850 109426
rect 6018 109334 6402 109426
rect 6570 109334 6954 109426
rect 7122 109334 7506 109426
rect 7674 109334 8058 109426
rect 8226 109334 8610 109426
rect 8778 109334 9162 109426
rect 9330 109334 9714 109426
rect 9882 109334 10266 109426
rect 10434 109334 10818 109426
rect 10986 109334 11370 109426
rect 11538 109334 11922 109426
rect 12090 109334 12474 109426
rect 12642 109334 13026 109426
rect 13194 109334 13578 109426
rect 13746 109334 14130 109426
rect 14298 109334 14682 109426
rect 14850 109334 15234 109426
rect 15402 109334 15786 109426
rect 15954 109334 16338 109426
rect 16506 109334 16890 109426
rect 17058 109334 17442 109426
rect 17610 109334 17994 109426
rect 18162 109334 18546 109426
rect 18714 109334 19098 109426
rect 19266 109334 19650 109426
rect 19818 109334 20202 109426
rect 20370 109334 20754 109426
rect 20922 109334 21306 109426
rect 21474 109334 21858 109426
rect 22026 109334 22410 109426
rect 22578 109334 22962 109426
rect 23130 109334 23514 109426
rect 23682 109334 24066 109426
rect 24234 109334 24618 109426
rect 24786 109334 25170 109426
rect 25338 109334 25722 109426
rect 25890 109334 26274 109426
rect 26442 109334 26826 109426
rect 26994 109334 27378 109426
rect 27546 109334 27930 109426
rect 28098 109334 28482 109426
rect 28650 109334 29034 109426
rect 29202 109334 29586 109426
rect 29754 109334 30138 109426
rect 30306 109334 30690 109426
rect 30858 109334 31242 109426
rect 31410 109334 31794 109426
rect 31962 109334 32346 109426
rect 32514 109334 32898 109426
rect 33066 109334 33450 109426
rect 33618 109334 34002 109426
rect 34170 109334 34554 109426
rect 34722 109334 35106 109426
rect 35274 109334 35658 109426
rect 35826 109334 36210 109426
rect 36378 109334 36762 109426
rect 36930 109334 37314 109426
rect 37482 109334 37866 109426
rect 38034 109334 38418 109426
rect 38586 109334 38970 109426
rect 39138 109334 39522 109426
rect 39690 109334 40074 109426
rect 40242 109334 40626 109426
rect 40794 109334 41178 109426
rect 41346 109334 41730 109426
rect 41898 109334 42282 109426
rect 42450 109334 42834 109426
rect 43002 109334 43386 109426
rect 43554 109334 43938 109426
rect 44106 109334 44490 109426
rect 44658 109334 45042 109426
rect 45210 109334 45594 109426
rect 45762 109334 46146 109426
rect 46314 109334 46698 109426
rect 46866 109334 47250 109426
rect 47418 109334 47802 109426
rect 47970 109334 48354 109426
rect 48522 109334 48906 109426
rect 49074 109334 49458 109426
rect 49626 109334 50010 109426
rect 50178 109334 50562 109426
rect 50730 109334 51114 109426
rect 51282 109334 51666 109426
rect 51834 109334 52218 109426
rect 52386 109334 52770 109426
rect 52938 109334 53322 109426
rect 53490 109334 53874 109426
rect 54042 109334 54426 109426
rect 54594 109334 54978 109426
rect 55146 109334 55530 109426
rect 55698 109334 56082 109426
rect 56250 109334 56634 109426
rect 56802 109334 57186 109426
rect 57354 109334 57738 109426
rect 57906 109334 58290 109426
rect 58458 109334 58842 109426
rect 59010 109334 59394 109426
rect 59562 109334 59946 109426
rect 60114 109334 60498 109426
rect 60666 109334 61050 109426
rect 61218 109334 61602 109426
rect 61770 109334 62154 109426
rect 62322 109334 62706 109426
rect 62874 109334 63258 109426
rect 63426 109334 63810 109426
rect 63978 109334 64362 109426
rect 64530 109334 64914 109426
rect 65082 109334 65466 109426
rect 65634 109334 66018 109426
rect 66186 109334 66570 109426
rect 66738 109334 67122 109426
rect 67290 109334 67674 109426
rect 67842 109334 68226 109426
rect 68394 109334 68778 109426
rect 68946 109334 69330 109426
rect 69498 109334 69882 109426
rect 70050 109334 70434 109426
rect 70602 109334 70986 109426
rect 71154 109334 71538 109426
rect 71706 109334 72090 109426
rect 72258 109334 72642 109426
rect 72810 109334 73194 109426
rect 73362 109334 73746 109426
rect 73914 109334 74298 109426
rect 74466 109334 74850 109426
rect 75018 109334 75402 109426
rect 75570 109334 75954 109426
rect 76122 109334 82032 109426
rect 1030 856 82032 109334
rect 1030 734 2814 856
rect 2982 734 3642 856
rect 3810 734 4470 856
rect 4638 734 5298 856
rect 5466 734 6126 856
rect 6294 734 6954 856
rect 7122 734 7782 856
rect 7950 734 8610 856
rect 8778 734 9438 856
rect 9606 734 10266 856
rect 10434 734 11094 856
rect 11262 734 11922 856
rect 12090 734 12750 856
rect 12918 734 13578 856
rect 13746 734 14406 856
rect 14574 734 15234 856
rect 15402 734 16062 856
rect 16230 734 16890 856
rect 17058 734 17718 856
rect 17886 734 18546 856
rect 18714 734 19374 856
rect 19542 734 20202 856
rect 20370 734 21030 856
rect 21198 734 21858 856
rect 22026 734 22686 856
rect 22854 734 23514 856
rect 23682 734 24342 856
rect 24510 734 25170 856
rect 25338 734 25998 856
rect 26166 734 26826 856
rect 26994 734 27654 856
rect 27822 734 28482 856
rect 28650 734 29310 856
rect 29478 734 30138 856
rect 30306 734 30966 856
rect 31134 734 31794 856
rect 31962 734 32622 856
rect 32790 734 33450 856
rect 33618 734 34278 856
rect 34446 734 35106 856
rect 35274 734 35934 856
rect 36102 734 36762 856
rect 36930 734 37590 856
rect 37758 734 38418 856
rect 38586 734 39246 856
rect 39414 734 40074 856
rect 40242 734 40902 856
rect 41070 734 41730 856
rect 41898 734 42558 856
rect 42726 734 43386 856
rect 43554 734 44214 856
rect 44382 734 45042 856
rect 45210 734 45870 856
rect 46038 734 46698 856
rect 46866 734 47526 856
rect 47694 734 48354 856
rect 48522 734 49182 856
rect 49350 734 50010 856
rect 50178 734 50838 856
rect 51006 734 51666 856
rect 51834 734 52494 856
rect 52662 734 53322 856
rect 53490 734 54150 856
rect 54318 734 54978 856
rect 55146 734 55806 856
rect 55974 734 56634 856
rect 56802 734 57462 856
rect 57630 734 58290 856
rect 58458 734 59118 856
rect 59286 734 59946 856
rect 60114 734 60774 856
rect 60942 734 61602 856
rect 61770 734 62430 856
rect 62598 734 63258 856
rect 63426 734 64086 856
rect 64254 734 64914 856
rect 65082 734 65742 856
rect 65910 734 66570 856
rect 66738 734 67398 856
rect 67566 734 68226 856
rect 68394 734 69054 856
rect 69222 734 69882 856
rect 70050 734 70710 856
rect 70878 734 71538 856
rect 71706 734 72366 856
rect 72534 734 73194 856
rect 73362 734 74022 856
rect 74190 734 74850 856
rect 75018 734 75678 856
rect 75846 734 76506 856
rect 76674 734 77334 856
rect 77502 734 78162 856
rect 78330 734 78990 856
rect 79158 734 82032 856
<< metal3 >>
rect 0 107992 800 108112
rect 81246 107176 82046 107296
rect 0 106360 800 106480
rect 81246 105544 82046 105664
rect 0 104728 800 104848
rect 81246 103912 82046 104032
rect 0 103096 800 103216
rect 81246 102280 82046 102400
rect 0 101464 800 101584
rect 81246 100648 82046 100768
rect 0 99832 800 99952
rect 81246 99016 82046 99136
rect 0 98200 800 98320
rect 81246 97384 82046 97504
rect 0 96568 800 96688
rect 81246 95752 82046 95872
rect 0 94936 800 95056
rect 81246 94120 82046 94240
rect 0 93304 800 93424
rect 81246 92488 82046 92608
rect 0 91672 800 91792
rect 81246 90856 82046 90976
rect 0 90040 800 90160
rect 81246 89224 82046 89344
rect 0 88408 800 88528
rect 81246 87592 82046 87712
rect 0 86776 800 86896
rect 81246 85960 82046 86080
rect 0 85144 800 85264
rect 81246 84328 82046 84448
rect 0 83512 800 83632
rect 81246 82696 82046 82816
rect 0 81880 800 82000
rect 81246 81064 82046 81184
rect 0 80248 800 80368
rect 81246 79432 82046 79552
rect 0 78616 800 78736
rect 81246 77800 82046 77920
rect 0 76984 800 77104
rect 81246 76168 82046 76288
rect 0 75352 800 75472
rect 81246 74536 82046 74656
rect 0 73720 800 73840
rect 81246 72904 82046 73024
rect 0 72088 800 72208
rect 81246 71272 82046 71392
rect 0 70456 800 70576
rect 81246 69640 82046 69760
rect 0 68824 800 68944
rect 81246 68008 82046 68128
rect 0 67192 800 67312
rect 81246 66376 82046 66496
rect 0 65560 800 65680
rect 81246 64744 82046 64864
rect 0 63928 800 64048
rect 81246 63112 82046 63232
rect 0 62296 800 62416
rect 81246 61480 82046 61600
rect 0 60664 800 60784
rect 81246 59848 82046 59968
rect 0 59032 800 59152
rect 81246 58216 82046 58336
rect 0 57400 800 57520
rect 81246 56584 82046 56704
rect 0 55768 800 55888
rect 81246 54952 82046 55072
rect 0 54136 800 54256
rect 81246 53320 82046 53440
rect 0 52504 800 52624
rect 81246 51688 82046 51808
rect 0 50872 800 50992
rect 81246 50056 82046 50176
rect 0 49240 800 49360
rect 81246 48424 82046 48544
rect 0 47608 800 47728
rect 81246 46792 82046 46912
rect 0 45976 800 46096
rect 81246 45160 82046 45280
rect 0 44344 800 44464
rect 81246 43528 82046 43648
rect 0 42712 800 42832
rect 81246 41896 82046 42016
rect 0 41080 800 41200
rect 81246 40264 82046 40384
rect 0 39448 800 39568
rect 81246 38632 82046 38752
rect 0 37816 800 37936
rect 81246 37000 82046 37120
rect 0 36184 800 36304
rect 81246 35368 82046 35488
rect 0 34552 800 34672
rect 81246 33736 82046 33856
rect 0 32920 800 33040
rect 81246 32104 82046 32224
rect 0 31288 800 31408
rect 81246 30472 82046 30592
rect 0 29656 800 29776
rect 81246 28840 82046 28960
rect 0 28024 800 28144
rect 81246 27208 82046 27328
rect 0 26392 800 26512
rect 81246 25576 82046 25696
rect 0 24760 800 24880
rect 81246 23944 82046 24064
rect 0 23128 800 23248
rect 81246 22312 82046 22432
rect 0 21496 800 21616
rect 81246 20680 82046 20800
rect 0 19864 800 19984
rect 81246 19048 82046 19168
rect 0 18232 800 18352
rect 81246 17416 82046 17536
rect 0 16600 800 16720
rect 81246 15784 82046 15904
rect 0 14968 800 15088
rect 81246 14152 82046 14272
rect 0 13336 800 13456
rect 81246 12520 82046 12640
rect 0 11704 800 11824
rect 81246 10888 82046 11008
rect 0 10072 800 10192
rect 81246 9256 82046 9376
rect 0 8440 800 8560
rect 81246 7624 82046 7744
rect 0 6808 800 6928
rect 81246 5992 82046 6112
rect 0 5176 800 5296
rect 81246 4360 82046 4480
rect 0 3544 800 3664
rect 81246 2728 82046 2848
rect 0 1912 800 2032
<< obsm3 >>
rect 880 107912 81959 108085
rect 800 107376 81959 107912
rect 800 107096 81166 107376
rect 800 106560 81959 107096
rect 880 106280 81959 106560
rect 800 105744 81959 106280
rect 800 105464 81166 105744
rect 800 104928 81959 105464
rect 880 104648 81959 104928
rect 800 104112 81959 104648
rect 800 103832 81166 104112
rect 800 103296 81959 103832
rect 880 103016 81959 103296
rect 800 102480 81959 103016
rect 800 102200 81166 102480
rect 800 101664 81959 102200
rect 880 101384 81959 101664
rect 800 100848 81959 101384
rect 800 100568 81166 100848
rect 800 100032 81959 100568
rect 880 99752 81959 100032
rect 800 99216 81959 99752
rect 800 98936 81166 99216
rect 800 98400 81959 98936
rect 880 98120 81959 98400
rect 800 97584 81959 98120
rect 800 97304 81166 97584
rect 800 96768 81959 97304
rect 880 96488 81959 96768
rect 800 95952 81959 96488
rect 800 95672 81166 95952
rect 800 95136 81959 95672
rect 880 94856 81959 95136
rect 800 94320 81959 94856
rect 800 94040 81166 94320
rect 800 93504 81959 94040
rect 880 93224 81959 93504
rect 800 92688 81959 93224
rect 800 92408 81166 92688
rect 800 91872 81959 92408
rect 880 91592 81959 91872
rect 800 91056 81959 91592
rect 800 90776 81166 91056
rect 800 90240 81959 90776
rect 880 89960 81959 90240
rect 800 89424 81959 89960
rect 800 89144 81166 89424
rect 800 88608 81959 89144
rect 880 88328 81959 88608
rect 800 87792 81959 88328
rect 800 87512 81166 87792
rect 800 86976 81959 87512
rect 880 86696 81959 86976
rect 800 86160 81959 86696
rect 800 85880 81166 86160
rect 800 85344 81959 85880
rect 880 85064 81959 85344
rect 800 84528 81959 85064
rect 800 84248 81166 84528
rect 800 83712 81959 84248
rect 880 83432 81959 83712
rect 800 82896 81959 83432
rect 800 82616 81166 82896
rect 800 82080 81959 82616
rect 880 81800 81959 82080
rect 800 81264 81959 81800
rect 800 80984 81166 81264
rect 800 80448 81959 80984
rect 880 80168 81959 80448
rect 800 79632 81959 80168
rect 800 79352 81166 79632
rect 800 78816 81959 79352
rect 880 78536 81959 78816
rect 800 78000 81959 78536
rect 800 77720 81166 78000
rect 800 77184 81959 77720
rect 880 76904 81959 77184
rect 800 76368 81959 76904
rect 800 76088 81166 76368
rect 800 75552 81959 76088
rect 880 75272 81959 75552
rect 800 74736 81959 75272
rect 800 74456 81166 74736
rect 800 73920 81959 74456
rect 880 73640 81959 73920
rect 800 73104 81959 73640
rect 800 72824 81166 73104
rect 800 72288 81959 72824
rect 880 72008 81959 72288
rect 800 71472 81959 72008
rect 800 71192 81166 71472
rect 800 70656 81959 71192
rect 880 70376 81959 70656
rect 800 69840 81959 70376
rect 800 69560 81166 69840
rect 800 69024 81959 69560
rect 880 68744 81959 69024
rect 800 68208 81959 68744
rect 800 67928 81166 68208
rect 800 67392 81959 67928
rect 880 67112 81959 67392
rect 800 66576 81959 67112
rect 800 66296 81166 66576
rect 800 65760 81959 66296
rect 880 65480 81959 65760
rect 800 64944 81959 65480
rect 800 64664 81166 64944
rect 800 64128 81959 64664
rect 880 63848 81959 64128
rect 800 63312 81959 63848
rect 800 63032 81166 63312
rect 800 62496 81959 63032
rect 880 62216 81959 62496
rect 800 61680 81959 62216
rect 800 61400 81166 61680
rect 800 60864 81959 61400
rect 880 60584 81959 60864
rect 800 60048 81959 60584
rect 800 59768 81166 60048
rect 800 59232 81959 59768
rect 880 58952 81959 59232
rect 800 58416 81959 58952
rect 800 58136 81166 58416
rect 800 57600 81959 58136
rect 880 57320 81959 57600
rect 800 56784 81959 57320
rect 800 56504 81166 56784
rect 800 55968 81959 56504
rect 880 55688 81959 55968
rect 800 55152 81959 55688
rect 800 54872 81166 55152
rect 800 54336 81959 54872
rect 880 54056 81959 54336
rect 800 53520 81959 54056
rect 800 53240 81166 53520
rect 800 52704 81959 53240
rect 880 52424 81959 52704
rect 800 51888 81959 52424
rect 800 51608 81166 51888
rect 800 51072 81959 51608
rect 880 50792 81959 51072
rect 800 50256 81959 50792
rect 800 49976 81166 50256
rect 800 49440 81959 49976
rect 880 49160 81959 49440
rect 800 48624 81959 49160
rect 800 48344 81166 48624
rect 800 47808 81959 48344
rect 880 47528 81959 47808
rect 800 46992 81959 47528
rect 800 46712 81166 46992
rect 800 46176 81959 46712
rect 880 45896 81959 46176
rect 800 45360 81959 45896
rect 800 45080 81166 45360
rect 800 44544 81959 45080
rect 880 44264 81959 44544
rect 800 43728 81959 44264
rect 800 43448 81166 43728
rect 800 42912 81959 43448
rect 880 42632 81959 42912
rect 800 42096 81959 42632
rect 800 41816 81166 42096
rect 800 41280 81959 41816
rect 880 41000 81959 41280
rect 800 40464 81959 41000
rect 800 40184 81166 40464
rect 800 39648 81959 40184
rect 880 39368 81959 39648
rect 800 38832 81959 39368
rect 800 38552 81166 38832
rect 800 38016 81959 38552
rect 880 37736 81959 38016
rect 800 37200 81959 37736
rect 800 36920 81166 37200
rect 800 36384 81959 36920
rect 880 36104 81959 36384
rect 800 35568 81959 36104
rect 800 35288 81166 35568
rect 800 34752 81959 35288
rect 880 34472 81959 34752
rect 800 33936 81959 34472
rect 800 33656 81166 33936
rect 800 33120 81959 33656
rect 880 32840 81959 33120
rect 800 32304 81959 32840
rect 800 32024 81166 32304
rect 800 31488 81959 32024
rect 880 31208 81959 31488
rect 800 30672 81959 31208
rect 800 30392 81166 30672
rect 800 29856 81959 30392
rect 880 29576 81959 29856
rect 800 29040 81959 29576
rect 800 28760 81166 29040
rect 800 28224 81959 28760
rect 880 27944 81959 28224
rect 800 27408 81959 27944
rect 800 27128 81166 27408
rect 800 26592 81959 27128
rect 880 26312 81959 26592
rect 800 25776 81959 26312
rect 800 25496 81166 25776
rect 800 24960 81959 25496
rect 880 24680 81959 24960
rect 800 24144 81959 24680
rect 800 23864 81166 24144
rect 800 23328 81959 23864
rect 880 23048 81959 23328
rect 800 22512 81959 23048
rect 800 22232 81166 22512
rect 800 21696 81959 22232
rect 880 21416 81959 21696
rect 800 20880 81959 21416
rect 800 20600 81166 20880
rect 800 20064 81959 20600
rect 880 19784 81959 20064
rect 800 19248 81959 19784
rect 800 18968 81166 19248
rect 800 18432 81959 18968
rect 880 18152 81959 18432
rect 800 17616 81959 18152
rect 800 17336 81166 17616
rect 800 16800 81959 17336
rect 880 16520 81959 16800
rect 800 15984 81959 16520
rect 800 15704 81166 15984
rect 800 15168 81959 15704
rect 880 14888 81959 15168
rect 800 14352 81959 14888
rect 800 14072 81166 14352
rect 800 13536 81959 14072
rect 880 13256 81959 13536
rect 800 12720 81959 13256
rect 800 12440 81166 12720
rect 800 11904 81959 12440
rect 880 11624 81959 11904
rect 800 11088 81959 11624
rect 800 10808 81166 11088
rect 800 10272 81959 10808
rect 880 9992 81959 10272
rect 800 9456 81959 9992
rect 800 9176 81166 9456
rect 800 8640 81959 9176
rect 880 8360 81959 8640
rect 800 7824 81959 8360
rect 800 7544 81166 7824
rect 800 7008 81959 7544
rect 880 6728 81959 7008
rect 800 6192 81959 6728
rect 800 5912 81166 6192
rect 800 5376 81959 5912
rect 880 5096 81959 5376
rect 800 4560 81959 5096
rect 800 4280 81166 4560
rect 800 3744 81959 4280
rect 880 3464 81959 3744
rect 800 2928 81959 3464
rect 800 2648 81166 2928
rect 800 2112 81959 2648
rect 880 1939 81959 2112
<< metal4 >>
rect 4208 2128 4528 107760
rect 11888 2128 12208 107760
rect 19568 2128 19888 107760
rect 27248 2128 27568 107760
rect 34928 2128 35248 107760
rect 42608 2128 42928 107760
rect 50288 2128 50608 107760
rect 57968 2128 58288 107760
rect 65648 2128 65968 107760
rect 73328 2128 73648 107760
<< obsm4 >>
rect 1899 2347 4128 106997
rect 4608 2347 11808 106997
rect 12288 2347 19488 106997
rect 19968 2347 27168 106997
rect 27648 2347 34848 106997
rect 35328 2347 42528 106997
rect 43008 2347 50208 106997
rect 50688 2347 57888 106997
rect 58368 2347 65568 106997
rect 66048 2347 73248 106997
rect 73728 2347 79981 106997
<< labels >>
rlabel metal4 s 11888 2128 12208 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27248 2128 27568 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 42608 2128 42928 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 57968 2128 58288 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 73328 2128 73648 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 1912 800 2032 6 debug_in
port 3 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 debug_mode
port 4 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 debug_oeb
port 5 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 debug_out
port 6 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 irq[0]
port 7 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 irq[1]
port 8 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 irq[2]
port 9 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 mask_rev_in[0]
port 10 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 mask_rev_in[10]
port 11 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 mask_rev_in[11]
port 12 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 mask_rev_in[12]
port 13 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 mask_rev_in[13]
port 14 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 mask_rev_in[14]
port 15 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 mask_rev_in[15]
port 16 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 mask_rev_in[16]
port 17 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 mask_rev_in[17]
port 18 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 mask_rev_in[18]
port 19 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 mask_rev_in[19]
port 20 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 mask_rev_in[1]
port 21 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 mask_rev_in[20]
port 22 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 mask_rev_in[21]
port 23 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 mask_rev_in[22]
port 24 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 mask_rev_in[23]
port 25 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 mask_rev_in[24]
port 26 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 mask_rev_in[25]
port 27 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 mask_rev_in[26]
port 28 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 mask_rev_in[27]
port 29 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 mask_rev_in[28]
port 30 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 mask_rev_in[29]
port 31 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 mask_rev_in[2]
port 32 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 mask_rev_in[30]
port 33 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 mask_rev_in[31]
port 34 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 mask_rev_in[3]
port 35 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 mask_rev_in[4]
port 36 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 mask_rev_in[5]
port 37 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 mask_rev_in[6]
port 38 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 mask_rev_in[7]
port 39 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 mask_rev_in[8]
port 40 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 mask_rev_in[9]
port 41 nsew signal input
rlabel metal3 s 81246 10888 82046 11008 6 mgmt_gpio_in[0]
port 42 nsew signal input
rlabel metal3 s 81246 59848 82046 59968 6 mgmt_gpio_in[10]
port 43 nsew signal input
rlabel metal3 s 81246 64744 82046 64864 6 mgmt_gpio_in[11]
port 44 nsew signal input
rlabel metal3 s 81246 69640 82046 69760 6 mgmt_gpio_in[12]
port 45 nsew signal input
rlabel metal3 s 81246 74536 82046 74656 6 mgmt_gpio_in[13]
port 46 nsew signal input
rlabel metal3 s 81246 79432 82046 79552 6 mgmt_gpio_in[14]
port 47 nsew signal input
rlabel metal3 s 81246 84328 82046 84448 6 mgmt_gpio_in[15]
port 48 nsew signal input
rlabel metal3 s 81246 89224 82046 89344 6 mgmt_gpio_in[16]
port 49 nsew signal input
rlabel metal3 s 81246 94120 82046 94240 6 mgmt_gpio_in[17]
port 50 nsew signal input
rlabel metal3 s 81246 99016 82046 99136 6 mgmt_gpio_in[18]
port 51 nsew signal input
rlabel metal3 s 81246 103912 82046 104032 6 mgmt_gpio_in[19]
port 52 nsew signal input
rlabel metal3 s 81246 15784 82046 15904 6 mgmt_gpio_in[1]
port 53 nsew signal input
rlabel metal2 s 46754 109390 46810 110190 6 mgmt_gpio_in[20]
port 54 nsew signal input
rlabel metal2 s 48410 109390 48466 110190 6 mgmt_gpio_in[21]
port 55 nsew signal input
rlabel metal2 s 50066 109390 50122 110190 6 mgmt_gpio_in[22]
port 56 nsew signal input
rlabel metal2 s 51722 109390 51778 110190 6 mgmt_gpio_in[23]
port 57 nsew signal input
rlabel metal2 s 53378 109390 53434 110190 6 mgmt_gpio_in[24]
port 58 nsew signal input
rlabel metal2 s 55034 109390 55090 110190 6 mgmt_gpio_in[25]
port 59 nsew signal input
rlabel metal2 s 56690 109390 56746 110190 6 mgmt_gpio_in[26]
port 60 nsew signal input
rlabel metal2 s 58346 109390 58402 110190 6 mgmt_gpio_in[27]
port 61 nsew signal input
rlabel metal2 s 60002 109390 60058 110190 6 mgmt_gpio_in[28]
port 62 nsew signal input
rlabel metal2 s 61658 109390 61714 110190 6 mgmt_gpio_in[29]
port 63 nsew signal input
rlabel metal3 s 81246 20680 82046 20800 6 mgmt_gpio_in[2]
port 64 nsew signal input
rlabel metal2 s 63314 109390 63370 110190 6 mgmt_gpio_in[30]
port 65 nsew signal input
rlabel metal2 s 64970 109390 65026 110190 6 mgmt_gpio_in[31]
port 66 nsew signal input
rlabel metal2 s 66626 109390 66682 110190 6 mgmt_gpio_in[32]
port 67 nsew signal input
rlabel metal2 s 68282 109390 68338 110190 6 mgmt_gpio_in[33]
port 68 nsew signal input
rlabel metal2 s 69938 109390 69994 110190 6 mgmt_gpio_in[34]
port 69 nsew signal input
rlabel metal2 s 71594 109390 71650 110190 6 mgmt_gpio_in[35]
port 70 nsew signal input
rlabel metal2 s 73250 109390 73306 110190 6 mgmt_gpio_in[36]
port 71 nsew signal input
rlabel metal2 s 74906 109390 74962 110190 6 mgmt_gpio_in[37]
port 72 nsew signal input
rlabel metal3 s 81246 25576 82046 25696 6 mgmt_gpio_in[3]
port 73 nsew signal input
rlabel metal3 s 81246 30472 82046 30592 6 mgmt_gpio_in[4]
port 74 nsew signal input
rlabel metal3 s 81246 35368 82046 35488 6 mgmt_gpio_in[5]
port 75 nsew signal input
rlabel metal3 s 81246 40264 82046 40384 6 mgmt_gpio_in[6]
port 76 nsew signal input
rlabel metal3 s 81246 45160 82046 45280 6 mgmt_gpio_in[7]
port 77 nsew signal input
rlabel metal3 s 81246 50056 82046 50176 6 mgmt_gpio_in[8]
port 78 nsew signal input
rlabel metal3 s 81246 54952 82046 55072 6 mgmt_gpio_in[9]
port 79 nsew signal input
rlabel metal3 s 81246 12520 82046 12640 6 mgmt_gpio_oeb[0]
port 80 nsew signal output
rlabel metal3 s 81246 61480 82046 61600 6 mgmt_gpio_oeb[10]
port 81 nsew signal output
rlabel metal3 s 81246 66376 82046 66496 6 mgmt_gpio_oeb[11]
port 82 nsew signal output
rlabel metal3 s 81246 71272 82046 71392 6 mgmt_gpio_oeb[12]
port 83 nsew signal output
rlabel metal3 s 81246 76168 82046 76288 6 mgmt_gpio_oeb[13]
port 84 nsew signal output
rlabel metal3 s 81246 81064 82046 81184 6 mgmt_gpio_oeb[14]
port 85 nsew signal output
rlabel metal3 s 81246 85960 82046 86080 6 mgmt_gpio_oeb[15]
port 86 nsew signal output
rlabel metal3 s 81246 90856 82046 90976 6 mgmt_gpio_oeb[16]
port 87 nsew signal output
rlabel metal3 s 81246 95752 82046 95872 6 mgmt_gpio_oeb[17]
port 88 nsew signal output
rlabel metal3 s 81246 100648 82046 100768 6 mgmt_gpio_oeb[18]
port 89 nsew signal output
rlabel metal3 s 81246 105544 82046 105664 6 mgmt_gpio_oeb[19]
port 90 nsew signal output
rlabel metal3 s 81246 17416 82046 17536 6 mgmt_gpio_oeb[1]
port 91 nsew signal output
rlabel metal2 s 47306 109390 47362 110190 6 mgmt_gpio_oeb[20]
port 92 nsew signal output
rlabel metal2 s 48962 109390 49018 110190 6 mgmt_gpio_oeb[21]
port 93 nsew signal output
rlabel metal2 s 50618 109390 50674 110190 6 mgmt_gpio_oeb[22]
port 94 nsew signal output
rlabel metal2 s 52274 109390 52330 110190 6 mgmt_gpio_oeb[23]
port 95 nsew signal output
rlabel metal2 s 53930 109390 53986 110190 6 mgmt_gpio_oeb[24]
port 96 nsew signal output
rlabel metal2 s 55586 109390 55642 110190 6 mgmt_gpio_oeb[25]
port 97 nsew signal output
rlabel metal2 s 57242 109390 57298 110190 6 mgmt_gpio_oeb[26]
port 98 nsew signal output
rlabel metal2 s 58898 109390 58954 110190 6 mgmt_gpio_oeb[27]
port 99 nsew signal output
rlabel metal2 s 60554 109390 60610 110190 6 mgmt_gpio_oeb[28]
port 100 nsew signal output
rlabel metal2 s 62210 109390 62266 110190 6 mgmt_gpio_oeb[29]
port 101 nsew signal output
rlabel metal3 s 81246 22312 82046 22432 6 mgmt_gpio_oeb[2]
port 102 nsew signal output
rlabel metal2 s 63866 109390 63922 110190 6 mgmt_gpio_oeb[30]
port 103 nsew signal output
rlabel metal2 s 65522 109390 65578 110190 6 mgmt_gpio_oeb[31]
port 104 nsew signal output
rlabel metal2 s 67178 109390 67234 110190 6 mgmt_gpio_oeb[32]
port 105 nsew signal output
rlabel metal2 s 68834 109390 68890 110190 6 mgmt_gpio_oeb[33]
port 106 nsew signal output
rlabel metal2 s 70490 109390 70546 110190 6 mgmt_gpio_oeb[34]
port 107 nsew signal output
rlabel metal2 s 72146 109390 72202 110190 6 mgmt_gpio_oeb[35]
port 108 nsew signal output
rlabel metal2 s 73802 109390 73858 110190 6 mgmt_gpio_oeb[36]
port 109 nsew signal output
rlabel metal2 s 75458 109390 75514 110190 6 mgmt_gpio_oeb[37]
port 110 nsew signal output
rlabel metal3 s 81246 27208 82046 27328 6 mgmt_gpio_oeb[3]
port 111 nsew signal output
rlabel metal3 s 81246 32104 82046 32224 6 mgmt_gpio_oeb[4]
port 112 nsew signal output
rlabel metal3 s 81246 37000 82046 37120 6 mgmt_gpio_oeb[5]
port 113 nsew signal output
rlabel metal3 s 81246 41896 82046 42016 6 mgmt_gpio_oeb[6]
port 114 nsew signal output
rlabel metal3 s 81246 46792 82046 46912 6 mgmt_gpio_oeb[7]
port 115 nsew signal output
rlabel metal3 s 81246 51688 82046 51808 6 mgmt_gpio_oeb[8]
port 116 nsew signal output
rlabel metal3 s 81246 56584 82046 56704 6 mgmt_gpio_oeb[9]
port 117 nsew signal output
rlabel metal3 s 81246 14152 82046 14272 6 mgmt_gpio_out[0]
port 118 nsew signal output
rlabel metal3 s 81246 63112 82046 63232 6 mgmt_gpio_out[10]
port 119 nsew signal output
rlabel metal3 s 81246 68008 82046 68128 6 mgmt_gpio_out[11]
port 120 nsew signal output
rlabel metal3 s 81246 72904 82046 73024 6 mgmt_gpio_out[12]
port 121 nsew signal output
rlabel metal3 s 81246 77800 82046 77920 6 mgmt_gpio_out[13]
port 122 nsew signal output
rlabel metal3 s 81246 82696 82046 82816 6 mgmt_gpio_out[14]
port 123 nsew signal output
rlabel metal3 s 81246 87592 82046 87712 6 mgmt_gpio_out[15]
port 124 nsew signal output
rlabel metal3 s 81246 92488 82046 92608 6 mgmt_gpio_out[16]
port 125 nsew signal output
rlabel metal3 s 81246 97384 82046 97504 6 mgmt_gpio_out[17]
port 126 nsew signal output
rlabel metal3 s 81246 102280 82046 102400 6 mgmt_gpio_out[18]
port 127 nsew signal output
rlabel metal3 s 81246 107176 82046 107296 6 mgmt_gpio_out[19]
port 128 nsew signal output
rlabel metal3 s 81246 19048 82046 19168 6 mgmt_gpio_out[1]
port 129 nsew signal output
rlabel metal2 s 47858 109390 47914 110190 6 mgmt_gpio_out[20]
port 130 nsew signal output
rlabel metal2 s 49514 109390 49570 110190 6 mgmt_gpio_out[21]
port 131 nsew signal output
rlabel metal2 s 51170 109390 51226 110190 6 mgmt_gpio_out[22]
port 132 nsew signal output
rlabel metal2 s 52826 109390 52882 110190 6 mgmt_gpio_out[23]
port 133 nsew signal output
rlabel metal2 s 54482 109390 54538 110190 6 mgmt_gpio_out[24]
port 134 nsew signal output
rlabel metal2 s 56138 109390 56194 110190 6 mgmt_gpio_out[25]
port 135 nsew signal output
rlabel metal2 s 57794 109390 57850 110190 6 mgmt_gpio_out[26]
port 136 nsew signal output
rlabel metal2 s 59450 109390 59506 110190 6 mgmt_gpio_out[27]
port 137 nsew signal output
rlabel metal2 s 61106 109390 61162 110190 6 mgmt_gpio_out[28]
port 138 nsew signal output
rlabel metal2 s 62762 109390 62818 110190 6 mgmt_gpio_out[29]
port 139 nsew signal output
rlabel metal3 s 81246 23944 82046 24064 6 mgmt_gpio_out[2]
port 140 nsew signal output
rlabel metal2 s 64418 109390 64474 110190 6 mgmt_gpio_out[30]
port 141 nsew signal output
rlabel metal2 s 66074 109390 66130 110190 6 mgmt_gpio_out[31]
port 142 nsew signal output
rlabel metal2 s 67730 109390 67786 110190 6 mgmt_gpio_out[32]
port 143 nsew signal output
rlabel metal2 s 69386 109390 69442 110190 6 mgmt_gpio_out[33]
port 144 nsew signal output
rlabel metal2 s 71042 109390 71098 110190 6 mgmt_gpio_out[34]
port 145 nsew signal output
rlabel metal2 s 72698 109390 72754 110190 6 mgmt_gpio_out[35]
port 146 nsew signal output
rlabel metal2 s 74354 109390 74410 110190 6 mgmt_gpio_out[36]
port 147 nsew signal output
rlabel metal2 s 76010 109390 76066 110190 6 mgmt_gpio_out[37]
port 148 nsew signal output
rlabel metal3 s 81246 28840 82046 28960 6 mgmt_gpio_out[3]
port 149 nsew signal output
rlabel metal3 s 81246 33736 82046 33856 6 mgmt_gpio_out[4]
port 150 nsew signal output
rlabel metal3 s 81246 38632 82046 38752 6 mgmt_gpio_out[5]
port 151 nsew signal output
rlabel metal3 s 81246 43528 82046 43648 6 mgmt_gpio_out[6]
port 152 nsew signal output
rlabel metal3 s 81246 48424 82046 48544 6 mgmt_gpio_out[7]
port 153 nsew signal output
rlabel metal3 s 81246 53320 82046 53440 6 mgmt_gpio_out[8]
port 154 nsew signal output
rlabel metal3 s 81246 58216 82046 58336 6 mgmt_gpio_out[9]
port 155 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 pad_flash_clk
port 156 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 pad_flash_clk_oeb
port 157 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 pad_flash_csb
port 158 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 pad_flash_csb_oeb
port 159 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 pad_flash_io0_di
port 160 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 pad_flash_io0_do
port 161 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 pad_flash_io0_ieb
port 162 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 pad_flash_io0_oeb
port 163 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 pad_flash_io1_di
port 164 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 pad_flash_io1_do
port 165 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 pad_flash_io1_ieb
port 166 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 pad_flash_io1_oeb
port 167 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 pll90_sel[0]
port 168 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 pll90_sel[1]
port 169 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 pll90_sel[2]
port 170 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 pll_bypass
port 171 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 pll_dco_ena
port 172 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 pll_div[0]
port 173 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 pll_div[1]
port 174 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 pll_div[2]
port 175 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 pll_div[3]
port 176 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 pll_div[4]
port 177 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 pll_ena
port 178 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 pll_sel[0]
port 179 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 pll_sel[1]
port 180 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 pll_sel[2]
port 181 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 pll_trim[0]
port 182 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 pll_trim[10]
port 183 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 pll_trim[11]
port 184 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 pll_trim[12]
port 185 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 pll_trim[13]
port 186 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 pll_trim[14]
port 187 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 pll_trim[15]
port 188 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 pll_trim[16]
port 189 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 pll_trim[17]
port 190 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 pll_trim[18]
port 191 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 pll_trim[19]
port 192 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 pll_trim[1]
port 193 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 pll_trim[20]
port 194 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 pll_trim[21]
port 195 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 pll_trim[22]
port 196 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 pll_trim[23]
port 197 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 pll_trim[24]
port 198 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 pll_trim[25]
port 199 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 pll_trim[2]
port 200 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 pll_trim[3]
port 201 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 pll_trim[4]
port 202 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 pll_trim[5]
port 203 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 pll_trim[6]
port 204 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 pll_trim[7]
port 205 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 pll_trim[8]
port 206 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 pll_trim[9]
port 207 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 porb
port 208 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 pwr_ctrl_out[0]
port 209 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 pwr_ctrl_out[1]
port 210 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 pwr_ctrl_out[2]
port 211 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 pwr_ctrl_out[3]
port 212 nsew signal output
rlabel metal3 s 0 26392 800 26512 6 qspi_enabled
port 213 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 reset
port 214 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 ser_rx
port 215 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 ser_tx
port 216 nsew signal input
rlabel metal3 s 81246 2728 82046 2848 6 serial_clock
port 217 nsew signal output
rlabel metal3 s 81246 7624 82046 7744 6 serial_data_1
port 218 nsew signal output
rlabel metal3 s 81246 9256 82046 9376 6 serial_data_2
port 219 nsew signal output
rlabel metal3 s 81246 5992 82046 6112 6 serial_load
port 220 nsew signal output
rlabel metal3 s 81246 4360 82046 4480 6 serial_resetn
port 221 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 spi_csb
port 222 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 spi_enabled
port 223 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 spi_sck
port 224 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 spi_sdi
port 225 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 spi_sdo
port 226 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 spi_sdoenb
port 227 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 spimemio_flash_clk
port 228 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 spimemio_flash_csb
port 229 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 spimemio_flash_io0_di
port 230 nsew signal output
rlabel metal3 s 0 91672 800 91792 6 spimemio_flash_io0_do
port 231 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 spimemio_flash_io0_oeb
port 232 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 spimemio_flash_io1_di
port 233 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 spimemio_flash_io1_do
port 234 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 spimemio_flash_io1_oeb
port 235 nsew signal input
rlabel metal3 s 0 99832 800 99952 6 spimemio_flash_io2_di
port 236 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 spimemio_flash_io2_do
port 237 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 spimemio_flash_io2_oeb
port 238 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 spimemio_flash_io3_di
port 239 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 spimemio_flash_io3_do
port 240 nsew signal input
rlabel metal3 s 0 107992 800 108112 6 spimemio_flash_io3_oeb
port 241 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 trap
port 242 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 uart_enabled
port 243 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 user_clock
port 244 nsew signal input
rlabel metal2 s 44546 109390 44602 110190 6 usr1_vcc_pwrgood
port 245 nsew signal input
rlabel metal2 s 45650 109390 45706 110190 6 usr1_vdd_pwrgood
port 246 nsew signal input
rlabel metal2 s 45098 109390 45154 110190 6 usr2_vcc_pwrgood
port 247 nsew signal input
rlabel metal2 s 46202 109390 46258 110190 6 usr2_vdd_pwrgood
port 248 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 wb_ack_o
port 249 nsew signal output
rlabel metal2 s 5906 109390 5962 110190 6 wb_adr_i[0]
port 250 nsew signal input
rlabel metal2 s 11426 109390 11482 110190 6 wb_adr_i[10]
port 251 nsew signal input
rlabel metal2 s 11978 109390 12034 110190 6 wb_adr_i[11]
port 252 nsew signal input
rlabel metal2 s 12530 109390 12586 110190 6 wb_adr_i[12]
port 253 nsew signal input
rlabel metal2 s 13082 109390 13138 110190 6 wb_adr_i[13]
port 254 nsew signal input
rlabel metal2 s 13634 109390 13690 110190 6 wb_adr_i[14]
port 255 nsew signal input
rlabel metal2 s 14186 109390 14242 110190 6 wb_adr_i[15]
port 256 nsew signal input
rlabel metal2 s 14738 109390 14794 110190 6 wb_adr_i[16]
port 257 nsew signal input
rlabel metal2 s 15290 109390 15346 110190 6 wb_adr_i[17]
port 258 nsew signal input
rlabel metal2 s 15842 109390 15898 110190 6 wb_adr_i[18]
port 259 nsew signal input
rlabel metal2 s 16394 109390 16450 110190 6 wb_adr_i[19]
port 260 nsew signal input
rlabel metal2 s 6458 109390 6514 110190 6 wb_adr_i[1]
port 261 nsew signal input
rlabel metal2 s 16946 109390 17002 110190 6 wb_adr_i[20]
port 262 nsew signal input
rlabel metal2 s 17498 109390 17554 110190 6 wb_adr_i[21]
port 263 nsew signal input
rlabel metal2 s 18050 109390 18106 110190 6 wb_adr_i[22]
port 264 nsew signal input
rlabel metal2 s 18602 109390 18658 110190 6 wb_adr_i[23]
port 265 nsew signal input
rlabel metal2 s 19154 109390 19210 110190 6 wb_adr_i[24]
port 266 nsew signal input
rlabel metal2 s 19706 109390 19762 110190 6 wb_adr_i[25]
port 267 nsew signal input
rlabel metal2 s 20258 109390 20314 110190 6 wb_adr_i[26]
port 268 nsew signal input
rlabel metal2 s 20810 109390 20866 110190 6 wb_adr_i[27]
port 269 nsew signal input
rlabel metal2 s 21362 109390 21418 110190 6 wb_adr_i[28]
port 270 nsew signal input
rlabel metal2 s 21914 109390 21970 110190 6 wb_adr_i[29]
port 271 nsew signal input
rlabel metal2 s 7010 109390 7066 110190 6 wb_adr_i[2]
port 272 nsew signal input
rlabel metal2 s 22466 109390 22522 110190 6 wb_adr_i[30]
port 273 nsew signal input
rlabel metal2 s 23018 109390 23074 110190 6 wb_adr_i[31]
port 274 nsew signal input
rlabel metal2 s 7562 109390 7618 110190 6 wb_adr_i[3]
port 275 nsew signal input
rlabel metal2 s 8114 109390 8170 110190 6 wb_adr_i[4]
port 276 nsew signal input
rlabel metal2 s 8666 109390 8722 110190 6 wb_adr_i[5]
port 277 nsew signal input
rlabel metal2 s 9218 109390 9274 110190 6 wb_adr_i[6]
port 278 nsew signal input
rlabel metal2 s 9770 109390 9826 110190 6 wb_adr_i[7]
port 279 nsew signal input
rlabel metal2 s 10322 109390 10378 110190 6 wb_adr_i[8]
port 280 nsew signal input
rlabel metal2 s 10874 109390 10930 110190 6 wb_adr_i[9]
port 281 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 wb_clk_i
port 282 nsew signal input
rlabel metal2 s 43994 109390 44050 110190 6 wb_cyc_i
port 283 nsew signal input
rlabel metal2 s 23570 109390 23626 110190 6 wb_dat_i[0]
port 284 nsew signal input
rlabel metal2 s 29090 109390 29146 110190 6 wb_dat_i[10]
port 285 nsew signal input
rlabel metal2 s 29642 109390 29698 110190 6 wb_dat_i[11]
port 286 nsew signal input
rlabel metal2 s 30194 109390 30250 110190 6 wb_dat_i[12]
port 287 nsew signal input
rlabel metal2 s 30746 109390 30802 110190 6 wb_dat_i[13]
port 288 nsew signal input
rlabel metal2 s 31298 109390 31354 110190 6 wb_dat_i[14]
port 289 nsew signal input
rlabel metal2 s 31850 109390 31906 110190 6 wb_dat_i[15]
port 290 nsew signal input
rlabel metal2 s 32402 109390 32458 110190 6 wb_dat_i[16]
port 291 nsew signal input
rlabel metal2 s 32954 109390 33010 110190 6 wb_dat_i[17]
port 292 nsew signal input
rlabel metal2 s 33506 109390 33562 110190 6 wb_dat_i[18]
port 293 nsew signal input
rlabel metal2 s 34058 109390 34114 110190 6 wb_dat_i[19]
port 294 nsew signal input
rlabel metal2 s 24122 109390 24178 110190 6 wb_dat_i[1]
port 295 nsew signal input
rlabel metal2 s 34610 109390 34666 110190 6 wb_dat_i[20]
port 296 nsew signal input
rlabel metal2 s 35162 109390 35218 110190 6 wb_dat_i[21]
port 297 nsew signal input
rlabel metal2 s 35714 109390 35770 110190 6 wb_dat_i[22]
port 298 nsew signal input
rlabel metal2 s 36266 109390 36322 110190 6 wb_dat_i[23]
port 299 nsew signal input
rlabel metal2 s 36818 109390 36874 110190 6 wb_dat_i[24]
port 300 nsew signal input
rlabel metal2 s 37370 109390 37426 110190 6 wb_dat_i[25]
port 301 nsew signal input
rlabel metal2 s 37922 109390 37978 110190 6 wb_dat_i[26]
port 302 nsew signal input
rlabel metal2 s 38474 109390 38530 110190 6 wb_dat_i[27]
port 303 nsew signal input
rlabel metal2 s 39026 109390 39082 110190 6 wb_dat_i[28]
port 304 nsew signal input
rlabel metal2 s 39578 109390 39634 110190 6 wb_dat_i[29]
port 305 nsew signal input
rlabel metal2 s 24674 109390 24730 110190 6 wb_dat_i[2]
port 306 nsew signal input
rlabel metal2 s 40130 109390 40186 110190 6 wb_dat_i[30]
port 307 nsew signal input
rlabel metal2 s 40682 109390 40738 110190 6 wb_dat_i[31]
port 308 nsew signal input
rlabel metal2 s 25226 109390 25282 110190 6 wb_dat_i[3]
port 309 nsew signal input
rlabel metal2 s 25778 109390 25834 110190 6 wb_dat_i[4]
port 310 nsew signal input
rlabel metal2 s 26330 109390 26386 110190 6 wb_dat_i[5]
port 311 nsew signal input
rlabel metal2 s 26882 109390 26938 110190 6 wb_dat_i[6]
port 312 nsew signal input
rlabel metal2 s 27434 109390 27490 110190 6 wb_dat_i[7]
port 313 nsew signal input
rlabel metal2 s 27986 109390 28042 110190 6 wb_dat_i[8]
port 314 nsew signal input
rlabel metal2 s 28538 109390 28594 110190 6 wb_dat_i[9]
port 315 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 wb_dat_o[0]
port 316 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 wb_dat_o[10]
port 317 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 wb_dat_o[11]
port 318 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 wb_dat_o[12]
port 319 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 wb_dat_o[13]
port 320 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 wb_dat_o[14]
port 321 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 wb_dat_o[15]
port 322 nsew signal output
rlabel metal3 s 0 60664 800 60784 6 wb_dat_o[16]
port 323 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 wb_dat_o[17]
port 324 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 wb_dat_o[18]
port 325 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 wb_dat_o[19]
port 326 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 wb_dat_o[1]
port 327 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 wb_dat_o[20]
port 328 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 wb_dat_o[21]
port 329 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 wb_dat_o[22]
port 330 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 wb_dat_o[23]
port 331 nsew signal output
rlabel metal3 s 0 73720 800 73840 6 wb_dat_o[24]
port 332 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 wb_dat_o[25]
port 333 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 wb_dat_o[26]
port 334 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 wb_dat_o[27]
port 335 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 wb_dat_o[28]
port 336 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 wb_dat_o[29]
port 337 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 wb_dat_o[2]
port 338 nsew signal output
rlabel metal3 s 0 83512 800 83632 6 wb_dat_o[30]
port 339 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 wb_dat_o[31]
port 340 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 wb_dat_o[3]
port 341 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 wb_dat_o[4]
port 342 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 wb_dat_o[5]
port 343 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 wb_dat_o[6]
port 344 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 wb_dat_o[7]
port 345 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 wb_dat_o[8]
port 346 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 wb_dat_o[9]
port 347 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 wb_rstn_i
port 348 nsew signal input
rlabel metal2 s 41234 109390 41290 110190 6 wb_sel_i[0]
port 349 nsew signal input
rlabel metal2 s 41786 109390 41842 110190 6 wb_sel_i[1]
port 350 nsew signal input
rlabel metal2 s 42338 109390 42394 110190 6 wb_sel_i[2]
port 351 nsew signal input
rlabel metal2 s 42890 109390 42946 110190 6 wb_sel_i[3]
port 352 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 wb_stb_i
port 353 nsew signal input
rlabel metal2 s 43442 109390 43498 110190 6 wb_we_i
port 354 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 82046 110190
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27092910
string GDS_FILE /home/hosni/caravel-redesign-2/caravel/openlane/housekeeping/runs/23_04_09_06_22/results/signoff/housekeeping.magic.gds
string GDS_START 1217680
<< end >>

