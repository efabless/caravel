magic
tech sky130A
timestamp 1608325192
<< checkpaint >>
rect 7176 6798 15816 6886
rect 6615 6791 15816 6798
rect 6306 3466 15816 6791
rect 6306 3371 15698 3466
rect 6486 3367 15698 3371
rect 6486 3339 15126 3367
rect -630 -630 8010 2790
<< metal5 >>
rect 3060 7740 3960 7920
rect 1440 7200 1980 7380
rect 1260 7020 2340 7200
rect 2880 7020 4140 7740
rect 5040 7200 5580 7380
rect 4680 7020 5760 7200
rect 1260 6840 2520 7020
rect 2700 6840 4320 7020
rect 4500 6840 5760 7020
rect 1260 6660 5760 6840
rect 1440 6300 5580 6660
rect 1620 6120 5400 6300
rect 1800 5940 5280 6120
rect 7056 6101 7356 6161
rect 7776 6101 8076 6161
rect 8436 6101 8856 6161
rect 9096 6101 9516 6161
rect 10296 6101 10716 6161
rect 11016 6101 11316 6161
rect 6996 6041 7416 6101
rect 7716 6041 8136 6101
rect 1620 5760 3060 5940
rect 3960 5760 5400 5940
rect 6936 5921 7476 6041
rect 900 5580 2880 5760
rect 4140 5580 6120 5760
rect 540 4680 2700 5580
rect 4320 4680 6300 5580
rect 6936 5501 7116 5921
rect 7296 5501 7476 5921
rect 6936 5381 7476 5501
rect 7656 5921 8196 6041
rect 7656 5501 7836 5921
rect 8016 5501 8196 5921
rect 7656 5381 8196 5501
rect 8376 5981 8916 6101
rect 8376 5801 8556 5981
rect 8736 5801 8916 5981
rect 8376 5681 8916 5801
rect 9096 6041 9576 6101
rect 10236 6041 10716 6101
rect 10956 6041 11376 6101
rect 9096 5921 9636 6041
rect 8376 5621 8856 5681
rect 8376 5441 8556 5621
rect 6996 5321 7416 5381
rect 7656 5321 8136 5381
rect 8376 5321 8916 5441
rect 7056 5261 7356 5321
rect 7656 5261 8076 5321
rect 8436 5261 8916 5321
rect 9096 5261 9276 5921
rect 9456 5261 9636 5921
rect 10176 5981 10716 6041
rect 10176 5801 10416 5981
rect 10896 5921 11436 6041
rect 10176 5741 10596 5801
rect 10236 5681 10656 5741
rect 10296 5621 10716 5681
rect 10476 5441 10716 5621
rect 10176 5381 10716 5441
rect 10896 5501 11076 5921
rect 11256 5501 11436 5921
rect 10896 5381 11436 5501
rect 11616 5501 11796 6161
rect 11976 5501 12156 6161
rect 11616 5381 12156 5501
rect 12336 6101 12756 6161
rect 13176 6101 13476 6161
rect 13836 6101 14256 6161
rect 12336 6041 12816 6101
rect 13116 6041 13536 6101
rect 12336 5921 12876 6041
rect 10176 5321 10656 5381
rect 10956 5321 11376 5381
rect 11676 5321 12096 5381
rect 10176 5261 10596 5321
rect 11016 5261 11316 5321
rect 11736 5261 12036 5321
rect 12336 5261 12516 5921
rect 12696 5801 12876 5921
rect 13056 5921 13596 6041
rect 13056 5501 13236 5921
rect 13416 5801 13596 5921
rect 13776 5981 14316 6101
rect 13776 5801 13956 5981
rect 14136 5801 14316 5981
rect 13776 5681 14316 5801
rect 13776 5621 14256 5681
rect 13416 5501 13596 5621
rect 13056 5381 13596 5501
rect 13776 5441 13956 5621
rect 13116 5321 13536 5381
rect 13776 5321 14316 5441
rect 13176 5261 13476 5321
rect 13836 5261 14316 5321
rect 7656 4901 7836 5261
rect 10176 4901 10356 5261
rect 7656 4841 8076 4901
rect 8376 4841 8856 4901
rect 9096 4841 9516 4901
rect 9936 4841 10356 4901
rect 7656 4781 8136 4841
rect 900 4500 2880 4680
rect 4140 4500 6120 4680
rect 7656 4661 8196 4781
rect 8376 4721 8916 4841
rect 1620 4320 3060 4500
rect 1800 4140 3060 4320
rect 3960 4320 5400 4500
rect 3960 4140 5220 4320
rect 1620 3960 2880 4140
rect 1440 3780 2880 3960
rect 4140 3960 5400 4140
rect 7656 4001 7836 4661
rect 8016 4001 8196 4661
rect 8736 4541 8916 4721
rect 8376 4361 8916 4541
rect 8376 4181 8556 4361
rect 8736 4181 8916 4361
rect 8376 4061 8916 4181
rect 8436 4001 8916 4061
rect 9096 4781 9576 4841
rect 9876 4781 10356 4841
rect 9096 4661 9636 4781
rect 9096 4001 9276 4661
rect 9456 4541 9636 4661
rect 9816 4661 10356 4781
rect 9816 4241 9996 4661
rect 10176 4241 10356 4661
rect 9816 4121 10356 4241
rect 10536 4241 10716 4901
rect 10896 4241 11076 4901
rect 11256 4241 11436 4901
rect 11616 4841 12096 4901
rect 12336 4841 12756 4901
rect 13116 4841 13536 4901
rect 11616 4721 12156 4841
rect 11976 4541 12156 4721
rect 11676 4481 12156 4541
rect 10536 4121 11436 4241
rect 11616 4361 12156 4481
rect 11616 4181 11796 4361
rect 11976 4181 12156 4361
rect 9876 4061 10356 4121
rect 10596 4061 11376 4121
rect 11616 4061 12156 4181
rect 9936 4001 10356 4061
rect 10656 4001 10896 4061
rect 11076 4001 11316 4061
rect 11676 4001 12156 4061
rect 12336 4781 12816 4841
rect 12336 4661 12876 4781
rect 12336 4001 12516 4661
rect 12696 4541 12876 4661
rect 13056 4721 13596 4841
rect 13056 4541 13236 4721
rect 13416 4541 13596 4721
rect 13056 4361 13596 4541
rect 13056 4181 13236 4361
rect 13056 4061 13596 4181
rect 13116 4001 13596 4061
rect 4140 3780 5580 3960
rect 1440 3600 2700 3780
rect 1260 3420 2700 3600
rect 4320 3660 5580 3780
rect 4320 3600 5640 3660
rect 4320 3420 5760 3600
rect 1260 3240 2520 3420
rect 4500 3240 5760 3420
rect 1260 3060 2340 3240
rect 4680 3060 5760 3240
rect 1440 2880 1980 3060
rect 5040 2880 5580 3060
<< fillblock >>
rect 376 2582 6603 8121
rect 6796 3824 14515 6352
<< end >>
