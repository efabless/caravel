magic
tech sky130A
magscale 1 2
timestamp 1666101711
<< checkpaint >>
rect 675407 99896 675887 115709
<< metal1 >>
rect 675682 113371 675734 115709
rect 675586 112665 675638 112671
rect 675586 112487 675638 112493
rect 675490 109630 675542 109636
rect 675490 109452 675542 109458
rect 675492 101631 675540 109452
rect 675588 108347 675636 112487
rect 675682 109050 675734 113199
rect 675586 108341 675638 108347
rect 675586 108163 675638 108169
rect 675490 101625 675542 101631
rect 675490 101567 675542 101573
rect 675492 100265 675540 101567
rect 675588 100462 675636 108163
rect 675586 100456 675638 100462
rect 675586 100278 675638 100284
rect 675588 100265 675636 100278
rect 675682 99896 675734 108866
<< via1 >>
rect 675682 113199 675734 113371
rect 675586 112493 675638 112665
rect 675490 109458 675542 109630
rect 675682 108866 675734 109050
rect 675586 108169 675638 108341
rect 675490 101573 675542 101625
rect 675586 100284 675638 100456
<< metal2 >>
rect 675676 113311 675682 113371
rect 675407 113255 675682 113311
rect 675676 113199 675682 113255
rect 675734 113311 675740 113371
rect 675734 113255 675887 113311
rect 675734 113199 675740 113255
rect 675407 112665 675887 112667
rect 675407 112611 675586 112665
rect 675580 112493 675586 112611
rect 675638 112611 675887 112665
rect 675638 112493 675644 112611
rect 675407 109630 675887 109631
rect 675407 109575 675490 109630
rect 675484 109458 675490 109575
rect 675542 109575 675887 109630
rect 675542 109458 675548 109575
rect 675676 108866 675682 109050
rect 675734 108866 675740 109050
rect 675407 108341 675887 108343
rect 675407 108287 675586 108341
rect 675580 108169 675586 108287
rect 675638 108287 675887 108341
rect 675638 108169 675644 108287
rect 675407 101625 675887 101627
rect 675407 101573 675490 101625
rect 675542 101573 675887 101625
rect 675407 101571 675887 101573
rect 675580 100339 675586 100456
rect 675407 100284 675586 100339
rect 675638 100339 675644 100456
rect 675638 100284 675887 100339
rect 675407 100283 675887 100284
<< properties >>
string flatten true
<< end >>
