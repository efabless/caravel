magic
tech sky130A
magscale 1 2
timestamp 1680214558
<< checkpaint >>
rect 26979 955052 29560 955590
rect 26977 954895 29568 955052
rect 26197 954869 29568 954895
rect 26197 951926 30892 954869
rect 26977 951900 30892 951926
rect 26977 951808 29568 951900
rect -1684 906704 1316 928403
rect -1726 904113 1518 906704
rect -1684 736704 1316 904113
rect -1726 734113 1518 736704
rect -1684 693704 1316 734113
rect -1726 691113 1518 693704
rect -1684 650704 1316 691113
rect -1726 648113 1518 650704
rect -1684 607704 1316 648113
rect -1726 605113 1518 607704
rect -1684 564704 1316 605113
rect -1726 562113 1518 564704
rect -1684 521704 1316 562113
rect -1726 519113 1518 521704
rect -1684 478704 1316 519113
rect -1726 476113 1518 478704
rect -1684 349704 1316 476113
rect -1726 347113 1518 349704
rect -1684 306704 1316 347113
rect -1726 304113 1518 306704
rect -1684 263704 1316 304113
rect -1726 261113 1518 263704
rect -1684 220704 1316 261113
rect -1726 218113 1518 220704
rect -1684 177704 1316 218113
rect -1726 175113 1518 177704
rect -1684 134704 1316 175113
rect -1726 132113 1518 134704
rect -1684 51887 1316 132113
rect 40340 94018 43565 970540
rect 78177 954952 80768 955052
rect 77380 954895 80768 954952
rect 129377 954916 131968 955052
rect 77380 951983 82080 954895
rect 78177 951926 82080 951983
rect 128579 954880 131968 954916
rect 180577 954895 183168 955052
rect 231777 955031 234368 955052
rect 231002 955000 234368 955031
rect 336177 955020 338768 955052
rect 231002 954983 235720 955000
rect 230894 954979 235720 954983
rect 180577 954880 184472 954895
rect 128579 951947 133274 954880
rect 78177 951808 80768 951926
rect 129377 951911 133274 951947
rect 179767 951926 184472 954880
rect 230874 951928 235720 954979
rect 336177 954964 340085 955020
rect 425177 954995 427768 955052
rect 335372 951948 340085 954964
rect 424333 954969 427768 954995
rect 179767 951911 183168 951926
rect 129377 951808 131968 951911
rect 180577 951808 183168 951911
rect 230874 951907 234368 951928
rect 230894 951815 234368 951907
rect 335372 951892 338768 951948
rect 424333 951923 429056 954969
rect 476377 954948 478968 955052
rect 575777 955042 578368 955052
rect 575777 954995 579629 955042
rect 231777 951808 234368 951815
rect 336177 951808 338768 951892
rect 425177 951897 429056 951923
rect 475540 954938 478968 954948
rect 574935 954979 579629 954995
rect 425177 951808 427768 951897
rect 475540 951876 480310 954938
rect 574935 951923 579679 954979
rect 476377 951866 480310 951876
rect 575777 951907 579679 951923
rect 476377 951808 478968 951866
rect 575777 951817 579629 951907
rect 575777 951808 578368 951817
rect 632010 929589 634850 930329
rect 631808 926997 635052 929589
rect 632010 839589 635010 926433
rect 631808 836997 635052 839589
rect 632010 750589 635010 836997
rect 631808 747997 635052 750589
rect 632010 705589 635010 747997
rect 631808 702997 635052 705589
rect 632010 660589 635010 702997
rect 631808 657997 635052 660589
rect 632010 615589 635010 657997
rect 631827 612997 635033 615589
rect 632010 570589 635010 612997
rect 631827 567997 635033 570589
rect 632010 525589 635010 567997
rect 631827 522997 635033 525589
rect 632010 348589 635010 522997
rect 631827 345997 635033 348589
rect 632010 303589 635010 345997
rect 631827 300997 635033 303589
rect 632010 258589 635010 300997
rect 631827 255997 635033 258589
rect 632010 213589 635010 255997
rect 631827 210997 635033 213589
rect 632010 168589 635010 210997
rect 631827 165997 635033 168589
rect 632010 123589 635010 165997
rect 631827 120997 635033 123589
rect 632010 78589 635010 120997
rect 674034 99654 677259 968570
rect 631827 75997 635033 78589
rect 632010 57523 635010 75997
rect -43397 -43397 -40876 -40876
<< metal2 >>
rect 27497 953270 27558 953590
rect 29498 953270 29559 953590
rect 34360 953270 34416 953750
rect 34912 953270 34968 953750
rect 35556 953270 35612 953750
rect 36200 953270 36256 953750
rect 38040 953270 38096 953750
rect 38592 953270 38648 953750
rect 39236 953270 39292 953750
rect 39880 953270 39936 953750
rect 42364 953270 42420 953750
rect 42916 953270 42972 953750
rect 43560 953270 43616 953750
rect 44204 953270 44260 953750
rect 44756 953270 44812 953750
rect 45400 953270 45456 953750
rect 46596 953270 46652 953750
rect 47240 953270 47296 953750
rect 47884 953270 47940 953750
rect 49080 953270 49136 953750
rect 78697 953270 78758 953590
rect 80698 953270 80759 953590
rect 85760 953270 85816 953750
rect 86312 953270 86368 953750
rect 86956 953270 87012 953750
rect 87600 953270 87656 953750
rect 89440 953270 89496 953750
rect 89992 953270 90048 953750
rect 90636 953270 90692 953750
rect 91280 953270 91336 953750
rect 93764 953270 93820 953750
rect 94316 953270 94372 953750
rect 94960 953270 95016 953750
rect 95604 953270 95660 953750
rect 96156 953270 96212 953750
rect 96800 953270 96856 953750
rect 97996 953270 98052 953750
rect 98640 953270 98696 953750
rect 99284 953270 99340 953750
rect 100480 953270 100536 953750
rect 129897 953270 129958 953590
rect 131898 953270 131959 953590
rect 137160 953270 137216 953750
rect 137712 953270 137768 953750
rect 138356 953270 138412 953750
rect 139000 953270 139056 953750
rect 140840 953270 140896 953750
rect 141392 953270 141448 953750
rect 142036 953270 142092 953750
rect 142680 953270 142736 953750
rect 145164 953270 145220 953750
rect 145716 953270 145772 953750
rect 146360 953270 146416 953750
rect 147004 953270 147060 953750
rect 147556 953270 147612 953750
rect 148200 953270 148256 953750
rect 149396 953270 149452 953750
rect 150040 953270 150096 953750
rect 150684 953270 150740 953750
rect 151880 953270 151936 953750
rect 181097 953270 181158 953590
rect 183098 953270 183159 953590
rect 188560 953270 188616 953750
rect 189112 953270 189168 953750
rect 189756 953270 189812 953750
rect 190400 953270 190456 953750
rect 192240 953270 192296 953750
rect 192792 953270 192848 953750
rect 193436 953270 193492 953750
rect 194080 953270 194136 953750
rect 196564 953270 196620 953750
rect 197116 953270 197172 953750
rect 197760 953270 197816 953750
rect 198404 953270 198460 953750
rect 198956 953270 199012 953750
rect 199600 953270 199656 953750
rect 200796 953270 200852 953750
rect 201440 953270 201496 953750
rect 202084 953270 202140 953750
rect 203280 953270 203336 953750
rect 232297 953270 232358 953590
rect 234298 953270 234359 953590
rect 240160 953270 240216 953750
rect 240712 953270 240768 953750
rect 241356 953270 241412 953750
rect 242000 953270 242056 953750
rect 243840 953270 243896 953750
rect 244392 953270 244448 953750
rect 245036 953270 245092 953750
rect 245680 953270 245736 953750
rect 248164 953270 248220 953750
rect 248716 953270 248772 953750
rect 249360 953270 249416 953750
rect 250004 953270 250060 953750
rect 250556 953270 250612 953750
rect 251200 953270 251256 953750
rect 252396 953270 252452 953750
rect 253040 953270 253096 953750
rect 253684 953270 253740 953750
rect 254880 953270 254936 953750
rect 336697 953270 336758 953590
rect 338698 953270 338759 953590
rect 341960 953270 342016 953750
rect 342512 953270 342568 953750
rect 343156 953270 343212 953750
rect 343800 953270 343856 953750
rect 345640 953270 345696 953750
rect 346192 953270 346248 953750
rect 346836 953270 346892 953750
rect 347480 953270 347536 953750
rect 349964 953270 350020 953750
rect 350516 953270 350572 953750
rect 351160 953270 351216 953750
rect 351804 953270 351860 953750
rect 352356 953270 352412 953750
rect 353000 953270 353056 953750
rect 354196 953270 354252 953750
rect 354840 953270 354896 953750
rect 355484 953270 355540 953750
rect 356680 953270 356736 953750
rect 425697 953270 425758 953590
rect 427698 953270 427759 953590
rect 430960 953270 431016 953750
rect 431512 953270 431568 953750
rect 432156 953270 432212 953750
rect 432800 953270 432856 953750
rect 434640 953270 434696 953750
rect 435192 953270 435248 953750
rect 435836 953270 435892 953750
rect 436480 953270 436536 953750
rect 438964 953270 439020 953750
rect 439516 953270 439572 953750
rect 440160 953270 440216 953750
rect 440804 953270 440860 953750
rect 441356 953270 441412 953750
rect 442000 953270 442056 953750
rect 443196 953270 443252 953750
rect 443840 953270 443896 953750
rect 444484 953270 444540 953750
rect 445680 953270 445736 953750
rect 476897 953270 476958 953590
rect 478898 953270 478959 953590
rect 482360 953270 482416 953750
rect 482912 953270 482968 953750
rect 483556 953270 483612 953750
rect 484200 953270 484256 953750
rect 486040 953270 486096 953750
rect 486592 953270 486648 953750
rect 487236 953270 487292 953750
rect 487880 953270 487936 953750
rect 490364 953270 490420 953750
rect 490916 953270 490972 953750
rect 491560 953270 491616 953750
rect 492204 953270 492260 953750
rect 492756 953270 492812 953750
rect 493400 953270 493456 953750
rect 494596 953270 494652 953750
rect 495240 953270 495296 953750
rect 495884 953270 495940 953750
rect 497080 953270 497136 953750
rect 576297 953270 576358 953590
rect 578298 953270 578359 953590
rect 584160 953270 584216 953750
rect 584712 953270 584768 953750
rect 585356 953270 585412 953750
rect 586000 953270 586056 953750
rect 587840 953270 587896 953750
rect 588392 953270 588448 953750
rect 589036 953270 589092 953750
rect 589680 953270 589736 953750
rect 592164 953270 592220 953750
rect 592716 953270 592772 953750
rect 593360 953270 593416 953750
rect 594004 953270 594060 953750
rect 594556 953270 594612 953750
rect 595200 953270 595256 953750
rect 596396 953270 596452 953750
rect 597040 953270 597096 953750
rect 597684 953270 597740 953750
rect 598880 953270 598936 953750
rect -274 141656 56 141663
rect -424 141600 56 141656
rect -274 141593 56 141600
rect 99571 -90 99637 56
rect 110164 -116 110220 56
rect 145190 -424 145246 56
rect 146386 -424 146442 56
rect 147030 -424 147086 56
rect 147674 -424 147730 56
rect 148870 -424 148926 56
rect 149514 -424 149570 56
rect 150066 -274 150123 56
rect 150066 -424 150122 -274
rect 150710 -424 150766 56
rect 151354 -424 151410 56
rect 151906 -424 151962 56
rect 154390 -424 154446 56
rect 155034 -424 155090 56
rect 155678 -424 155734 56
rect 156230 -424 156286 56
rect 158070 -424 158126 56
rect 158714 -424 158770 56
rect 159358 -424 159414 56
rect 159910 -424 159966 56
rect 160580 -260 160632 56
rect 163791 -259 163843 56
rect 253790 -424 253846 56
rect 254986 -424 255042 56
rect 255630 -424 255686 56
rect 256274 -424 256330 56
rect 257470 -424 257526 56
rect 258114 -424 258170 56
rect 258666 -424 258722 56
rect 259310 -424 259366 56
rect 259954 -424 260010 56
rect 260506 -424 260562 56
rect 262990 -424 263046 56
rect 263634 -424 263690 56
rect 264278 -424 264334 56
rect 264830 -424 264886 56
rect 266670 -424 266726 56
rect 267314 -424 267370 56
rect 267958 -424 268014 56
rect 268510 -424 268566 56
rect 269180 -260 269232 56
rect 273360 -260 273412 56
rect 308590 -424 308646 56
rect 309786 -424 309842 56
rect 310430 -424 310486 56
rect 311074 -424 311130 56
rect 312270 -424 312326 56
rect 312914 -424 312970 56
rect 313466 -424 313522 56
rect 314110 -424 314166 56
rect 314754 -424 314810 56
rect 315306 -424 315362 56
rect 317790 -424 317846 56
rect 318434 -424 318490 56
rect 319078 -424 319134 56
rect 319630 -424 319686 56
rect 321470 -424 321526 56
rect 322114 -424 322170 56
rect 322758 -424 322814 56
rect 323310 -424 323366 56
rect 323980 -260 324032 56
rect 328165 -282 328217 34
rect 363390 -424 363446 56
rect 364586 -424 364642 56
rect 365230 -424 365286 56
rect 365874 -424 365930 56
rect 367070 -424 367126 56
rect 367714 -424 367770 56
rect 368266 -424 368322 56
rect 368910 -424 368966 56
rect 369554 -424 369610 56
rect 370106 -424 370162 56
rect 372590 -424 372646 56
rect 373234 -424 373290 56
rect 373878 -424 373934 56
rect 374430 -424 374486 56
rect 376270 -424 376326 56
rect 376914 -424 376970 56
rect 377558 -424 377614 56
rect 378110 -424 378166 56
rect 378780 -260 378832 56
rect 382978 -260 383030 56
rect 418190 -424 418246 56
rect 419386 -424 419442 56
rect 420030 -424 420086 56
rect 420674 -424 420730 56
rect 421870 -424 421926 56
rect 422514 -424 422570 56
rect 423066 -424 423122 56
rect 423710 -424 423766 56
rect 424354 -424 424410 56
rect 424906 -424 424962 56
rect 427390 -424 427446 56
rect 428034 -424 428090 56
rect 428678 -424 428734 56
rect 429230 -424 429286 56
rect 431070 -424 431126 56
rect 431714 -424 431770 56
rect 432358 -424 432414 56
rect 432910 -424 432966 56
rect 433580 -260 433632 56
rect 437778 -260 437830 56
rect 472990 -424 473046 56
rect 474186 -424 474242 56
rect 474830 -424 474886 56
rect 475474 -424 475530 56
rect 476670 -424 476726 56
rect 477314 -424 477370 56
rect 477866 -424 477922 56
rect 478510 -424 478566 56
rect 479154 -424 479210 56
rect 479706 -424 479762 56
rect 482190 -424 482246 56
rect 482834 -424 482890 56
rect 483478 -424 483534 56
rect 484030 -424 484086 56
rect 485870 -424 485926 56
rect 486514 -424 486570 56
rect 487158 -424 487214 56
rect 487710 -424 487766 56
rect 488380 -260 488432 56
rect 492635 -260 492687 56
rect 605082 -260 605134 56
rect 605306 -260 605358 56
rect 605530 -260 605582 56
rect 605754 -260 605806 56
rect 605978 -260 606030 56
rect 606202 -260 606254 56
rect 606426 -260 606478 56
rect 606650 -260 606702 56
rect 606874 -260 606926 56
rect 607098 -260 607150 56
rect 607322 -260 607374 56
rect 607546 -260 607598 56
rect 607770 -260 607822 56
rect 607994 -260 608046 56
rect 608218 -260 608270 56
rect 608442 -260 608494 56
rect 608666 -260 608718 56
rect 608890 -260 608942 56
rect 609114 -260 609166 56
rect 609338 -260 609390 56
rect 609562 -260 609614 56
rect 609786 -260 609838 56
rect 610010 -260 610062 56
rect 610234 -260 610286 56
rect 610458 -260 610510 56
rect 610682 -260 610734 56
rect 610906 -260 610958 56
rect 611130 -260 611182 56
rect 611354 -260 611406 56
rect 611578 -260 611630 56
rect 611802 -260 611854 56
rect 612026 -260 612078 56
<< metal3 >>
rect 291362 953270 296142 953770
rect 301341 953270 306121 953770
rect 533562 953270 538342 953770
rect 543541 953270 548321 953770
rect 633270 929007 633590 929069
rect -424 927073 56 927143
rect 633270 927005 633590 927067
rect -424 925877 56 925947
rect -424 925233 56 925303
rect 633270 925103 633750 925173
rect -424 924589 56 924659
rect 633270 924551 633750 924621
rect 633270 923907 633750 923977
rect -424 923393 56 923463
rect 633270 923263 633750 923333
rect -424 922749 56 922819
rect -424 922197 56 922267
rect -424 921553 56 921623
rect 633270 921423 633750 921493
rect -424 920909 56 920979
rect 633270 920871 633750 920941
rect -424 920357 56 920427
rect 633270 920227 633750 920297
rect 633270 919583 633750 919653
rect -424 917873 56 917943
rect -424 917229 56 917299
rect 633270 917099 633750 917169
rect -424 916585 56 916655
rect 633270 916547 633750 916617
rect -424 916033 56 916103
rect 633270 915903 633750 915973
rect 633270 915259 633750 915329
rect 633270 914707 633750 914777
rect -424 914193 56 914263
rect 633270 914063 633750 914133
rect -424 913549 56 913619
rect -424 912905 56 912975
rect 633270 912867 633750 912937
rect -424 912353 56 912423
rect 633270 912223 633750 912293
rect 633270 911579 633750 911649
rect 633270 910383 633750 910453
rect -264 906644 56 906704
rect -264 904644 56 904704
rect -444 880014 56 884803
rect -444 875053 56 879715
rect 633270 875563 633770 880363
rect -444 869963 56 874763
rect 633270 870611 633770 875273
rect 633270 865523 633770 870312
rect -444 837741 56 842521
rect 633270 839007 633590 839069
rect 633270 837005 633590 837067
rect 633270 835903 633750 835973
rect 633270 835351 633750 835421
rect 633270 834707 633750 834777
rect 633270 834063 633750 834133
rect -444 827762 56 832542
rect 633270 832223 633750 832293
rect 633270 831671 633750 831741
rect 633270 831027 633750 831097
rect 633270 830383 633750 830453
rect 633270 827899 633750 827969
rect 633270 827347 633750 827417
rect 633270 826703 633750 826773
rect 633270 826059 633750 826129
rect 633270 825507 633750 825577
rect 633270 824863 633750 824933
rect 633270 823667 633750 823737
rect 633270 823023 633750 823093
rect 633270 822379 633750 822449
rect 633270 821183 633750 821253
rect -444 795541 56 800321
rect -444 785562 56 790342
rect 633270 786384 633770 791164
rect 633270 776405 633770 781185
rect -424 757273 56 757343
rect -424 756077 56 756147
rect -424 755433 56 755503
rect -424 754789 56 754859
rect -424 753593 56 753663
rect -424 752949 56 753019
rect -424 752397 56 752467
rect -424 751753 56 751823
rect -424 751109 56 751179
rect -424 750557 56 750627
rect 633270 750007 633590 750069
rect -424 748073 56 748143
rect 633270 748005 633590 748067
rect -424 747429 56 747499
rect -424 746785 56 746855
rect 633270 746703 633750 746773
rect -424 746233 56 746303
rect 633270 746151 633750 746221
rect 633270 745507 633750 745577
rect 633270 744863 633750 744933
rect -424 744393 56 744463
rect -424 743749 56 743819
rect -424 743105 56 743175
rect 633270 743023 633750 743093
rect -424 742553 56 742623
rect 633270 742471 633750 742541
rect 633270 741827 633750 741897
rect 633270 741183 633750 741253
rect 633270 738699 633750 738769
rect 633270 738147 633750 738217
rect 633270 737503 633750 737573
rect 633270 736859 633750 736929
rect -264 736644 56 736704
rect 633270 736307 633750 736377
rect 633270 735663 633750 735733
rect -264 734644 56 734704
rect 633270 734467 633750 734537
rect 633270 733823 633750 733893
rect 633270 733179 633750 733249
rect 633270 731983 633750 732053
rect -424 714073 56 714143
rect -424 712877 56 712947
rect -424 712233 56 712303
rect -424 711589 56 711659
rect -424 710393 56 710463
rect -424 709749 56 709819
rect -424 709197 56 709267
rect -424 708553 56 708623
rect -424 707909 56 707979
rect -424 707357 56 707427
rect 633270 705007 633590 705069
rect -424 704873 56 704943
rect -424 704229 56 704299
rect -424 703585 56 703655
rect -424 703033 56 703103
rect 633270 703005 633590 703067
rect 633270 701703 633750 701773
rect -424 701193 56 701263
rect 633270 701151 633750 701221
rect -424 700549 56 700619
rect 633270 700507 633750 700577
rect -424 699905 56 699975
rect 633270 699863 633750 699933
rect -424 699353 56 699423
rect 633270 698023 633750 698093
rect 633270 697471 633750 697541
rect 633270 696827 633750 696897
rect 633270 696183 633750 696253
rect -264 693644 56 693704
rect 633270 693699 633750 693769
rect 633270 693147 633750 693217
rect 633270 692503 633750 692573
rect 633270 691859 633750 691929
rect -264 691644 56 691704
rect 633270 691307 633750 691377
rect 633270 690663 633750 690733
rect 633270 689467 633750 689537
rect 633270 688823 633750 688893
rect 633270 688179 633750 688249
rect 633270 686983 633750 687053
rect -424 670873 56 670943
rect -424 669677 56 669747
rect -424 669033 56 669103
rect -424 668389 56 668459
rect -424 667193 56 667263
rect -424 666549 56 666619
rect -424 665997 56 666067
rect -424 665353 56 665423
rect -424 664709 56 664779
rect -424 664157 56 664227
rect -424 661673 56 661743
rect -424 661029 56 661099
rect -424 660385 56 660455
rect 633270 660007 633590 660069
rect -424 659833 56 659903
rect -424 657993 56 658063
rect 633270 658005 633590 658067
rect -424 657349 56 657419
rect -424 656705 56 656775
rect 633270 656703 633750 656773
rect -424 656153 56 656223
rect 633270 656151 633750 656221
rect 633270 655507 633750 655577
rect 633270 654863 633750 654933
rect 633270 653023 633750 653093
rect 633270 652471 633750 652541
rect 633270 651827 633750 651897
rect 633270 651183 633750 651253
rect -264 650644 56 650704
rect -264 648644 56 648704
rect 633270 648699 633750 648769
rect 633270 648147 633750 648217
rect 633270 647503 633750 647573
rect 633270 646859 633750 646929
rect 633270 646307 633750 646377
rect 633270 645663 633750 645733
rect 633270 644467 633750 644537
rect 633270 643823 633750 643893
rect 633270 643179 633750 643249
rect 633270 641983 633750 642053
rect -424 627673 56 627743
rect -424 626477 56 626547
rect -424 625833 56 625903
rect -424 625189 56 625259
rect -424 623993 56 624063
rect -424 623349 56 623419
rect -424 622797 56 622867
rect -424 622153 56 622223
rect -424 621509 56 621579
rect -424 620957 56 621027
rect -424 618473 56 618543
rect -424 617829 56 617899
rect -424 617185 56 617255
rect -424 616633 56 616703
rect 633270 615007 633590 615069
rect -424 614793 56 614863
rect -424 614149 56 614219
rect -424 613505 56 613575
rect -424 612953 56 613023
rect 633270 613005 633590 613067
rect 633270 611503 633750 611573
rect 633270 610951 633750 611021
rect 633270 610307 633750 610377
rect 633270 609663 633750 609733
rect 633270 607823 633750 607893
rect -264 607644 56 607704
rect 633270 607271 633750 607341
rect 633270 606627 633750 606697
rect 633270 605983 633750 606053
rect -264 605644 56 605704
rect 633270 603499 633750 603569
rect 633270 602947 633750 603017
rect 633270 602303 633750 602373
rect 633270 601659 633750 601729
rect 633270 601107 633750 601177
rect 633270 600463 633750 600533
rect 633270 599267 633750 599337
rect 633270 598623 633750 598693
rect 633270 597979 633750 598049
rect 633270 596783 633750 596853
rect -424 584473 56 584543
rect -424 583277 56 583347
rect -424 582633 56 582703
rect -424 581989 56 582059
rect -424 580793 56 580863
rect -424 580149 56 580219
rect -424 579597 56 579667
rect -424 578953 56 579023
rect -424 578309 56 578379
rect -424 577757 56 577827
rect -424 575273 56 575343
rect -424 574629 56 574699
rect -424 573985 56 574055
rect -424 573433 56 573503
rect -424 571593 56 571663
rect -424 570949 56 571019
rect -424 570305 56 570375
rect 633270 570007 633590 570069
rect -424 569753 56 569823
rect 633270 568005 633590 568067
rect 633270 566503 633750 566573
rect 633270 565951 633750 566021
rect 633270 565307 633750 565377
rect -264 564644 56 564704
rect 633270 564663 633750 564733
rect 633270 562823 633750 562893
rect -264 562644 56 562704
rect 633270 562271 633750 562341
rect 633270 561627 633750 561697
rect 633270 560983 633750 561053
rect 633270 558499 633750 558569
rect 633270 557947 633750 558017
rect 633270 557303 633750 557373
rect 633270 556659 633750 556729
rect 633270 556107 633750 556177
rect 633270 555463 633750 555533
rect 633270 554267 633750 554337
rect 633270 553623 633750 553693
rect 633270 552979 633750 553049
rect 633270 551783 633750 551853
rect -424 541273 56 541343
rect -424 540077 56 540147
rect -424 539433 56 539503
rect -424 538789 56 538859
rect -424 537593 56 537663
rect -424 536949 56 537019
rect -424 536397 56 536467
rect -424 535753 56 535823
rect -424 535109 56 535179
rect -424 534557 56 534627
rect -424 532073 56 532143
rect -424 531429 56 531499
rect -424 530785 56 530855
rect -424 530233 56 530303
rect -424 528393 56 528463
rect -424 527749 56 527819
rect -424 527105 56 527175
rect -424 526553 56 526623
rect 633270 525007 633590 525069
rect 633270 523005 633590 523067
rect -264 521644 56 521704
rect 633270 521303 633750 521373
rect 633270 520751 633750 520821
rect 633270 520107 633750 520177
rect -264 519644 56 519704
rect 633270 519463 633750 519533
rect 633270 517623 633750 517693
rect 633270 517071 633750 517141
rect 633270 516427 633750 516497
rect 633270 515783 633750 515853
rect 633270 513299 633750 513369
rect 633270 512747 633750 512817
rect 633270 512103 633750 512173
rect 633270 511459 633750 511529
rect 633270 510907 633750 510977
rect 633270 510263 633750 510333
rect 633270 509067 633750 509137
rect 633270 508423 633750 508493
rect 633270 507779 633750 507849
rect 633270 506583 633750 506653
rect -424 498073 56 498143
rect -424 496877 56 496947
rect -424 496233 56 496303
rect -424 495589 56 495659
rect -424 494393 56 494463
rect -424 493749 56 493819
rect -424 493197 56 493267
rect -424 492553 56 492623
rect -424 491909 56 491979
rect -424 491357 56 491427
rect -424 488873 56 488943
rect -424 488229 56 488299
rect -424 487585 56 487655
rect -424 487033 56 487103
rect -424 485193 56 485263
rect -424 484549 56 484619
rect -424 483905 56 483975
rect -424 483353 56 483423
rect -264 478644 56 478704
rect -264 476644 56 476704
rect 633270 471784 633770 476564
rect 633270 461805 633770 466585
rect -444 450941 56 455721
rect -444 440962 56 445742
rect 633270 427763 633770 432563
rect 633270 422812 633770 427463
rect 633270 417723 633770 422512
rect -444 408814 56 413603
rect -444 403863 56 408514
rect -444 398763 56 403563
rect 633270 383584 633770 388364
rect 633270 373605 633770 378385
rect -424 370473 56 370543
rect -424 369277 56 369347
rect -424 368633 56 368703
rect -424 367989 56 368059
rect -424 366793 56 366863
rect -424 366149 56 366219
rect -424 365597 56 365667
rect -424 364953 56 365023
rect -424 364309 56 364379
rect -424 363757 56 363827
rect -424 361273 56 361343
rect -424 360629 56 360699
rect -424 359985 56 360055
rect -424 359433 56 359503
rect -424 357593 56 357663
rect -424 356949 56 357019
rect -424 356305 56 356375
rect -424 355753 56 355823
rect -264 349644 56 349704
rect 633270 348007 633590 348069
rect -264 347644 56 347704
rect 633270 346005 633590 346067
rect 633270 344103 633750 344173
rect 633270 343551 633750 343621
rect 633270 342907 633750 342977
rect 633270 342263 633750 342333
rect 633270 340423 633750 340493
rect 633270 339871 633750 339941
rect 633270 339227 633750 339297
rect 633270 338583 633750 338653
rect 633270 336099 633750 336169
rect 633270 335547 633750 335617
rect 633270 334903 633750 334973
rect 633270 334259 633750 334329
rect 633270 333707 633750 333777
rect 633270 333063 633750 333133
rect 633270 331867 633750 331937
rect 633270 331223 633750 331293
rect 633270 330579 633750 330649
rect 633270 329383 633750 329453
rect -424 327273 56 327343
rect -424 326077 56 326147
rect -424 325433 56 325503
rect -424 324789 56 324859
rect -424 323593 56 323663
rect -424 322949 56 323019
rect -424 322397 56 322467
rect -424 321753 56 321823
rect -424 321109 56 321179
rect -424 320557 56 320627
rect -424 318073 56 318143
rect -424 317429 56 317499
rect -424 316785 56 316855
rect -424 316233 56 316303
rect -424 314393 56 314463
rect -424 313749 56 313819
rect -424 313105 56 313175
rect -424 312553 56 312623
rect -264 306644 56 306704
rect -264 304644 56 304704
rect 633270 303007 633590 303069
rect 633270 301005 633590 301067
rect 633270 298903 633750 298973
rect 633270 298351 633750 298421
rect 633270 297707 633750 297777
rect 633270 297063 633750 297133
rect 633270 295223 633750 295293
rect 633270 294671 633750 294741
rect 633270 294027 633750 294097
rect 633270 293383 633750 293453
rect 633270 290899 633750 290969
rect 633270 290347 633750 290417
rect 633270 289703 633750 289773
rect 633270 289059 633750 289129
rect 633270 288507 633750 288577
rect 633270 287863 633750 287933
rect 633270 286667 633750 286737
rect 633270 286023 633750 286093
rect 633270 285379 633750 285449
rect 633270 284183 633750 284253
rect -424 284073 56 284143
rect -424 282877 56 282947
rect -424 282233 56 282303
rect -424 281589 56 281659
rect -424 280393 56 280463
rect -424 279749 56 279819
rect -424 279197 56 279267
rect -424 278553 56 278623
rect -424 277909 56 277979
rect -424 277357 56 277427
rect -424 274873 56 274943
rect -424 274229 56 274299
rect -424 273585 56 273655
rect -424 273033 56 273103
rect -424 271193 56 271263
rect -424 270549 56 270619
rect -424 269905 56 269975
rect -424 269353 56 269423
rect -264 263644 56 263704
rect -264 261644 56 261704
rect 633270 258007 633590 258069
rect 633270 256005 633590 256067
rect 633270 253903 633750 253973
rect 633270 253351 633750 253421
rect 633270 252707 633750 252777
rect 633270 252063 633750 252133
rect 633270 250223 633750 250293
rect 633270 249671 633750 249741
rect 633270 249027 633750 249097
rect 633270 248383 633750 248453
rect 633270 245899 633750 245969
rect 633270 245347 633750 245417
rect 633270 244703 633750 244773
rect 633270 244059 633750 244129
rect 633270 243507 633750 243577
rect 633270 242863 633750 242933
rect 633270 241667 633750 241737
rect 633270 241023 633750 241093
rect -424 240873 56 240943
rect 633270 240379 633750 240449
rect -424 239677 56 239747
rect 633270 239183 633750 239253
rect -424 239033 56 239103
rect -424 238389 56 238459
rect -424 237193 56 237263
rect -424 236549 56 236619
rect -424 235997 56 236067
rect -424 235353 56 235423
rect -424 234709 56 234779
rect -424 234157 56 234227
rect -424 231673 56 231743
rect -424 231029 56 231099
rect -424 230385 56 230455
rect -424 229833 56 229903
rect -424 227993 56 228063
rect -424 227349 56 227419
rect -424 226705 56 226775
rect -424 226153 56 226223
rect -264 220644 56 220704
rect -264 218644 56 218704
rect 633270 213007 633590 213069
rect 633270 211005 633590 211067
rect 633270 208903 633750 208973
rect 633270 208351 633750 208421
rect 633270 207707 633750 207777
rect 633270 207063 633750 207133
rect 633270 205223 633750 205293
rect 633270 204671 633750 204741
rect 633270 204027 633750 204097
rect 633270 203383 633750 203453
rect 633270 200899 633750 200969
rect 633270 200347 633750 200417
rect 633270 199703 633750 199773
rect 633270 199059 633750 199129
rect 633270 198507 633750 198577
rect 633270 197863 633750 197933
rect -424 197673 56 197744
rect 633270 196667 633750 196737
rect -424 196477 56 196548
rect 633270 196023 633750 196093
rect -424 195833 56 195904
rect 633270 195379 633750 195449
rect -424 195189 56 195260
rect 633270 194183 633750 194253
rect -424 193993 56 194064
rect -424 193349 56 193420
rect -424 192797 56 192868
rect -424 192153 56 192224
rect -424 191509 56 191580
rect -424 190957 56 191028
rect -424 188473 56 188544
rect -424 187829 56 187900
rect -424 187185 56 187256
rect -424 186633 56 186704
rect -424 184793 56 184864
rect -424 184149 56 184220
rect -424 183505 56 183576
rect -424 182953 56 183024
rect -264 177644 56 177704
rect -264 175644 56 175704
rect 633270 168007 633590 168069
rect 633270 166005 633590 166067
rect 633270 163703 633750 163773
rect 633270 163151 633750 163221
rect 633270 162507 633750 162577
rect 633270 161863 633750 161933
rect 633270 160023 633750 160093
rect 633270 159471 633750 159541
rect 633270 158827 633750 158897
rect 633270 158183 633750 158253
rect 633270 155699 633750 155769
rect 633270 155147 633750 155217
rect -424 154473 56 154544
rect 633270 154503 633750 154573
rect 633270 153859 633750 153929
rect -424 153277 56 153348
rect 633270 153307 633750 153377
rect -424 152633 56 152704
rect 633270 152663 633750 152733
rect -424 151989 56 152060
rect 633270 151467 633750 151537
rect -424 150793 56 150864
rect 633270 150823 633750 150893
rect -424 150149 56 150220
rect 633270 150179 633750 150249
rect -424 149597 56 149668
rect -424 148953 56 149024
rect 633270 148983 633750 149053
rect -424 148309 56 148380
rect -424 147757 56 147828
rect -424 145273 56 145344
rect -424 144629 56 144700
rect -424 143985 56 144056
rect -424 143433 56 143504
rect -424 140949 56 141020
rect -424 140305 56 140376
rect -424 139753 56 139824
rect -264 134644 56 134704
rect -264 132644 56 132704
rect 633270 123007 633590 123069
rect 633270 121005 633590 121067
rect 633270 118703 633750 118773
rect 633270 118151 633750 118221
rect 633270 117507 633750 117577
rect 633270 116863 633750 116933
rect 633270 115023 633750 115093
rect 633270 114471 633750 114541
rect 633270 113827 633750 113897
rect 633270 113183 633750 113253
rect 633270 110699 633750 110769
rect 633270 110147 633750 110217
rect 633270 109503 633750 109573
rect 633270 108859 633750 108929
rect 633270 108307 633750 108377
rect 633270 107663 633750 107733
rect 633270 106467 633750 106537
rect 633270 105823 633750 105893
rect 633270 105179 633750 105249
rect 633270 103983 633750 104053
rect -444 78141 56 82921
rect 633270 78007 633590 78069
rect 633270 76005 633590 76067
rect 633270 73503 633750 73573
rect 633270 72951 633750 73021
rect -444 68162 56 72942
rect 633270 72307 633750 72377
rect 633270 71663 633750 71733
rect 633270 69823 633750 69893
rect 633270 69271 633750 69341
rect 633270 68627 633750 68697
rect 633270 67983 633750 68053
rect 633270 65499 633750 65569
rect 633270 64947 633750 65017
rect 633270 64303 633750 64373
rect 633270 63659 633750 63729
rect 633270 63107 633750 63177
rect 633270 62463 633750 62533
rect 633270 61267 633750 61337
rect 633270 60623 633750 60693
rect 633270 59979 633750 60049
rect 633270 58783 633750 58853
rect -283 53595 56 53665
rect -283 53372 56 53442
rect -283 53147 56 53217
rect -444 36014 56 40803
rect -444 25963 56 30763
rect 36805 -444 41585 56
rect 46784 -444 51564 57
rect 199283 -444 203912 56
rect 209163 -444 213963 56
rect 527005 -444 531785 56
rect 536984 -444 541764 56
rect 580805 -444 585585 56
rect 590784 -444 595564 56
<< comment >>
rect -400 953326 633726 953726
rect -400 0 0 953326
rect 633326 0 633726 953326
rect -400 -400 633726 0
<< labels >>
flabel metal3 -264 906644 56 906704 0 FreeSans 400 0 0 0 gpio_loopback_one[24]
port 837 nsew
flabel metal2 485870 -424 485926 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[43]
port 290 nsew
flabel metal2 s 594004 953270 594060 953750 0 FreeSans 400 90 0 0 gpio_analog_en[15]
port 450 nsew
flabel metal2 s 592716 953270 592772 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[15]
port 538 nsew
flabel metal2 s 589680 953270 589736 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[15]
port 494 nsew
flabel metal2 s 593360 953270 593416 953750 0 FreeSans 400 90 0 0 gpio_dm0[15]
port 582 nsew
flabel metal2 s 595200 953270 595256 953750 0 FreeSans 400 90 0 0 gpio_dm1[15]
port 626 nsew
flabel metal2 s 589036 953270 589092 953750 0 FreeSans 400 90 0 0 gpio_dm2[15]
port 670 nsew
flabel metal2 s 588392 953270 588448 953750 0 FreeSans 400 90 0 0 gpio_holdover[15]
port 406 nsew
flabel metal2 s 585356 953270 585412 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[15]
port 274 nsew
flabel metal2 s 592164 953270 592220 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[15]
port 230 nsew
flabel metal2 s 584712 953270 584768 953750 0 FreeSans 400 90 0 0 gpio_oeb[15]
port 186 nsew
flabel metal2 s 587840 953270 587896 953750 0 FreeSans 400 90 0 0 gpio_out[15]
port 142 nsew
flabel metal2 s 597040 953270 597096 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[15]
port 362 nsew
flabel metal2 s 586000 953270 586056 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[15]
port 318 nsew
flabel metal2 s 598880 953270 598936 953750 0 FreeSans 400 90 0 0 gpio_in[15]
port 714 nsew
flabel metal2 s 492204 953270 492260 953750 0 FreeSans 400 90 0 0 gpio_analog_en[16]
port 449 nsew
flabel metal2 s 490916 953270 490972 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[16]
port 537 nsew
flabel metal2 s 487880 953270 487936 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[16]
port 493 nsew
flabel metal2 s 491560 953270 491616 953750 0 FreeSans 400 90 0 0 gpio_dm0[16]
port 581 nsew
flabel metal2 s 493400 953270 493456 953750 0 FreeSans 400 90 0 0 gpio_dm1[16]
port 625 nsew
flabel metal2 s 487236 953270 487292 953750 0 FreeSans 400 90 0 0 gpio_dm2[16]
port 669 nsew
flabel metal2 s 486592 953270 486648 953750 0 FreeSans 400 90 0 0 gpio_holdover[16]
port 405 nsew
flabel metal2 s 483556 953270 483612 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[16]
port 273 nsew
flabel metal2 s 490364 953270 490420 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[16]
port 229 nsew
flabel metal2 s 482912 953270 482968 953750 0 FreeSans 400 90 0 0 gpio_oeb[16]
port 185 nsew
flabel metal2 s 486040 953270 486096 953750 0 FreeSans 400 90 0 0 gpio_out[16]
port 141 nsew
flabel metal2 s 495240 953270 495296 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[16]
port 361 nsew
flabel metal2 s 484200 953270 484256 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[16]
port 317 nsew
flabel metal2 s 497080 953270 497136 953750 0 FreeSans 400 90 0 0 gpio_in[16]
port 713 nsew
flabel metal2 s 597684 953270 597740 953750 0 FreeSans 400 90 0 0 gpio_loopback_one[15]
port 846 nsew
flabel metal2 s 495884 953270 495940 953750 0 FreeSans 400 90 0 0 gpio_loopback_one[16]
port 845 nsew
flabel metal2 s 442000 953270 442056 953750 0 FreeSans 400 90 0 0 gpio_dm1[17]
port 624 nsew
flabel metal2 s 435836 953270 435892 953750 0 FreeSans 400 90 0 0 gpio_dm2[17]
port 668 nsew
flabel metal2 s 435192 953270 435248 953750 0 FreeSans 400 90 0 0 gpio_holdover[17]
port 404 nsew
flabel metal2 s 432156 953270 432212 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[17]
port 272 nsew
flabel metal2 s 438964 953270 439020 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[17]
port 228 nsew
flabel metal2 s 431512 953270 431568 953750 0 FreeSans 400 90 0 0 gpio_oeb[17]
port 184 nsew
flabel metal2 s 434640 953270 434696 953750 0 FreeSans 400 90 0 0 gpio_out[17]
port 140 nsew
flabel metal2 s 443840 953270 443896 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[17]
port 360 nsew
flabel metal2 s 432800 953270 432856 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[17]
port 316 nsew
flabel metal2 s 445680 953270 445736 953750 0 FreeSans 400 90 0 0 gpio_in[17]
port 712 nsew
flabel metal2 s 351804 953270 351860 953750 0 FreeSans 400 90 0 0 gpio_analog_en[18]
port 447 nsew
flabel metal2 s 350516 953270 350572 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[18]
port 535 nsew
flabel metal2 s 347480 953270 347536 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[18]
port 491 nsew
flabel metal2 s 351160 953270 351216 953750 0 FreeSans 400 90 0 0 gpio_dm0[18]
port 579 nsew
flabel metal2 s 353000 953270 353056 953750 0 FreeSans 400 90 0 0 gpio_dm1[18]
port 623 nsew
flabel metal2 s 346836 953270 346892 953750 0 FreeSans 400 90 0 0 gpio_dm2[18]
port 667 nsew
flabel metal2 s 346192 953270 346248 953750 0 FreeSans 400 90 0 0 gpio_holdover[18]
port 403 nsew
flabel metal2 s 343156 953270 343212 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[18]
port 271 nsew
flabel metal2 s 349964 953270 350020 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[18]
port 227 nsew
flabel metal2 s 342512 953270 342568 953750 0 FreeSans 400 90 0 0 gpio_oeb[18]
port 183 nsew
flabel metal2 s 345640 953270 345696 953750 0 FreeSans 400 90 0 0 gpio_out[18]
port 139 nsew
flabel metal2 s 354840 953270 354896 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[18]
port 359 nsew
flabel metal2 s 343800 953270 343856 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[18]
port 315 nsew
flabel metal2 s 356680 953270 356736 953750 0 FreeSans 400 90 0 0 gpio_in[18]
port 711 nsew
flabel metal2 s 440804 953270 440860 953750 0 FreeSans 400 90 0 0 gpio_analog_en[17]
port 448 nsew
flabel metal2 s 439516 953270 439572 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[17]
port 536 nsew
flabel metal2 s 436480 953270 436536 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[17]
port 492 nsew
flabel metal2 s 440160 953270 440216 953750 0 FreeSans 400 90 0 0 gpio_dm0[17]
port 580 nsew
flabel metal2 s 444484 953270 444540 953750 0 FreeSans 400 90 0 0 gpio_loopback_one[17]
port 844 nsew
flabel metal2 s 355484 953270 355540 953750 0 FreeSans 400 90 0 0 gpio_loopback_one[18]
port 843 nsew
flabel metal2 s 253040 953270 253096 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[19]
port 358 nsew
flabel metal2 s 242000 953270 242056 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[19]
port 314 nsew
flabel metal2 s 254880 953270 254936 953750 0 FreeSans 400 90 0 0 gpio_in[19]
port 710 nsew
flabel metal2 s 198404 953270 198460 953750 0 FreeSans 400 90 0 0 gpio_analog_en[20]
port 445 nsew
flabel metal2 s 197116 953270 197172 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[20]
port 533 nsew
flabel metal2 s 194080 953270 194136 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[20]
port 489 nsew
flabel metal2 s 197760 953270 197816 953750 0 FreeSans 400 90 0 0 gpio_dm0[20]
port 577 nsew
flabel metal2 s 199600 953270 199656 953750 0 FreeSans 400 90 0 0 gpio_dm1[20]
port 621 nsew
flabel metal2 s 193436 953270 193492 953750 0 FreeSans 400 90 0 0 gpio_dm2[20]
port 665 nsew
flabel metal2 s 192792 953270 192848 953750 0 FreeSans 400 90 0 0 gpio_holdover[20]
port 401 nsew
flabel metal2 s 189756 953270 189812 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[20]
port 269 nsew
flabel metal2 s 196564 953270 196620 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[20]
port 225 nsew
flabel metal2 s 189112 953270 189168 953750 0 FreeSans 400 90 0 0 gpio_oeb[20]
port 181 nsew
flabel metal2 s 192240 953270 192296 953750 0 FreeSans 400 90 0 0 gpio_out[20]
port 137 nsew
flabel metal2 s 201440 953270 201496 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[20]
port 357 nsew
flabel metal2 s 190400 953270 190456 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[20]
port 313 nsew
flabel metal2 s 203280 953270 203336 953750 0 FreeSans 400 90 0 0 gpio_in[20]
port 709 nsew
flabel metal2 s 250004 953270 250060 953750 0 FreeSans 400 90 0 0 gpio_analog_en[19]
port 446 nsew
flabel metal2 s 248716 953270 248772 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[19]
port 534 nsew
flabel metal2 s 245680 953270 245736 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[19]
port 490 nsew
flabel metal2 s 249360 953270 249416 953750 0 FreeSans 400 90 0 0 gpio_dm0[19]
port 578 nsew
flabel metal2 s 251200 953270 251256 953750 0 FreeSans 400 90 0 0 gpio_dm1[19]
port 622 nsew
flabel metal2 s 245036 953270 245092 953750 0 FreeSans 400 90 0 0 gpio_dm2[19]
port 666 nsew
flabel metal2 s 244392 953270 244448 953750 0 FreeSans 400 90 0 0 gpio_holdover[19]
port 402 nsew
flabel metal2 s 241356 953270 241412 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[19]
port 270 nsew
flabel metal2 s 248164 953270 248220 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[19]
port 226 nsew
flabel metal2 s 240712 953270 240768 953750 0 FreeSans 400 90 0 0 gpio_oeb[19]
port 182 nsew
flabel metal2 s 243840 953270 243896 953750 0 FreeSans 400 90 0 0 gpio_out[19]
port 138 nsew
flabel metal2 s 253684 953270 253740 953750 0 FreeSans 400 90 0 0 gpio_loopback_one[19]
port 842 nsew
flabel metal2 s 202084 953270 202140 953750 0 FreeSans 400 90 0 0 gpio_loopback_one[20]
port 841 nsew
flabel metal2 s 151880 953270 151936 953750 0 FreeSans 400 90 0 0 gpio_in[21]
port 708 nsew
flabel metal2 s 95604 953270 95660 953750 0 FreeSans 400 90 0 0 gpio_analog_en[22]
port 443 nsew
flabel metal2 s 94316 953270 94372 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[22]
port 531 nsew
flabel metal2 s 91280 953270 91336 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[22]
port 487 nsew
flabel metal2 s 94960 953270 95016 953750 0 FreeSans 400 90 0 0 gpio_dm0[22]
port 575 nsew
flabel metal2 s 96800 953270 96856 953750 0 FreeSans 400 90 0 0 gpio_dm1[22]
port 619 nsew
flabel metal2 s 90636 953270 90692 953750 0 FreeSans 400 90 0 0 gpio_dm2[22]
port 663 nsew
flabel metal2 s 89992 953270 90048 953750 0 FreeSans 400 90 0 0 gpio_holdover[22]
port 399 nsew
flabel metal2 s 86956 953270 87012 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[22]
port 267 nsew
flabel metal2 s 93764 953270 93820 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[22]
port 223 nsew
flabel metal2 s 86312 953270 86368 953750 0 FreeSans 400 90 0 0 gpio_oeb[22]
port 179 nsew
flabel metal2 s 89440 953270 89496 953750 0 FreeSans 400 90 0 0 gpio_out[22]
port 135 nsew
flabel metal2 s 98640 953270 98696 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[22]
port 355 nsew
flabel metal2 s 87600 953270 87656 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[22]
port 311 nsew
flabel metal2 s 100480 953270 100536 953750 0 FreeSans 400 90 0 0 gpio_in[22]
port 707 nsew
flabel metal2 s 44204 953270 44260 953750 0 FreeSans 400 90 0 0 gpio_analog_en[23]
port 442 nsew
flabel metal2 s 42916 953270 42972 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[23]
port 530 nsew
flabel metal2 s 39880 953270 39936 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[23]
port 486 nsew
flabel metal2 s 43560 953270 43616 953750 0 FreeSans 400 90 0 0 gpio_dm0[23]
port 574 nsew
flabel metal2 s 45400 953270 45456 953750 0 FreeSans 400 90 0 0 gpio_dm1[23]
port 618 nsew
flabel metal2 s 39236 953270 39292 953750 0 FreeSans 400 90 0 0 gpio_dm2[23]
port 662 nsew
flabel metal2 s 38592 953270 38648 953750 0 FreeSans 400 90 0 0 gpio_holdover[23]
port 398 nsew
flabel metal2 s 35556 953270 35612 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[23]
port 266 nsew
flabel metal2 s 42364 953270 42420 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[23]
port 222 nsew
flabel metal2 s 34912 953270 34968 953750 0 FreeSans 400 90 0 0 gpio_oeb[23]
port 178 nsew
flabel metal2 s 38040 953270 38096 953750 0 FreeSans 400 90 0 0 gpio_out[23]
port 134 nsew
flabel metal2 s 47240 953270 47296 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[23]
port 354 nsew
flabel metal2 s 36200 953270 36256 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[23]
port 310 nsew
flabel metal2 s 49080 953270 49136 953750 0 FreeSans 400 90 0 0 gpio_in[23]
port 706 nsew
flabel metal2 s 147004 953270 147060 953750 0 FreeSans 400 90 0 0 gpio_analog_en[21]
port 444 nsew
flabel metal2 s 145716 953270 145772 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[21]
port 532 nsew
flabel metal2 s 142680 953270 142736 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[21]
port 488 nsew
flabel metal2 s 146360 953270 146416 953750 0 FreeSans 400 90 0 0 gpio_dm0[21]
port 576 nsew
flabel metal2 s 148200 953270 148256 953750 0 FreeSans 400 90 0 0 gpio_dm1[21]
port 620 nsew
flabel metal2 s 142036 953270 142092 953750 0 FreeSans 400 90 0 0 gpio_dm2[21]
port 664 nsew
flabel metal2 s 141392 953270 141448 953750 0 FreeSans 400 90 0 0 gpio_holdover[21]
port 400 nsew
flabel metal2 s 138356 953270 138412 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[21]
port 268 nsew
flabel metal2 s 145164 953270 145220 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[21]
port 224 nsew
flabel metal2 s 137712 953270 137768 953750 0 FreeSans 400 90 0 0 gpio_oeb[21]
port 180 nsew
flabel metal2 s 140840 953270 140896 953750 0 FreeSans 400 90 0 0 gpio_out[21]
port 136 nsew
flabel metal2 s 150040 953270 150096 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[21]
port 356 nsew
flabel metal2 s 139000 953270 139056 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[21]
port 312 nsew
flabel metal2 s 150684 953270 150740 953750 0 FreeSans 400 90 0 0 gpio_loopback_one[21]
port 840 nsew
flabel metal2 s 99284 953270 99340 953750 0 FreeSans 400 90 0 0 gpio_loopback_one[22]
port 839 nsew
flabel metal2 s 47884 953270 47940 953750 0 FreeSans 400 90 0 0 gpio_loopback_one[23]
port 838 nsew
flabel metal2 145190 -424 145246 56 0 FreeSans 400 270 0 0 gpio_in[38]
port 691 nsew
flabel metal2 146386 -424 146442 56 0 FreeSans 400 270 0 0 gpio_loopback_one[38]
port 823 nsew
flabel metal2 147030 -424 147086 56 0 FreeSans 400 270 0 0 gpio_slow_sel[38]
port 339 nsew
flabel metal2 148870 -424 148926 56 0 FreeSans 400 270 0 0 gpio_dm0[38]
port 559 nsew
flabel metal2 150710 -424 150766 56 0 FreeSans 400 270 0 0 gpio_dm1[38]
port 603 nsew
flabel metal2 151354 -424 151410 56 0 FreeSans 400 270 0 0 gpio_analog_pol[38]
port 515 nsew
flabel metal2 150066 -424 150122 56 0 FreeSans 400 270 0 0 gpio_analog_en[38]
port 427 nsew
flabel metal2 151906 -424 151962 56 0 FreeSans 400 270 0 0 gpio_inp_dis[38]
port 207 nsew
flabel metal2 154390 -424 154446 56 0 FreeSans 400 270 0 0 gpio_analog_sel[38]
port 471 nsew
flabel metal2 155034 -424 155090 56 0 FreeSans 400 270 0 0 gpio_dm2[38]
port 647 nsew
flabel metal2 155678 -424 155734 56 0 FreeSans 400 270 0 0 gpio_holdover[38]
port 383 nsew
flabel metal2 156230 -424 156286 56 0 FreeSans 400 270 0 0 gpio_out[38]
port 119 nsew
flabel metal2 158070 -424 158126 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[38]
port 295 nsew
flabel metal2 158714 -424 158770 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[38]
port 251 nsew
flabel metal2 159358 -424 159414 56 0 FreeSans 400 270 0 0 gpio_oeb[38]
port 163 nsew
flabel metal2 253790 -424 253846 56 0 FreeSans 400 270 0 0 gpio_in[39]
port 690 nsew
flabel metal2 254986 -424 255042 56 0 FreeSans 400 270 0 0 gpio_loopback_one[39]
port 822 nsew
flabel metal2 255630 -424 255686 56 0 FreeSans 400 270 0 0 gpio_slow_sel[39]
port 338 nsew
flabel metal2 257470 -424 257526 56 0 FreeSans 400 270 0 0 gpio_dm1[39]
port 602 nsew
flabel metal2 259310 -424 259366 56 0 FreeSans 400 270 0 0 gpio_dm0[39]
port 558 nsew
flabel metal2 259954 -424 260010 56 0 FreeSans 400 270 0 0 gpio_analog_pol[39]
port 514 nsew
flabel metal2 258666 -424 258722 56 0 FreeSans 400 270 0 0 gpio_analog_en[39]
port 426 nsew
flabel metal2 260506 -424 260562 56 0 FreeSans 400 270 0 0 gpio_inp_dis[39]
port 206 nsew
flabel metal2 262990 -424 263046 56 0 FreeSans 400 270 0 0 gpio_analog_sel[39]
port 470 nsew
flabel metal2 263634 -424 263690 56 0 FreeSans 400 270 0 0 gpio_dm2[39]
port 646 nsew
flabel metal2 264278 -424 264334 56 0 FreeSans 400 270 0 0 gpio_holdover[39]
port 382 nsew
flabel metal2 264830 -424 264886 56 0 FreeSans 400 270 0 0 gpio_out[39]
port 118 nsew
flabel metal2 266670 -424 266726 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[39]
port 294 nsew
flabel metal2 267314 -424 267370 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[39]
port 250 nsew
flabel metal2 267958 -424 268014 56 0 FreeSans 400 270 0 0 gpio_oeb[39]
port 162 nsew
flabel metal2 308590 -424 308646 56 0 FreeSans 400 270 0 0 gpio_in[40]
port 689 nsew
flabel metal2 309786 -424 309842 56 0 FreeSans 400 270 0 0 gpio_loopback_one[40]
port 821 nsew
flabel metal2 310430 -424 310486 56 0 FreeSans 400 270 0 0 gpio_slow_sel[40]
port 337 nsew
flabel metal2 312270 -424 312326 56 0 FreeSans 400 270 0 0 gpio_dm1[40]
port 601 nsew
flabel metal2 314110 -424 314166 56 0 FreeSans 400 270 0 0 gpio_dm0[40]
port 557 nsew
flabel metal2 314754 -424 314810 56 0 FreeSans 400 270 0 0 gpio_analog_pol[40]
port 513 nsew
flabel metal2 313466 -424 313522 56 0 FreeSans 400 270 0 0 gpio_analog_en[40]
port 425 nsew
flabel metal2 315306 -424 315362 56 0 FreeSans 400 270 0 0 gpio_inp_dis[40]
port 205 nsew
flabel metal2 317790 -424 317846 56 0 FreeSans 400 270 0 0 gpio_analog_sel[40]
port 469 nsew
flabel metal2 318434 -424 318490 56 0 FreeSans 400 270 0 0 gpio_dm2[40]
port 645 nsew
flabel metal2 319078 -424 319134 56 0 FreeSans 400 270 0 0 gpio_holdover[40]
port 381 nsew
flabel metal2 319630 -424 319686 56 0 FreeSans 400 270 0 0 gpio_out[40]
port 117 nsew
flabel metal2 321470 -424 321526 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[40]
port 293 nsew
flabel metal2 322114 -424 322170 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[40]
port 249 nsew
flabel metal2 322758 -424 322814 56 0 FreeSans 400 270 0 0 gpio_oeb[40]
port 161 nsew
flabel metal2 363390 -424 363446 56 0 FreeSans 400 270 0 0 gpio_in[41]
port 688 nsew
flabel metal2 364586 -424 364642 56 0 FreeSans 400 270 0 0 gpio_loopback_one[41]
port 820 nsew
flabel metal2 365230 -424 365286 56 0 FreeSans 400 270 0 0 gpio_slow_sel[41]
port 336 nsew
flabel metal2 367070 -424 367126 56 0 FreeSans 400 270 0 0 gpio_dm1[41]
port 600 nsew
flabel metal2 368910 -424 368966 56 0 FreeSans 400 270 0 0 gpio_dm0[41]
port 556 nsew
flabel metal2 369554 -424 369610 56 0 FreeSans 400 270 0 0 gpio_analog_pol[41]
port 512 nsew
flabel metal2 368266 -424 368322 56 0 FreeSans 400 270 0 0 gpio_analog_en[41]
port 424 nsew
flabel metal2 370106 -424 370162 56 0 FreeSans 400 270 0 0 gpio_inp_dis[41]
port 204 nsew
flabel metal2 372590 -424 372646 56 0 FreeSans 400 270 0 0 gpio_analog_sel[41]
port 468 nsew
flabel metal2 373234 -424 373290 56 0 FreeSans 400 270 0 0 gpio_dm2[41]
port 644 nsew
flabel metal2 373878 -424 373934 56 0 FreeSans 400 270 0 0 gpio_holdover[41]
port 380 nsew
flabel metal2 374430 -424 374486 56 0 FreeSans 400 270 0 0 gpio_out[41]
port 116 nsew
flabel metal2 376270 -424 376326 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[41]
port 292 nsew
flabel metal2 376914 -424 376970 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[41]
port 248 nsew
flabel metal2 377558 -424 377614 56 0 FreeSans 400 270 0 0 gpio_oeb[41]
port 160 nsew
flabel metal2 418190 -424 418246 56 0 FreeSans 400 270 0 0 gpio_in[42]
port 687 nsew
flabel metal2 419386 -424 419442 56 0 FreeSans 400 270 0 0 gpio_loopback_one[42]
port 819 nsew
flabel metal2 420030 -424 420086 56 0 FreeSans 400 270 0 0 gpio_slow_sel[42]
port 335 nsew
flabel metal2 421870 -424 421926 56 0 FreeSans 400 270 0 0 gpio_dm1[42]
port 599 nsew
flabel metal2 423710 -424 423766 56 0 FreeSans 400 270 0 0 gpio_dm0[42]
port 555 nsew
flabel metal2 424354 -424 424410 56 0 FreeSans 400 270 0 0 gpio_analog_pol[42]
port 511 nsew
flabel metal2 423066 -424 423122 56 0 FreeSans 400 270 0 0 gpio_analog_en[42]
port 423 nsew
flabel metal2 424906 -424 424962 56 0 FreeSans 400 270 0 0 gpio_inp_dis[42]
port 203 nsew
flabel metal2 427390 -424 427446 56 0 FreeSans 400 270 0 0 gpio_analog_sel[42]
port 467 nsew
flabel metal2 428034 -424 428090 56 0 FreeSans 400 270 0 0 gpio_dm2[42]
port 643 nsew
flabel metal2 428678 -424 428734 56 0 FreeSans 400 270 0 0 gpio_holdover[42]
port 379 nsew
flabel metal2 429230 -424 429286 56 0 FreeSans 400 270 0 0 gpio_out[42]
port 115 nsew
flabel metal2 431070 -424 431126 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[42]
port 291 nsew
flabel metal2 431714 -424 431770 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[42]
port 247 nsew
flabel metal2 432358 -424 432414 56 0 FreeSans 400 270 0 0 gpio_oeb[42]
port 159 nsew
flabel metal2 472990 -424 473046 56 0 FreeSans 400 270 0 0 gpio_in[43]
port 686 nsew
flabel metal2 474186 -424 474242 56 0 FreeSans 400 270 0 0 gpio_loopback_one[43]
port 818 nsew
flabel metal2 474830 -424 474886 56 0 FreeSans 400 270 0 0 gpio_slow_sel[43]
port 334 nsew
flabel metal2 476670 -424 476726 56 0 FreeSans 400 270 0 0 gpio_dm1[43]
port 598 nsew
flabel metal2 478510 -424 478566 56 0 FreeSans 400 270 0 0 gpio_dm0[43]
port 554 nsew
flabel metal2 479154 -424 479210 56 0 FreeSans 400 270 0 0 gpio_analog_pol[43]
port 510 nsew
flabel metal2 477866 -424 477922 56 0 FreeSans 400 270 0 0 gpio_analog_en[43]
port 422 nsew
flabel metal2 479706 -424 479762 56 0 FreeSans 400 270 0 0 gpio_inp_dis[43]
port 202 nsew
flabel metal2 482190 -424 482246 56 0 FreeSans 400 270 0 0 gpio_analog_sel[43]
port 466 nsew
flabel metal2 482834 -424 482890 56 0 FreeSans 400 270 0 0 gpio_dm2[43]
port 642 nsew
flabel metal2 483478 -424 483534 56 0 FreeSans 400 270 0 0 gpio_holdover[43]
port 378 nsew
flabel metal2 484030 -424 484086 56 0 FreeSans 400 270 0 0 gpio_out[43]
port 114 nsew
flabel metal2 486514 -424 486570 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[43]
port 246 nsew
flabel metal2 487158 -424 487214 56 0 FreeSans 400 270 0 0 gpio_oeb[43]
port 158 nsew
flabel metal2 s 584160 953270 584216 953750 0 FreeSans 400 90 0 0 gpio_in_h[15]
port 758 nsew
flabel metal2 s 482360 953270 482416 953750 0 FreeSans 400 90 0 0 gpio_in_h[16]
port 757 nsew
flabel metal2 s 430960 953270 431016 953750 0 FreeSans 400 90 0 0 gpio_in_h[17]
port 756 nsew
flabel metal2 s 341960 953270 342016 953750 0 FreeSans 400 90 0 0 gpio_in_h[18]
port 755 nsew
flabel metal2 s 240160 953270 240216 953750 0 FreeSans 400 90 0 0 gpio_in_h[19]
port 754 nsew
flabel metal2 s 188560 953270 188616 953750 0 FreeSans 400 90 0 0 gpio_in_h[20]
port 753 nsew
flabel metal2 s 137160 953270 137216 953750 0 FreeSans 400 90 0 0 gpio_in_h[21]
port 752 nsew
flabel metal2 s 85760 953270 85816 953750 0 FreeSans 400 90 0 0 gpio_in_h[22]
port 751 nsew
flabel metal2 s 34360 953270 34416 953750 0 FreeSans 400 90 0 0 gpio_in_h[23]
port 750 nsew
flabel metal2 s 159910 -424 159966 56 0 FreeSans 400 90 0 0 gpio_in_h[38]
port 735 nsew
flabel metal2 s 268510 -424 268566 56 0 FreeSans 400 90 0 0 gpio_in_h[39]
port 734 nsew
flabel metal2 s 323310 -424 323366 56 0 FreeSans 400 90 0 0 gpio_in_h[40]
port 733 nsew
flabel metal2 s 378110 -424 378166 56 0 FreeSans 400 90 0 0 gpio_in_h[41]
port 732 nsew
flabel metal2 s 432910 -424 432966 56 0 FreeSans 400 90 0 0 gpio_in_h[42]
port 731 nsew
flabel metal2 s 487710 -424 487766 56 0 FreeSans 400 90 0 0 gpio_in_h[43]
port 730 nsew
flabel metal2 s 596396 953270 596452 953750 0 FreeSans 400 90 0 0 analog_io[15]
port 890 nsew
flabel metal2 s 494596 953270 494652 953750 0 FreeSans 400 90 0 0 analog_io[16]
port 889 nsew
flabel metal2 s 443196 953270 443252 953750 0 FreeSans 400 90 0 0 analog_io[17]
port 888 nsew
flabel metal2 s 354196 953270 354252 953750 0 FreeSans 400 90 0 0 analog_io[18]
port 887 nsew
flabel metal2 s 252396 953270 252452 953750 0 FreeSans 400 90 0 0 analog_io[19]
port 886 nsew
flabel metal2 s 200796 953270 200852 953750 0 FreeSans 400 90 0 0 analog_io[20]
port 885 nsew
flabel metal2 s 149396 953270 149452 953750 0 FreeSans 400 90 0 0 analog_io[21]
port 884 nsew
flabel metal2 s 97996 953270 98052 953750 0 FreeSans 400 90 0 0 analog_io[22]
port 883 nsew
flabel metal2 s 46596 953270 46652 953750 0 FreeSans 400 90 0 0 analog_io[23]
port 882 nsew
flabel metal2 s 147674 -424 147730 56 0 FreeSans 400 90 0 0 analog_io[38]
port 867 nsew
flabel metal2 s 256274 -424 256330 56 0 FreeSans 400 90 0 0 analog_io[39]
port 866 nsew
flabel metal2 s 311074 -424 311130 56 0 FreeSans 400 90 0 0 analog_io[40]
port 865 nsew
flabel metal2 s 365874 -424 365930 56 0 FreeSans 400 90 0 0 analog_io[41]
port 864 nsew
flabel metal2 s 420674 -424 420730 56 0 FreeSans 400 90 0 0 analog_io[42]
port 863 nsew
flabel metal2 s 475474 -424 475530 56 0 FreeSans 400 90 0 0 analog_io[43]
port 862 nsew
flabel metal2 s 594556 953270 594612 953750 0 FreeSans 400 90 0 0 analog_noesd_io[15]
port 934 nsew
flabel metal2 s 492756 953270 492812 953750 0 FreeSans 400 90 0 0 analog_noesd_io[16]
port 933 nsew
flabel metal2 s 441356 953270 441412 953750 0 FreeSans 400 90 0 0 analog_noesd_io[17]
port 932 nsew
flabel metal2 s 352356 953270 352412 953750 0 FreeSans 400 90 0 0 analog_noesd_io[18]
port 931 nsew
flabel metal2 s 250556 953270 250612 953750 0 FreeSans 400 90 0 0 analog_noesd_io[19]
port 930 nsew
flabel metal2 s 198956 953270 199012 953750 0 FreeSans 400 90 0 0 analog_noesd_io[20]
port 929 nsew
flabel metal2 s 147556 953270 147612 953750 0 FreeSans 400 90 0 0 analog_noesd_io[21]
port 928 nsew
flabel metal2 s 96156 953270 96212 953750 0 FreeSans 400 90 0 0 analog_noesd_io[22]
port 927 nsew
flabel metal2 s 44756 953270 44812 953750 0 FreeSans 400 90 0 0 analog_noesd_io[23]
port 926 nsew
flabel metal2 s 149514 -424 149570 56 0 FreeSans 400 90 0 0 analog_noesd_io[38]
port 911 nsew
flabel metal2 s 258114 -424 258170 56 0 FreeSans 400 90 0 0 analog_noesd_io[39]
port 910 nsew
flabel metal2 s 312914 -424 312970 56 0 FreeSans 400 90 0 0 analog_noesd_io[40]
port 909 nsew
flabel metal2 s 367714 -424 367770 56 0 FreeSans 400 90 0 0 analog_noesd_io[41]
port 908 nsew
flabel metal2 s 422514 -424 422570 56 0 FreeSans 400 90 0 0 analog_noesd_io[42]
port 907 nsew
flabel metal2 s 477314 -424 477370 56 0 FreeSans 400 90 0 0 analog_noesd_io[43]
port 906 nsew
flabel metal2 s 488380 -260 488432 56 0 FreeSans 400 90 0 0 gpio_loopback_one[43]
port 818 nsew
flabel metal2 s 492635 -260 492687 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[43]
port 774 nsew
flabel metal2 s 433580 -260 433632 56 0 FreeSans 400 90 0 0 gpio_loopback_one[42]
port 819 nsew
flabel metal2 s 437778 -260 437830 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[42]
port 775 nsew
flabel metal2 s 378780 -260 378832 56 0 FreeSans 400 90 0 0 gpio_loopback_one[41]
port 820 nsew
flabel metal2 s 382978 -260 383030 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[41]
port 776 nsew
flabel metal2 s 323980 -260 324032 56 0 FreeSans 400 90 0 0 gpio_loopback_one[40]
port 821 nsew
flabel metal2 s 328165 -282 328217 34 0 FreeSans 400 90 0 0 gpio_loopback_zero[40]
port 777 nsew
flabel metal2 s 269180 -260 269232 56 0 FreeSans 400 90 0 0 gpio_loopback_one[39]
port 822 nsew
flabel metal2 s 273360 -260 273412 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[39]
port 778 nsew
flabel metal2 s 160580 -260 160632 56 0 FreeSans 400 90 0 0 gpio_loopback_one[38]
port 823 nsew
flabel metal2 s 163791 -259 163843 57 0 FreeSans 400 90 0 0 gpio_loopback_zero[38]
port 779 nsew
flabel metal2 s 110164 -116 110220 56 0 FreeSans 400 90 0 0 resetb_l
port 37 nsew
flabel metal2 s 99571 -90 99637 56 0 FreeSans 400 90 0 0 resetb_h
port 36 nsew
flabel metal2 s 605082 -260 605134 56 0 FreeSans 400 90 0 0 mask_rev[0]
port 69 nsew
flabel metal2 s 605978 -260 606030 56 0 FreeSans 400 90 0 0 mask_rev[4]
port 65 nsew
flabel metal2 s 606202 -260 606254 56 0 FreeSans 400 90 0 0 mask_rev[5]
port 64 nsew
flabel metal2 s 606426 -260 606478 56 0 FreeSans 400 90 0 0 mask_rev[6]
port 63 nsew
flabel metal2 s 606650 -260 606702 56 0 FreeSans 400 90 0 0 mask_rev[7]
port 62 nsew
flabel metal2 s 606874 -260 606926 56 0 FreeSans 400 90 0 0 mask_rev[8]
port 61 nsew
flabel metal2 s 607098 -260 607150 56 0 FreeSans 400 90 0 0 mask_rev[9]
port 60 nsew
flabel metal2 s 607322 -260 607374 56 0 FreeSans 400 90 0 0 mask_rev[10]
port 59 nsew
flabel metal2 s 607546 -260 607598 56 0 FreeSans 400 90 0 0 mask_rev[11]
port 58 nsew
flabel metal2 s 607770 -260 607822 56 0 FreeSans 400 90 0 0 mask_rev[12]
port 57 nsew
flabel metal2 s 607994 -260 608046 56 0 FreeSans 400 90 0 0 mask_rev[13]
port 56 nsew
flabel metal2 s 608218 -260 608270 56 0 FreeSans 400 90 0 0 mask_rev[14]
port 55 nsew
flabel metal2 s 608442 -260 608494 56 0 FreeSans 400 90 0 0 mask_rev[15]
port 54 nsew
flabel metal2 s 608666 -260 608718 56 0 FreeSans 400 90 0 0 mask_rev[16]
port 53 nsew
flabel metal2 s 608890 -260 608942 56 0 FreeSans 400 90 0 0 mask_rev[17]
port 52 nsew
flabel metal2 s 609114 -260 609166 56 0 FreeSans 400 90 0 0 mask_rev[18]
port 51 nsew
flabel metal2 s 609338 -260 609390 56 0 FreeSans 400 90 0 0 mask_rev[19]
port 50 nsew
flabel metal2 s 609562 -260 609614 56 0 FreeSans 400 90 0 0 mask_rev[20]
port 49 nsew
flabel metal2 s 609786 -260 609838 56 0 FreeSans 400 90 0 0 mask_rev[21]
port 48 nsew
flabel metal2 s 610010 -260 610062 56 0 FreeSans 400 90 0 0 mask_rev[22]
port 47 nsew
flabel metal2 s 610234 -260 610286 56 0 FreeSans 400 90 0 0 mask_rev[23]
port 46 nsew
flabel metal2 s 610458 -260 610510 56 0 FreeSans 400 90 0 0 mask_rev[24]
port 45 nsew
flabel metal2 s 610682 -260 610734 56 0 FreeSans 400 90 0 0 mask_rev[25]
port 44 nsew
flabel metal2 s 610906 -260 610958 56 0 FreeSans 400 90 0 0 mask_rev[26]
port 43 nsew
flabel metal2 s 611130 -260 611182 56 0 FreeSans 400 90 0 0 mask_rev[27]
port 42 nsew
flabel metal2 s 611354 -260 611406 56 0 FreeSans 400 90 0 0 mask_rev[28]
port 41 nsew
flabel metal2 s 611578 -260 611630 56 0 FreeSans 400 90 0 0 mask_rev[29]
port 40 nsew
flabel metal2 s 611802 -260 611854 56 0 FreeSans 400 90 0 0 mask_rev[30]
port 39 nsew
flabel metal2 s 612026 -260 612078 56 0 FreeSans 400 90 0 0 mask_rev[31]
port 38 nsew
flabel metal2 s 605754 -260 605806 56 0 FreeSans 400 90 0 0 mask_rev[3]
port 66 nsew
flabel metal2 s 605530 -260 605582 56 0 FreeSans 400 90 0 0 mask_rev[2]
port 67 nsew
flabel metal2 s 605306 -260 605358 56 0 FreeSans 400 90 0 0 mask_rev[1]
port 68 nsew
flabel metal2 s -424 141600 56 141656 0 FreeSans 400 0 0 0 gpio_vtrip_sel[37]
port 296 nsew
flabel metal3 633270 422812 633770 427463 0 FreeSans 3200 90 0 0 vccd1
port 28 nsew
flabel metal3 633270 427763 633770 432563 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 633270 417723 633770 422512 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 s 633270 870611 633770 875273 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 s 633270 875563 633770 880363 0 FreeSans 3200 90 0 0 vccd1
port 28 nsew
flabel metal3 s 633270 865523 633770 870312 0 FreeSans 3200 90 0 0 vccd1
port 28 nsew
flabel metal3 s 633270 786384 633770 791164 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633270 776405 633770 781185 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633270 471784 633770 476564 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633270 461805 633770 466585 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633270 383584 633770 388364 0 FreeSans 3200 90 0 0 vssa1
port 26 nsew
flabel metal3 s 633270 373605 633770 378385 0 FreeSans 3200 90 0 0 vssa1
port 26 nsew
flabel metal3 s 543541 953270 548321 953770 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 s 533562 953270 538342 953770 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 301341 953270 306121 953770 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 291362 953270 296142 953770 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 -444 875053 56 879715 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -444 880014 56 884803 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -444 869963 56 874763 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -444 837741 56 842521 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -444 827762 56 832542 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -444 795541 56 800321 0 FreeSans 3200 90 0 0 vssa2
port 27 nsew
flabel metal3 -444 785562 56 790342 0 FreeSans 3200 90 0 0 vssa2
port 27 nsew
flabel metal3 -444 450941 56 455721 0 FreeSans 3200 90 0 0 vdda2
port 25 nsew
flabel metal3 -444 440962 56 445742 0 FreeSans 3200 90 0 0 vdda2
port 25 nsew
flabel metal3 -444 403863 56 408514 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -444 408814 56 413603 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -444 398763 56 403563 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -444 78141 56 82921 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -444 68162 56 72942 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -444 36014 56 40803 0 FreeSans 3200 90 0 0 vccd
port 20 nsew
flabel metal3 -444 25963 56 30763 0 FreeSans 3200 90 0 0 vccd
port 20 nsew
flabel metal3 46784 -443 51564 57 0 FreeSans 3200 0 0 0 vssa
port 23 nsew
flabel metal3 36805 -444 41585 56 0 FreeSans 3200 0 0 0 vssa
port 23 nsew
flabel metal3 209163 -444 213963 56 0 FreeSans 3200 0 0 0 vssd
port 21 nsew
flabel metal3 199283 -444 203912 56 0 FreeSans 3200 0 0 0 vssd
port 21 nsew
flabel metal3 536984 -444 541764 56 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 527005 -444 531785 56 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 580805 -444 585585 56 0 FreeSans 3200 0 0 0 vdda
port 22 nsew
flabel metal3 590784 -444 595564 56 0 FreeSans 3200 0 0 0 vdda
port 22 nsew
flabel metal3 633270 76005 633590 76067 0 FreeSans 400 0 0 0 gpio_loopback_one[0]
port 861 nsew
flabel metal3 633270 121005 633590 121067 0 FreeSans 400 0 0 0 gpio_loopback_one[1]
port 860 nsew
flabel metal3 633270 166005 633590 166067 0 FreeSans 400 0 0 0 gpio_loopback_one[2]
port 859 nsew
flabel metal3 633270 211005 633590 211067 0 FreeSans 400 0 0 0 gpio_loopback_one[3]
port 858 nsew
flabel metal3 633270 256005 633590 256067 0 FreeSans 400 0 0 0 gpio_loopback_one[4]
port 857 nsew
flabel metal3 633270 301005 633590 301067 0 FreeSans 400 0 0 0 gpio_loopback_one[5]
port 856 nsew
flabel metal3 633270 346005 633590 346067 0 FreeSans 400 0 0 0 gpio_loopback_one[6]
port 855 nsew
flabel metal3 633270 523005 633590 523067 0 FreeSans 400 0 0 0 gpio_loopback_one[7]
port 854 nsew
flabel metal3 633270 568005 633590 568067 0 FreeSans 400 0 0 0 gpio_loopback_one[8]
port 853 nsew
flabel metal3 633270 613005 633590 613067 0 FreeSans 400 0 0 0 gpio_loopback_one[9]
port 852 nsew
flabel metal3 633270 658005 633590 658067 0 FreeSans 400 0 0 0 gpio_loopback_one[10]
port 851 nsew
flabel metal3 633270 703005 633590 703067 0 FreeSans 400 0 0 0 gpio_loopback_one[11]
port 850 nsew
flabel metal3 633270 748005 633590 748067 0 FreeSans 400 0 0 0 gpio_loopback_one[12]
port 849 nsew
flabel metal3 633270 837005 633590 837067 0 FreeSans 400 0 0 0 gpio_loopback_one[13]
port 848 nsew
flabel metal3 633270 927005 633590 927067 0 FreeSans 400 0 0 0 gpio_loopback_one[14]
port 847 nsew
flabel metal3 -264 134644 56 134704 0 FreeSans 400 0 0 0 gpio_loopback_one[37]
port 824 nsew
flabel metal3 -264 177644 56 177704 0 FreeSans 400 0 0 0 gpio_loopback_one[36]
port 825 nsew
flabel metal3 -264 220644 56 220704 0 FreeSans 400 0 0 0 gpio_loopback_one[35]
port 826 nsew
flabel metal3 -264 263644 56 263704 0 FreeSans 400 0 0 0 gpio_loopback_one[34]
port 827 nsew
flabel metal3 -264 306644 56 306704 0 FreeSans 400 0 0 0 gpio_loopback_one[33]
port 828 nsew
flabel metal3 -264 349644 56 349704 0 FreeSans 400 0 0 0 gpio_loopback_one[32]
port 829 nsew
flabel metal3 -264 478644 56 478704 0 FreeSans 400 0 0 0 gpio_loopback_one[31]
port 830 nsew
flabel metal3 -264 521644 56 521704 0 FreeSans 400 0 0 0 gpio_loopback_one[30]
port 831 nsew
flabel metal3 -264 564644 56 564704 0 FreeSans 400 0 0 0 gpio_loopback_one[29]
port 832 nsew
flabel metal3 -264 607644 56 607704 0 FreeSans 400 0 0 0 gpio_loopback_one[28]
port 833 nsew
flabel metal3 -264 650644 56 650704 0 FreeSans 400 0 0 0 gpio_loopback_one[27]
port 834 nsew
flabel metal3 -264 693644 56 693704 0 FreeSans 400 0 0 0 gpio_loopback_one[26]
port 835 nsew
flabel metal3 -264 736644 56 736704 0 FreeSans 400 0 0 0 gpio_loopback_one[25]
port 836 nsew
flabel comment s 107715 141850 108715 141850 0 FreeSans 1120000 60 0 0 example
flabel metal3 -264 261644 56 261704 0 FreeSans 400 0 0 0 gpio_loopback_zero[34]
port 783 nsew
flabel metal3 -264 218644 56 218704 0 FreeSans 400 0 0 0 gpio_loopback_zero[35]
port 782 nsew
flabel metal3 -264 175644 56 175704 0 FreeSans 400 0 0 0 gpio_loopback_zero[36]
port 781 nsew
flabel metal3 -264 132644 56 132704 0 FreeSans 400 0 0 0 gpio_loopback_zero[37]
port 780 nsew
flabel metal3 -264 304644 56 304704 0 FreeSans 400 0 0 0 gpio_loopback_zero[33]
port 784 nsew
flabel metal3 -264 347644 56 347704 0 FreeSans 400 0 0 0 gpio_loopback_zero[32]
port 785 nsew
flabel metal3 -264 476644 56 476704 0 FreeSans 400 0 0 0 gpio_loopback_zero[31]
port 786 nsew
flabel metal3 -264 519644 56 519704 0 FreeSans 400 0 0 0 gpio_loopback_zero[30]
port 787 nsew
flabel metal3 -264 562644 56 562704 0 FreeSans 400 0 0 0 gpio_loopback_zero[29]
port 788 nsew
flabel metal3 -264 605644 56 605704 0 FreeSans 400 0 0 0 gpio_loopback_zero[28]
port 789 nsew
flabel metal3 -264 648644 56 648704 0 FreeSans 400 0 0 0 gpio_loopback_zero[27]
port 790 nsew
flabel metal3 -264 691644 56 691704 0 FreeSans 400 0 0 0 gpio_loopback_zero[26]
port 791 nsew
flabel metal3 -264 734644 56 734704 0 FreeSans 400 0 0 0 gpio_loopback_zero[25]
port 792 nsew
flabel metal3 -264 904644 56 904704 0 FreeSans 400 0 0 0 gpio_loopback_zero[24]
port 793 nsew
flabel metal3 633270 929007 633590 929069 0 FreeSans 400 0 0 0 gpio_loopback_zero[14]
port 803 nsew
flabel metal3 633270 839007 633590 839069 0 FreeSans 400 0 0 0 gpio_loopback_zero[13]
port 804 nsew
flabel metal3 633270 750007 633590 750069 0 FreeSans 400 0 0 0 gpio_loopback_zero[12]
port 805 nsew
flabel metal3 633270 705007 633590 705069 0 FreeSans 400 0 0 0 gpio_loopback_zero[11]
port 806 nsew
flabel metal3 633270 660007 633590 660069 0 FreeSans 400 0 0 0 gpio_loopback_zero[10]
port 807 nsew
flabel metal3 633270 615007 633590 615069 0 FreeSans 400 0 0 0 gpio_loopback_zero[9]
port 808 nsew
flabel metal3 633270 570007 633590 570069 0 FreeSans 400 0 0 0 gpio_loopback_zero[8]
port 809 nsew
flabel metal3 633270 525007 633590 525069 0 FreeSans 400 0 0 0 gpio_loopback_zero[7]
port 810 nsew
flabel metal3 633270 348007 633590 348069 0 FreeSans 400 0 0 0 gpio_loopback_zero[6]
port 811 nsew
flabel metal3 633270 303007 633590 303069 0 FreeSans 400 0 0 0 gpio_loopback_zero[5]
port 812 nsew
flabel metal3 633270 258007 633590 258069 0 FreeSans 400 0 0 0 gpio_loopback_zero[4]
port 813 nsew
flabel metal3 633270 213007 633590 213069 0 FreeSans 400 0 0 0 gpio_loopback_zero[3]
port 814 nsew
flabel metal3 633270 168007 633590 168069 0 FreeSans 400 0 0 0 gpio_loopback_zero[2]
port 815 nsew
flabel metal3 633270 123007 633590 123069 0 FreeSans 400 0 0 0 gpio_loopback_zero[1]
port 816 nsew
flabel metal3 633270 78007 633590 78069 0 FreeSans 400 0 0 0 gpio_loopback_zero[0]
port 817 nsew
flabel metal3 s 633270 736859 633750 736929 0 FreeSans 400 0 0 0 gpio_analog_en[12]
port 453 nsew
flabel metal3 s 633270 738147 633750 738217 0 FreeSans 400 0 0 0 gpio_analog_pol[12]
port 541 nsew
flabel metal3 s 633270 741183 633750 741253 0 FreeSans 400 0 0 0 gpio_analog_sel[12]
port 497 nsew
flabel metal3 s 633270 737503 633750 737573 0 FreeSans 400 0 0 0 gpio_dm0[12]
port 585 nsew
flabel metal3 s 633270 735663 633750 735733 0 FreeSans 400 0 0 0 gpio_dm1[12]
port 629 nsew
flabel metal3 s 633270 741827 633750 741897 0 FreeSans 400 0 0 0 gpio_dm2[12]
port 673 nsew
flabel metal3 s 633270 742471 633750 742541 0 FreeSans 400 0 0 0 gpio_holdover[12]
port 409 nsew
flabel metal3 s 633270 745507 633750 745577 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[12]
port 277 nsew
flabel metal3 s 633270 738699 633750 738769 0 FreeSans 400 0 0 0 gpio_inp_dis[12]
port 233 nsew
flabel metal3 s 633270 746151 633750 746221 0 FreeSans 400 0 0 0 gpio_oeb[12]
port 189 nsew
flabel metal3 s 633270 743023 633750 743093 0 FreeSans 400 0 0 0 gpio_out[12]
port 145 nsew
flabel metal3 s 633270 733823 633750 733893 0 FreeSans 400 0 0 0 gpio_slow_sel[12]
port 365 nsew
flabel metal3 s 633270 744863 633750 744933 0 FreeSans 400 0 0 0 gpio_vtrip_sel[12]
port 321 nsew
flabel metal3 s 633270 731983 633750 732053 0 FreeSans 400 0 0 0 gpio_in[12]
port 717 nsew
flabel metal3 s 633270 826059 633750 826129 0 FreeSans 400 0 0 0 gpio_analog_en[13]
port 452 nsew
flabel metal3 s 633270 827347 633750 827417 0 FreeSans 400 0 0 0 gpio_analog_pol[13]
port 540 nsew
flabel metal3 s 633270 830383 633750 830453 0 FreeSans 400 0 0 0 gpio_analog_sel[13]
port 496 nsew
flabel metal3 s 633270 826703 633750 826773 0 FreeSans 400 0 0 0 gpio_dm0[13]
port 584 nsew
flabel metal3 s 633270 824863 633750 824933 0 FreeSans 400 0 0 0 gpio_dm1[13]
port 628 nsew
flabel metal3 s 633270 831027 633750 831097 0 FreeSans 400 0 0 0 gpio_dm2[13]
port 672 nsew
flabel metal3 s 633270 831671 633750 831741 0 FreeSans 400 0 0 0 gpio_holdover[13]
port 408 nsew
flabel metal3 s 633270 834707 633750 834777 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[13]
port 276 nsew
flabel metal3 s 633270 827899 633750 827969 0 FreeSans 400 0 0 0 gpio_inp_dis[13]
port 232 nsew
flabel metal3 s 633270 835351 633750 835421 0 FreeSans 400 0 0 0 gpio_oeb[13]
port 188 nsew
flabel metal3 s 633270 832223 633750 832293 0 FreeSans 400 0 0 0 gpio_out[13]
port 144 nsew
flabel metal3 s 633270 823023 633750 823093 0 FreeSans 400 0 0 0 gpio_slow_sel[13]
port 364 nsew
flabel metal3 s 633270 834063 633750 834133 0 FreeSans 400 0 0 0 gpio_vtrip_sel[13]
port 320 nsew
flabel metal3 s 633270 821183 633750 821253 0 FreeSans 400 0 0 0 gpio_in[13]
port 716 nsew
flabel metal3 s 633270 915259 633750 915329 0 FreeSans 400 0 0 0 gpio_analog_en[14]
port 451 nsew
flabel metal3 s 633270 916547 633750 916617 0 FreeSans 400 0 0 0 gpio_analog_pol[14]
port 539 nsew
flabel metal3 s 633270 919583 633750 919653 0 FreeSans 400 0 0 0 gpio_analog_sel[14]
port 495 nsew
flabel metal3 s 633270 915903 633750 915973 0 FreeSans 400 0 0 0 gpio_dm0[14]
port 583 nsew
flabel metal3 s 633270 914063 633750 914133 0 FreeSans 400 0 0 0 gpio_dm1[14]
port 627 nsew
flabel metal3 s 633270 920227 633750 920297 0 FreeSans 400 0 0 0 gpio_dm2[14]
port 671 nsew
flabel metal3 s 633270 920871 633750 920941 0 FreeSans 400 0 0 0 gpio_holdover[14]
port 407 nsew
flabel metal3 s 633270 923907 633750 923977 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[14]
port 275 nsew
flabel metal3 s 633270 917099 633750 917169 0 FreeSans 400 0 0 0 gpio_inp_dis[14]
port 231 nsew
flabel metal3 s 633270 924551 633750 924621 0 FreeSans 400 0 0 0 gpio_oeb[14]
port 187 nsew
flabel metal3 s 633270 921423 633750 921493 0 FreeSans 400 0 0 0 gpio_out[14]
port 143 nsew
flabel metal3 s 633270 912223 633750 912293 0 FreeSans 400 0 0 0 gpio_slow_sel[14]
port 363 nsew
flabel metal3 s 633270 923263 633750 923333 0 FreeSans 400 0 0 0 gpio_vtrip_sel[14]
port 319 nsew
flabel metal3 s 633270 910383 633750 910453 0 FreeSans 400 0 0 0 gpio_in[14]
port 715 nsew
flabel metal3 s 633270 733179 633750 733249 0 FreeSans 400 0 0 0 gpio_loopback_one[12]
port 849 nsew
flabel metal3 s 633270 822379 633750 822449 0 FreeSans 400 0 0 0 gpio_loopback_one[13]
port 848 nsew
flabel metal3 s 633270 911579 633750 911649 0 FreeSans 400 0 0 0 gpio_loopback_one[14]
port 847 nsew
flabel metal3 s 633270 697471 633750 697541 0 FreeSans 400 0 0 0 gpio_holdover[11]
port 410 nsew
flabel metal3 s 633270 700507 633750 700577 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[11]
port 278 nsew
flabel metal3 s 633270 693699 633750 693769 0 FreeSans 400 0 0 0 gpio_inp_dis[11]
port 234 nsew
flabel metal3 s 633270 701151 633750 701221 0 FreeSans 400 0 0 0 gpio_oeb[11]
port 190 nsew
flabel metal3 s 633270 698023 633750 698093 0 FreeSans 400 0 0 0 gpio_out[11]
port 146 nsew
flabel metal3 s 633270 688823 633750 688893 0 FreeSans 400 0 0 0 gpio_slow_sel[11]
port 366 nsew
flabel metal3 s 633270 699863 633750 699933 0 FreeSans 400 0 0 0 gpio_vtrip_sel[11]
port 322 nsew
flabel metal3 s 633270 686983 633750 687053 0 FreeSans 400 0 0 0 gpio_in[11]
port 718 nsew
flabel metal3 s 633270 646859 633750 646929 0 FreeSans 400 0 0 0 gpio_analog_en[10]
port 455 nsew
flabel metal3 s 633270 648147 633750 648217 0 FreeSans 400 0 0 0 gpio_analog_pol[10]
port 543 nsew
flabel metal3 s 633270 651183 633750 651253 0 FreeSans 400 0 0 0 gpio_analog_sel[10]
port 499 nsew
flabel metal3 s 633270 647503 633750 647573 0 FreeSans 400 0 0 0 gpio_dm0[10]
port 587 nsew
flabel metal3 s 633270 645663 633750 645733 0 FreeSans 400 0 0 0 gpio_dm1[10]
port 631 nsew
flabel metal3 s 633270 651827 633750 651897 0 FreeSans 400 0 0 0 gpio_dm2[10]
port 675 nsew
flabel metal3 s 633270 652471 633750 652541 0 FreeSans 400 0 0 0 gpio_holdover[10]
port 411 nsew
flabel metal3 s 633270 655507 633750 655577 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[10]
port 279 nsew
flabel metal3 s 633270 648699 633750 648769 0 FreeSans 400 0 0 0 gpio_inp_dis[10]
port 235 nsew
flabel metal3 s 633270 656151 633750 656221 0 FreeSans 400 0 0 0 gpio_oeb[10]
port 191 nsew
flabel metal3 s 633270 653023 633750 653093 0 FreeSans 400 0 0 0 gpio_out[10]
port 147 nsew
flabel metal3 s 633270 643823 633750 643893 0 FreeSans 400 0 0 0 gpio_slow_sel[10]
port 367 nsew
flabel metal3 s 633270 654863 633750 654933 0 FreeSans 400 0 0 0 gpio_vtrip_sel[10]
port 323 nsew
flabel metal3 s 633270 641983 633750 642053 0 FreeSans 400 0 0 0 gpio_in[10]
port 719 nsew
flabel metal3 s 633270 511459 633750 511529 0 FreeSans 400 0 0 0 gpio_analog_en[7]
port 458 nsew
flabel metal3 s 633270 512747 633750 512817 0 FreeSans 400 0 0 0 gpio_analog_pol[7]
port 546 nsew
flabel metal3 s 633270 515783 633750 515853 0 FreeSans 400 0 0 0 gpio_analog_sel[7]
port 502 nsew
flabel metal3 s 633270 512103 633750 512173 0 FreeSans 400 0 0 0 gpio_dm0[7]
port 590 nsew
flabel metal3 s 633270 510263 633750 510333 0 FreeSans 400 0 0 0 gpio_dm1[7]
port 634 nsew
flabel metal3 s 633270 516427 633750 516497 0 FreeSans 400 0 0 0 gpio_dm2[7]
port 678 nsew
flabel metal3 s 633270 517071 633750 517141 0 FreeSans 400 0 0 0 gpio_holdover[7]
port 414 nsew
flabel metal3 s 633270 520107 633750 520177 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[7]
port 282 nsew
flabel metal3 s 633270 513299 633750 513369 0 FreeSans 400 0 0 0 gpio_inp_dis[7]
port 238 nsew
flabel metal3 s 633270 520751 633750 520821 0 FreeSans 400 0 0 0 gpio_oeb[7]
port 194 nsew
flabel metal3 s 633270 517623 633750 517693 0 FreeSans 400 0 0 0 gpio_out[7]
port 150 nsew
flabel metal3 s 633270 508423 633750 508493 0 FreeSans 400 0 0 0 gpio_slow_sel[7]
port 370 nsew
flabel metal3 s 633270 519463 633750 519533 0 FreeSans 400 0 0 0 gpio_vtrip_sel[7]
port 326 nsew
flabel metal3 s 633270 506583 633750 506653 0 FreeSans 400 0 0 0 gpio_in[7]
port 722 nsew
flabel metal3 s 633270 556659 633750 556729 0 FreeSans 400 0 0 0 gpio_analog_en[8]
port 457 nsew
flabel metal3 s 633270 557947 633750 558017 0 FreeSans 400 0 0 0 gpio_analog_pol[8]
port 545 nsew
flabel metal3 s 633270 560983 633750 561053 0 FreeSans 400 0 0 0 gpio_analog_sel[8]
port 501 nsew
flabel metal3 s 633270 557303 633750 557373 0 FreeSans 400 0 0 0 gpio_dm0[8]
port 589 nsew
flabel metal3 s 633270 555463 633750 555533 0 FreeSans 400 0 0 0 gpio_dm1[8]
port 633 nsew
flabel metal3 s 633270 561627 633750 561697 0 FreeSans 400 0 0 0 gpio_dm2[8]
port 677 nsew
flabel metal3 s 633270 562271 633750 562341 0 FreeSans 400 0 0 0 gpio_holdover[8]
port 413 nsew
flabel metal3 s 633270 565307 633750 565377 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[8]
port 281 nsew
flabel metal3 s 633270 558499 633750 558569 0 FreeSans 400 0 0 0 gpio_inp_dis[8]
port 237 nsew
flabel metal3 s 633270 565951 633750 566021 0 FreeSans 400 0 0 0 gpio_oeb[8]
port 193 nsew
flabel metal3 s 633270 562823 633750 562893 0 FreeSans 400 0 0 0 gpio_out[8]
port 149 nsew
flabel metal3 s 633270 553623 633750 553693 0 FreeSans 400 0 0 0 gpio_slow_sel[8]
port 369 nsew
flabel metal3 s 633270 564663 633750 564733 0 FreeSans 400 0 0 0 gpio_vtrip_sel[8]
port 325 nsew
flabel metal3 s 633270 551783 633750 551853 0 FreeSans 400 0 0 0 gpio_in[8]
port 721 nsew
flabel metal3 s 633270 601659 633750 601729 0 FreeSans 400 0 0 0 gpio_analog_en[9]
port 456 nsew
flabel metal3 s 633270 602947 633750 603017 0 FreeSans 400 0 0 0 gpio_analog_pol[9]
port 544 nsew
flabel metal3 s 633270 605983 633750 606053 0 FreeSans 400 0 0 0 gpio_analog_sel[9]
port 500 nsew
flabel metal3 s 633270 602303 633750 602373 0 FreeSans 400 0 0 0 gpio_dm0[9]
port 588 nsew
flabel metal3 s 633270 600463 633750 600533 0 FreeSans 400 0 0 0 gpio_dm1[9]
port 632 nsew
flabel metal3 s 633270 606627 633750 606697 0 FreeSans 400 0 0 0 gpio_dm2[9]
port 676 nsew
flabel metal3 s 633270 607271 633750 607341 0 FreeSans 400 0 0 0 gpio_holdover[9]
port 412 nsew
flabel metal3 s 633270 610307 633750 610377 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[9]
port 280 nsew
flabel metal3 s 633270 603499 633750 603569 0 FreeSans 400 0 0 0 gpio_inp_dis[9]
port 236 nsew
flabel metal3 s 633270 610951 633750 611021 0 FreeSans 400 0 0 0 gpio_oeb[9]
port 192 nsew
flabel metal3 s 633270 607823 633750 607893 0 FreeSans 400 0 0 0 gpio_out[9]
port 148 nsew
flabel metal3 s 633270 598623 633750 598693 0 FreeSans 400 0 0 0 gpio_slow_sel[9]
port 368 nsew
flabel metal3 s 633270 609663 633750 609733 0 FreeSans 400 0 0 0 gpio_vtrip_sel[9]
port 324 nsew
flabel metal3 s 633270 596783 633750 596853 0 FreeSans 400 0 0 0 gpio_in[9]
port 720 nsew
flabel metal3 s 633270 507779 633750 507849 0 FreeSans 400 0 0 0 gpio_loopback_one[7]
port 854 nsew
flabel metal3 s 633270 552979 633750 553049 0 FreeSans 400 0 0 0 gpio_loopback_one[8]
port 853 nsew
flabel metal3 s 633270 597979 633750 598049 0 FreeSans 400 0 0 0 gpio_loopback_one[9]
port 852 nsew
flabel metal3 s 633270 643179 633750 643249 0 FreeSans 400 0 0 0 gpio_loopback_one[10]
port 851 nsew
flabel metal3 s 633270 688179 633750 688249 0 FreeSans 400 0 0 0 gpio_loopback_one[11]
port 850 nsew
flabel metal3 s 633270 691859 633750 691929 0 FreeSans 400 0 0 0 gpio_analog_en[11]
port 454 nsew
flabel metal3 s 633270 693147 633750 693217 0 FreeSans 400 0 0 0 gpio_analog_pol[11]
port 542 nsew
flabel metal3 s 633270 696183 633750 696253 0 FreeSans 400 0 0 0 gpio_analog_sel[11]
port 498 nsew
flabel metal3 s 633270 692503 633750 692573 0 FreeSans 400 0 0 0 gpio_dm0[11]
port 586 nsew
flabel metal3 s 633270 690663 633750 690733 0 FreeSans 400 0 0 0 gpio_dm1[11]
port 630 nsew
flabel metal3 s 633270 696827 633750 696897 0 FreeSans 400 0 0 0 gpio_dm2[11]
port 674 nsew
flabel metal3 s 633270 244059 633750 244129 0 FreeSans 400 0 0 0 gpio_analog_en[4]
port 461 nsew
flabel metal3 s 633270 245347 633750 245417 0 FreeSans 400 0 0 0 gpio_analog_pol[4]
port 549 nsew
flabel metal3 s 633270 248383 633750 248453 0 FreeSans 400 0 0 0 gpio_analog_sel[4]
port 505 nsew
flabel metal3 s 633270 244703 633750 244773 0 FreeSans 400 0 0 0 gpio_dm0[4]
port 593 nsew
flabel metal3 s 633270 242863 633750 242933 0 FreeSans 400 0 0 0 gpio_dm1[4]
port 637 nsew
flabel metal3 s 633270 249027 633750 249097 0 FreeSans 400 0 0 0 gpio_dm2[4]
port 681 nsew
flabel metal3 s 633270 249671 633750 249741 0 FreeSans 400 0 0 0 gpio_holdover[4]
port 417 nsew
flabel metal3 s 633270 252707 633750 252777 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[4]
port 285 nsew
flabel metal3 s 633270 245899 633750 245969 0 FreeSans 400 0 0 0 gpio_inp_dis[4]
port 241 nsew
flabel metal3 s 633270 253351 633750 253421 0 FreeSans 400 0 0 0 gpio_oeb[4]
port 197 nsew
flabel metal3 s 633270 250223 633750 250293 0 FreeSans 400 0 0 0 gpio_out[4]
port 153 nsew
flabel metal3 s 633270 241023 633750 241093 0 FreeSans 400 0 0 0 gpio_slow_sel[4]
port 373 nsew
flabel metal3 s 633270 252063 633750 252133 0 FreeSans 400 0 0 0 gpio_vtrip_sel[4]
port 329 nsew
flabel metal3 s 633270 239183 633750 239253 0 FreeSans 400 0 0 0 gpio_in[4]
port 725 nsew
flabel metal3 s 633270 289059 633750 289129 0 FreeSans 400 0 0 0 gpio_analog_en[5]
port 460 nsew
flabel metal3 s 633270 290347 633750 290417 0 FreeSans 400 0 0 0 gpio_analog_pol[5]
port 548 nsew
flabel metal3 s 633270 293383 633750 293453 0 FreeSans 400 0 0 0 gpio_analog_sel[5]
port 504 nsew
flabel metal3 s 633270 289703 633750 289773 0 FreeSans 400 0 0 0 gpio_dm0[5]
port 592 nsew
flabel metal3 s 633270 287863 633750 287933 0 FreeSans 400 0 0 0 gpio_dm1[5]
port 636 nsew
flabel metal3 s 633270 294027 633750 294097 0 FreeSans 400 0 0 0 gpio_dm2[5]
port 680 nsew
flabel metal3 s 633270 294671 633750 294741 0 FreeSans 400 0 0 0 gpio_holdover[5]
port 416 nsew
flabel metal3 s 633270 297707 633750 297777 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[5]
port 284 nsew
flabel metal3 s 633270 290899 633750 290969 0 FreeSans 400 0 0 0 gpio_inp_dis[5]
port 240 nsew
flabel metal3 s 633270 298351 633750 298421 0 FreeSans 400 0 0 0 gpio_oeb[5]
port 196 nsew
flabel metal3 s 633270 295223 633750 295293 0 FreeSans 400 0 0 0 gpio_out[5]
port 152 nsew
flabel metal3 s 633270 286023 633750 286093 0 FreeSans 400 0 0 0 gpio_slow_sel[5]
port 372 nsew
flabel metal3 s 633270 297063 633750 297133 0 FreeSans 400 0 0 0 gpio_vtrip_sel[5]
port 328 nsew
flabel metal3 s 633270 284183 633750 284253 0 FreeSans 400 0 0 0 gpio_in[5]
port 724 nsew
flabel metal3 s 633270 334259 633750 334329 0 FreeSans 400 0 0 0 gpio_analog_en[6]
port 459 nsew
flabel metal3 s 633270 240379 633750 240449 0 FreeSans 400 0 0 0 gpio_loopback_one[4]
port 857 nsew
flabel metal3 s 633270 285379 633750 285449 0 FreeSans 400 0 0 0 gpio_loopback_one[5]
port 856 nsew
flabel metal3 s 633270 330579 633750 330649 0 FreeSans 400 0 0 0 gpio_loopback_one[6]
port 855 nsew
flabel metal3 s 633270 335547 633750 335617 0 FreeSans 400 0 0 0 gpio_analog_pol[6]
port 547 nsew
flabel metal3 s 633270 338583 633750 338653 0 FreeSans 400 0 0 0 gpio_analog_sel[6]
port 503 nsew
flabel metal3 s 633270 334903 633750 334973 0 FreeSans 400 0 0 0 gpio_dm0[6]
port 591 nsew
flabel metal3 s 633270 333063 633750 333133 0 FreeSans 400 0 0 0 gpio_dm1[6]
port 635 nsew
flabel metal3 s 633270 339227 633750 339297 0 FreeSans 400 0 0 0 gpio_dm2[6]
port 679 nsew
flabel metal3 s 633270 339871 633750 339941 0 FreeSans 400 0 0 0 gpio_holdover[6]
port 415 nsew
flabel metal3 s 633270 342907 633750 342977 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[6]
port 283 nsew
flabel metal3 s 633270 336099 633750 336169 0 FreeSans 400 0 0 0 gpio_inp_dis[6]
port 239 nsew
flabel metal3 s 633270 343551 633750 343621 0 FreeSans 400 0 0 0 gpio_oeb[6]
port 195 nsew
flabel metal3 s 633270 340423 633750 340493 0 FreeSans 400 0 0 0 gpio_out[6]
port 151 nsew
flabel metal3 s 633270 331223 633750 331293 0 FreeSans 400 0 0 0 gpio_slow_sel[6]
port 371 nsew
flabel metal3 s 633270 342263 633750 342333 0 FreeSans 400 0 0 0 gpio_vtrip_sel[6]
port 327 nsew
flabel metal3 s 633270 329383 633750 329453 0 FreeSans 400 0 0 0 gpio_in[6]
port 723 nsew
flabel metal3 s 633270 108859 633750 108929 0 FreeSans 400 0 0 0 gpio_analog_en[1]
port 464 nsew
flabel metal3 s 633270 110147 633750 110217 0 FreeSans 400 0 0 0 gpio_analog_pol[1]
port 552 nsew
flabel metal3 s 633270 113183 633750 113253 0 FreeSans 400 0 0 0 gpio_analog_sel[1]
port 508 nsew
flabel metal3 s 633270 109503 633750 109573 0 FreeSans 400 0 0 0 gpio_dm0[1]
port 596 nsew
flabel metal3 s 633270 107663 633750 107733 0 FreeSans 400 0 0 0 gpio_dm1[1]
port 640 nsew
flabel metal3 s 633270 113827 633750 113897 0 FreeSans 400 0 0 0 gpio_dm2[1]
port 684 nsew
flabel metal3 s 633270 114471 633750 114541 0 FreeSans 400 0 0 0 gpio_holdover[1]
port 420 nsew
flabel metal3 s 633270 117507 633750 117577 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[1]
port 288 nsew
flabel metal3 s 633270 110699 633750 110769 0 FreeSans 400 0 0 0 gpio_inp_dis[1]
port 244 nsew
flabel metal3 s 633270 118151 633750 118221 0 FreeSans 400 0 0 0 gpio_oeb[1]
port 200 nsew
flabel metal3 s 633270 115023 633750 115093 0 FreeSans 400 0 0 0 gpio_out[1]
port 156 nsew
flabel metal3 s 633270 105823 633750 105893 0 FreeSans 400 0 0 0 gpio_slow_sel[1]
port 376 nsew
flabel metal3 s 633270 116863 633750 116933 0 FreeSans 400 0 0 0 gpio_vtrip_sel[1]
port 332 nsew
flabel metal3 s 633270 103983 633750 104053 0 FreeSans 400 0 0 0 gpio_in[1]
port 728 nsew
flabel metal3 s 633270 153859 633750 153929 0 FreeSans 400 0 0 0 gpio_analog_en[2]
port 463 nsew
flabel metal3 s 633270 155147 633750 155217 0 FreeSans 400 0 0 0 gpio_analog_pol[2]
port 551 nsew
flabel metal3 s 633270 158183 633750 158253 0 FreeSans 400 0 0 0 gpio_analog_sel[2]
port 507 nsew
flabel metal3 s 633270 154503 633750 154573 0 FreeSans 400 0 0 0 gpio_dm0[2]
port 595 nsew
flabel metal3 s 633270 152663 633750 152733 0 FreeSans 400 0 0 0 gpio_dm1[2]
port 639 nsew
flabel metal3 s 633270 158827 633750 158897 0 FreeSans 400 0 0 0 gpio_dm2[2]
port 683 nsew
flabel metal3 s 633270 159471 633750 159541 0 FreeSans 400 0 0 0 gpio_holdover[2]
port 419 nsew
flabel metal3 s 633270 162507 633750 162577 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[2]
port 287 nsew
flabel metal3 s 633270 155699 633750 155769 0 FreeSans 400 0 0 0 gpio_inp_dis[2]
port 243 nsew
flabel metal3 s 633270 163151 633750 163221 0 FreeSans 400 0 0 0 gpio_oeb[2]
port 199 nsew
flabel metal3 s 633270 160023 633750 160093 0 FreeSans 400 0 0 0 gpio_out[2]
port 155 nsew
flabel metal3 s 633270 59979 633750 60049 0 FreeSans 400 0 0 0 gpio_loopback_one[0]
port 861 nsew
flabel metal3 s 633270 105179 633750 105249 0 FreeSans 400 0 0 0 gpio_loopback_one[1]
port 860 nsew
flabel metal3 s 633270 150179 633750 150249 0 FreeSans 400 0 0 0 gpio_loopback_one[2]
port 859 nsew
flabel metal3 s 633270 195379 633750 195449 0 FreeSans 400 0 0 0 gpio_loopback_one[3]
port 858 nsew
flabel metal3 s 633270 150823 633750 150893 0 FreeSans 400 0 0 0 gpio_slow_sel[2]
port 375 nsew
flabel metal3 s 633270 161863 633750 161933 0 FreeSans 400 0 0 0 gpio_vtrip_sel[2]
port 331 nsew
flabel metal3 s 633270 148983 633750 149053 0 FreeSans 400 0 0 0 gpio_in[2]
port 727 nsew
flabel metal3 s 633270 199059 633750 199129 0 FreeSans 400 0 0 0 gpio_analog_en[3]
port 462 nsew
flabel metal3 s 633270 200347 633750 200417 0 FreeSans 400 0 0 0 gpio_analog_pol[3]
port 550 nsew
flabel metal3 s 633270 203383 633750 203453 0 FreeSans 400 0 0 0 gpio_analog_sel[3]
port 506 nsew
flabel metal3 s 633270 197863 633750 197933 0 FreeSans 400 0 0 0 gpio_dm1[3]
port 638 nsew
flabel metal3 s 633270 204027 633750 204097 0 FreeSans 400 0 0 0 gpio_dm2[3]
port 682 nsew
flabel metal3 s 633270 199703 633750 199773 0 FreeSans 400 0 0 0 gpio_dm0[3]
port 594 nsew
flabel metal3 s 633270 204671 633750 204741 0 FreeSans 400 0 0 0 gpio_holdover[3]
port 418 nsew
flabel metal3 s 633270 207707 633750 207777 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[3]
port 286 nsew
flabel metal3 s 633270 200899 633750 200969 0 FreeSans 400 0 0 0 gpio_inp_dis[3]
port 242 nsew
flabel metal3 s 633270 208351 633750 208421 0 FreeSans 400 0 0 0 gpio_oeb[3]
port 198 nsew
flabel metal3 s 633270 205223 633750 205293 0 FreeSans 400 0 0 0 gpio_out[3]
port 154 nsew
flabel metal3 s 633270 196023 633750 196093 0 FreeSans 400 0 0 0 gpio_slow_sel[3]
port 374 nsew
flabel metal3 s 633270 207063 633750 207133 0 FreeSans 400 0 0 0 gpio_vtrip_sel[3]
port 330 nsew
flabel metal3 s 633270 63659 633750 63729 0 FreeSans 400 0 0 0 gpio_analog_en[0]
port 465 nsew
flabel metal3 s 633270 64947 633750 65017 0 FreeSans 400 0 0 0 gpio_analog_pol[0]
port 553 nsew
flabel metal3 s 633270 67983 633750 68053 0 FreeSans 400 0 0 0 gpio_analog_sel[0]
port 509 nsew
flabel metal3 s 633270 64303 633750 64373 0 FreeSans 400 0 0 0 gpio_dm0[0]
port 597 nsew
flabel metal3 s 633270 62463 633750 62533 0 FreeSans 400 0 0 0 gpio_dm1[0]
port 641 nsew
flabel metal3 s 633270 68627 633750 68697 0 FreeSans 400 0 0 0 gpio_dm2[0]
port 685 nsew
flabel metal3 s 633270 69271 633750 69341 0 FreeSans 400 0 0 0 gpio_holdover[0]
port 421 nsew
flabel metal3 s 633270 72307 633750 72377 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[0]
port 289 nsew
flabel metal3 s 633270 65499 633750 65569 0 FreeSans 400 0 0 0 gpio_inp_dis[0]
port 245 nsew
flabel metal3 s 633270 72951 633750 73021 0 FreeSans 400 0 0 0 gpio_oeb[0]
port 201 nsew
flabel metal3 s 633270 69823 633750 69893 0 FreeSans 400 0 0 0 gpio_out[0]
port 157 nsew
flabel metal3 s 633270 60623 633750 60693 0 FreeSans 400 0 0 0 gpio_slow_sel[0]
port 377 nsew
flabel metal3 s 633270 71663 633750 71733 0 FreeSans 400 0 0 0 gpio_vtrip_sel[0]
port 333 nsew
flabel metal3 s 633270 58783 633750 58853 0 FreeSans 400 0 0 0 gpio_in[0]
port 729 nsew
flabel metal3 s 633270 194183 633750 194253 0 FreeSans 400 0 0 0 gpio_in[3]
port 726 nsew
flabel metal3 633270 61267 633750 61337 0 FreeSans 400 0 0 0 analog_io[0]
port 905 nsew
flabel metal3 633270 63107 633750 63177 0 FreeSans 400 0 0 0 analog_noesd_io[0]
port 949 nsew
flabel metal3 633270 108307 633750 108377 0 FreeSans 400 0 0 0 analog_noesd_io[1]
port 948 nsew
flabel metal3 633270 106467 633750 106537 0 FreeSans 400 0 0 0 analog_io[1]
port 904 nsew
flabel metal3 633270 73503 633750 73573 0 FreeSans 400 0 0 0 gpio_in_h[0]
port 773 nsew
flabel metal3 633270 118703 633750 118773 0 FreeSans 400 0 0 0 gpio_in_h[1]
port 772 nsew
flabel metal3 633270 151467 633750 151537 0 FreeSans 400 0 0 0 analog_io[2]
port 903 nsew
flabel metal3 633270 153307 633750 153377 0 FreeSans 400 0 0 0 analog_noesd_io[2]
port 947 nsew
flabel metal3 633270 163703 633750 163773 0 FreeSans 400 0 0 0 gpio_in_h[2]
port 771 nsew
flabel metal3 633270 196667 633750 196737 0 FreeSans 400 0 0 0 analog_io[3]
port 902 nsew
flabel metal3 633270 198507 633750 198577 0 FreeSans 400 0 0 0 analog_noesd_io[3]
port 946 nsew
flabel metal3 633270 208903 633750 208973 0 FreeSans 400 0 0 0 gpio_in_h[3]
port 770 nsew
flabel metal3 633270 241667 633750 241737 0 FreeSans 400 0 0 0 analog_io[4]
port 901 nsew
flabel metal3 633270 243507 633750 243577 0 FreeSans 400 0 0 0 analog_noesd_io[4]
port 945 nsew
flabel metal3 633270 253903 633750 253973 0 FreeSans 400 0 0 0 gpio_in_h[4]
port 769 nsew
flabel metal3 633270 286667 633750 286737 0 FreeSans 400 0 0 0 analog_io[5]
port 900 nsew
flabel metal3 633270 288507 633750 288577 0 FreeSans 400 0 0 0 analog_noesd_io[5]
port 944 nsew
flabel metal3 633270 298903 633750 298973 0 FreeSans 400 0 0 0 gpio_in_h[5]
port 768 nsew
flabel metal3 633270 331867 633750 331937 0 FreeSans 400 0 0 0 analog_io[6]
port 899 nsew
flabel metal3 633270 333707 633750 333777 0 FreeSans 400 0 0 0 analog_noesd_io[6]
port 943 nsew
flabel metal3 633270 344103 633750 344173 0 FreeSans 400 0 0 0 gpio_in_h[6]
port 767 nsew
flabel metal3 s 633270 509067 633750 509137 0 FreeSans 400 0 0 0 analog_io[7]
port 898 nsew
flabel metal3 s 633270 510907 633750 510977 0 FreeSans 400 0 0 0 analog_noesd_io[7]
port 942 nsew
flabel metal3 s 633270 521303 633750 521373 0 FreeSans 400 0 0 0 gpio_in_h[7]
port 766 nsew
flabel metal3 s 633270 554267 633750 554337 0 FreeSans 400 0 0 0 analog_io[8]
port 897 nsew
flabel metal3 s 633270 556107 633750 556177 0 FreeSans 400 0 0 0 analog_noesd_io[8]
port 941 nsew
flabel metal3 s 633270 566503 633750 566573 0 FreeSans 400 0 0 0 gpio_in_h[8]
port 765 nsew
flabel metal3 s 633270 599267 633750 599337 0 FreeSans 400 0 0 0 analog_io[9]
port 896 nsew
flabel metal3 s 633270 601107 633750 601177 0 FreeSans 400 0 0 0 analog_noesd_io[9]
port 940 nsew
flabel metal3 s 633270 611503 633750 611573 0 FreeSans 400 0 0 0 gpio_in_h[9]
port 764 nsew
flabel metal3 s 633270 644467 633750 644537 0 FreeSans 400 0 0 0 analog_io[10]
port 895 nsew
flabel metal3 s 633270 646307 633750 646377 0 FreeSans 400 0 0 0 analog_noesd_io[10]
port 939 nsew
flabel metal3 s 633270 656703 633750 656773 0 FreeSans 400 0 0 0 gpio_in_h[10]
port 763 nsew
flabel metal3 s 633270 689467 633750 689537 0 FreeSans 400 0 0 0 analog_io[11]
port 894 nsew
flabel metal3 s 633270 691307 633750 691377 0 FreeSans 400 0 0 0 analog_noesd_io[11]
port 938 nsew
flabel metal3 s 633270 701703 633750 701773 0 FreeSans 400 0 0 0 gpio_in_h[11]
port 762 nsew
flabel metal3 s 633270 746703 633750 746773 0 FreeSans 400 0 0 0 gpio_in_h[12]
port 761 nsew
flabel metal3 s 633270 835903 633750 835973 0 FreeSans 400 0 0 0 gpio_in_h[13]
port 760 nsew
flabel metal3 s 633270 925103 633750 925173 0 FreeSans 400 0 0 0 gpio_in_h[14]
port 759 nsew
flabel metal3 s 633270 734467 633750 734537 0 FreeSans 400 0 0 0 analog_io[12]
port 893 nsew
flabel metal3 s 633270 823667 633750 823737 0 FreeSans 400 0 0 0 analog_io[13]
port 892 nsew
flabel metal3 s 633270 912867 633750 912937 0 FreeSans 400 0 0 0 analog_io[14]
port 891 nsew
flabel metal3 s 633270 736307 633750 736377 0 FreeSans 400 0 0 0 analog_noesd_io[12]
port 937 nsew
flabel metal3 s 633270 825507 633750 825577 0 FreeSans 400 0 0 0 analog_noesd_io[13]
port 936 nsew
flabel metal3 s 633270 914707 633750 914777 0 FreeSans 400 0 0 0 analog_noesd_io[14]
port 935 nsew
flabel metal3 s -424 925877 56 925947 0 FreeSans 400 0 0 0 gpio_loopback_one[24]
port 837 nsew
flabel metal3 s -424 922197 56 922267 0 FreeSans 400 0 0 0 gpio_analog_en[24]
port 441 nsew
flabel metal3 s -424 920909 56 920979 0 FreeSans 400 0 0 0 gpio_analog_pol[24]
port 529 nsew
flabel metal3 s -424 917873 56 917943 0 FreeSans 400 0 0 0 gpio_analog_sel[24]
port 485 nsew
flabel metal3 s -424 921553 56 921623 0 FreeSans 400 0 0 0 gpio_dm0[24]
port 573 nsew
flabel metal3 s -424 923393 56 923463 0 FreeSans 400 0 0 0 gpio_dm1[24]
port 617 nsew
flabel metal3 s -424 917229 56 917299 0 FreeSans 400 0 0 0 gpio_dm2[24]
port 661 nsew
flabel metal3 s -424 916585 56 916655 0 FreeSans 400 0 0 0 gpio_holdover[24]
port 397 nsew
flabel metal3 s -424 913549 56 913619 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[24]
port 265 nsew
flabel metal3 s -424 920357 56 920427 0 FreeSans 400 0 0 0 gpio_inp_dis[24]
port 221 nsew
flabel metal3 s -424 912905 56 912975 0 FreeSans 400 0 0 0 gpio_oeb[24]
port 177 nsew
flabel metal3 s -424 916033 56 916103 0 FreeSans 400 0 0 0 gpio_out[24]
port 133 nsew
flabel metal3 s -424 925233 56 925303 0 FreeSans 400 0 0 0 gpio_slow_sel[24]
port 353 nsew
flabel metal3 s -424 914193 56 914263 0 FreeSans 400 0 0 0 gpio_vtrip_sel[24]
port 309 nsew
flabel metal3 s -424 927073 56 927143 0 FreeSans 400 0 0 0 gpio_in[24]
port 705 nsew
flabel metal3 s -424 912353 56 912423 0 FreeSans 400 0 0 0 gpio_in_h[24]
port 749 nsew
flabel metal3 s -424 924589 56 924659 0 FreeSans 400 0 0 0 analog_io[24]
port 881 nsew
flabel metal3 s -424 922749 56 922819 0 FreeSans 400 0 0 0 analog_noesd_io[24]
port 925 nsew
flabel metal3 -283 53372 56 53442 0 FreeSans 400 0 0 0 por_l
port 35 nsew
flabel metal3 -283 53595 56 53665 0 FreeSans 400 0 0 0 porb_l
port 34 nsew
flabel metal3 -283 53147 56 53217 0 FreeSans 400 0 0 0 porb_h
port 33 nsew
flabel metal3 s -424 752397 56 752467 0 FreeSans 400 0 0 0 gpio_analog_en[25]
port 440 nsew
flabel metal3 s -424 751109 56 751179 0 FreeSans 400 0 0 0 gpio_analog_pol[25]
port 528 nsew
flabel metal3 s -424 748073 56 748143 0 FreeSans 400 0 0 0 gpio_analog_sel[25]
port 484 nsew
flabel metal3 s -424 751753 56 751823 0 FreeSans 400 0 0 0 gpio_dm0[25]
port 572 nsew
flabel metal3 s -424 753593 56 753663 0 FreeSans 400 0 0 0 gpio_dm1[25]
port 616 nsew
flabel metal3 s -424 747429 56 747499 0 FreeSans 400 0 0 0 gpio_dm2[25]
port 660 nsew
flabel metal3 s -424 746785 56 746855 0 FreeSans 400 0 0 0 gpio_holdover[25]
port 396 nsew
flabel metal3 s -424 743749 56 743819 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[25]
port 264 nsew
flabel metal3 s -424 750557 56 750627 0 FreeSans 400 0 0 0 gpio_inp_dis[25]
port 220 nsew
flabel metal3 s -424 743105 56 743175 0 FreeSans 400 0 0 0 gpio_oeb[25]
port 176 nsew
flabel metal3 s -424 746233 56 746303 0 FreeSans 400 0 0 0 gpio_out[25]
port 132 nsew
flabel metal3 s -424 755433 56 755503 0 FreeSans 400 0 0 0 gpio_slow_sel[25]
port 352 nsew
flabel metal3 s -424 757273 56 757343 0 FreeSans 400 0 0 0 gpio_in[25]
port 704 nsew
flabel metal3 s -424 756077 56 756147 0 FreeSans 400 0 0 0 gpio_loopback_one[25]
port 836 nsew
flabel metal3 s -424 535753 56 535823 0 FreeSans 400 0 0 0 gpio_dm0[30]
port 567 nsew
flabel metal3 s -424 537593 56 537663 0 FreeSans 400 0 0 0 gpio_dm1[30]
port 611 nsew
flabel metal3 s -424 531429 56 531499 0 FreeSans 400 0 0 0 gpio_dm2[30]
port 655 nsew
flabel metal3 s -424 530785 56 530855 0 FreeSans 400 0 0 0 gpio_holdover[30]
port 391 nsew
flabel metal3 s -424 527749 56 527819 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[30]
port 259 nsew
flabel metal3 s -424 534557 56 534627 0 FreeSans 400 0 0 0 gpio_inp_dis[30]
port 215 nsew
flabel metal3 s -424 527105 56 527175 0 FreeSans 400 0 0 0 gpio_oeb[30]
port 171 nsew
flabel metal3 s -424 530233 56 530303 0 FreeSans 400 0 0 0 gpio_out[30]
port 127 nsew
flabel metal3 s -424 539433 56 539503 0 FreeSans 400 0 0 0 gpio_slow_sel[30]
port 347 nsew
flabel metal3 s -424 528393 56 528463 0 FreeSans 400 0 0 0 gpio_vtrip_sel[30]
port 303 nsew
flabel metal3 s -424 541273 56 541343 0 FreeSans 400 0 0 0 gpio_in[30]
port 699 nsew
flabel metal3 s -424 493197 56 493267 0 FreeSans 400 0 0 0 gpio_analog_en[31]
port 434 nsew
flabel metal3 s -424 491909 56 491979 0 FreeSans 400 0 0 0 gpio_analog_pol[31]
port 522 nsew
flabel metal3 s -424 488873 56 488943 0 FreeSans 400 0 0 0 gpio_analog_sel[31]
port 478 nsew
flabel metal3 s -424 492553 56 492623 0 FreeSans 400 0 0 0 gpio_dm0[31]
port 566 nsew
flabel metal3 s -424 494393 56 494463 0 FreeSans 400 0 0 0 gpio_dm1[31]
port 610 nsew
flabel metal3 s -424 488229 56 488299 0 FreeSans 400 0 0 0 gpio_dm2[31]
port 654 nsew
flabel metal3 s -424 487585 56 487655 0 FreeSans 400 0 0 0 gpio_holdover[31]
port 390 nsew
flabel metal3 s -424 484549 56 484619 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[31]
port 258 nsew
flabel metal3 s -424 491357 56 491427 0 FreeSans 400 0 0 0 gpio_inp_dis[31]
port 214 nsew
flabel metal3 s -424 483905 56 483975 0 FreeSans 400 0 0 0 gpio_oeb[31]
port 170 nsew
flabel metal3 s -424 487033 56 487103 0 FreeSans 400 0 0 0 gpio_out[31]
port 126 nsew
flabel metal3 s -424 496233 56 496303 0 FreeSans 400 0 0 0 gpio_slow_sel[31]
port 346 nsew
flabel metal3 s -424 485193 56 485263 0 FreeSans 400 0 0 0 gpio_vtrip_sel[31]
port 302 nsew
flabel metal3 s -424 498073 56 498143 0 FreeSans 400 0 0 0 gpio_in[31]
port 698 nsew
flabel metal3 s -424 709197 56 709267 0 FreeSans 400 0 0 0 gpio_analog_en[26]
port 439 nsew
flabel metal3 s -424 707909 56 707979 0 FreeSans 400 0 0 0 gpio_analog_pol[26]
port 527 nsew
flabel metal3 s -424 704873 56 704943 0 FreeSans 400 0 0 0 gpio_analog_sel[26]
port 483 nsew
flabel metal3 s -424 708553 56 708623 0 FreeSans 400 0 0 0 gpio_dm0[26]
port 571 nsew
flabel metal3 s -424 710393 56 710463 0 FreeSans 400 0 0 0 gpio_dm1[26]
port 615 nsew
flabel metal3 s -424 704229 56 704299 0 FreeSans 400 0 0 0 gpio_dm2[26]
port 659 nsew
flabel metal3 s -424 703585 56 703655 0 FreeSans 400 0 0 0 gpio_holdover[26]
port 395 nsew
flabel metal3 s -424 700549 56 700619 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[26]
port 263 nsew
flabel metal3 s -424 707357 56 707427 0 FreeSans 400 0 0 0 gpio_inp_dis[26]
port 219 nsew
flabel metal3 s -424 699905 56 699975 0 FreeSans 400 0 0 0 gpio_oeb[26]
port 175 nsew
flabel metal3 s -424 703033 56 703103 0 FreeSans 400 0 0 0 gpio_out[26]
port 131 nsew
flabel metal3 s -424 712233 56 712303 0 FreeSans 400 0 0 0 gpio_slow_sel[26]
port 351 nsew
flabel metal3 s -424 701193 56 701263 0 FreeSans 400 0 0 0 gpio_vtrip_sel[26]
port 307 nsew
flabel metal3 s -424 714073 56 714143 0 FreeSans 400 0 0 0 gpio_in[26]
port 703 nsew
flabel metal3 s -424 665997 56 666067 0 FreeSans 400 0 0 0 gpio_analog_en[27]
port 438 nsew
flabel metal3 s -424 664709 56 664779 0 FreeSans 400 0 0 0 gpio_analog_pol[27]
port 526 nsew
flabel metal3 s -424 661673 56 661743 0 FreeSans 400 0 0 0 gpio_analog_sel[27]
port 482 nsew
flabel metal3 s -424 665353 56 665423 0 FreeSans 400 0 0 0 gpio_dm0[27]
port 570 nsew
flabel metal3 s -424 667193 56 667263 0 FreeSans 400 0 0 0 gpio_dm1[27]
port 614 nsew
flabel metal3 s -424 661029 56 661099 0 FreeSans 400 0 0 0 gpio_dm2[27]
port 658 nsew
flabel metal3 s -424 660385 56 660455 0 FreeSans 400 0 0 0 gpio_holdover[27]
port 394 nsew
flabel metal3 s -424 657349 56 657419 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[27]
port 262 nsew
flabel metal3 s -424 664157 56 664227 0 FreeSans 400 0 0 0 gpio_inp_dis[27]
port 218 nsew
flabel metal3 s -424 656705 56 656775 0 FreeSans 400 0 0 0 gpio_oeb[27]
port 174 nsew
flabel metal3 s -424 659833 56 659903 0 FreeSans 400 0 0 0 gpio_out[27]
port 130 nsew
flabel metal3 s -424 669033 56 669103 0 FreeSans 400 0 0 0 gpio_slow_sel[27]
port 350 nsew
flabel metal3 s -424 657993 56 658063 0 FreeSans 400 0 0 0 gpio_vtrip_sel[27]
port 306 nsew
flabel metal3 s -424 670873 56 670943 0 FreeSans 400 0 0 0 gpio_in[27]
port 702 nsew
flabel metal3 s -424 622797 56 622867 0 FreeSans 400 0 0 0 gpio_analog_en[28]
port 437 nsew
flabel metal3 s -424 621509 56 621579 0 FreeSans 400 0 0 0 gpio_analog_pol[28]
port 525 nsew
flabel metal3 s -424 618473 56 618543 0 FreeSans 400 0 0 0 gpio_analog_sel[28]
port 481 nsew
flabel metal3 s -424 622153 56 622223 0 FreeSans 400 0 0 0 gpio_dm0[28]
port 569 nsew
flabel metal3 s -424 623993 56 624063 0 FreeSans 400 0 0 0 gpio_dm1[28]
port 613 nsew
flabel metal3 s -424 617829 56 617899 0 FreeSans 400 0 0 0 gpio_dm2[28]
port 657 nsew
flabel metal3 s -424 617185 56 617255 0 FreeSans 400 0 0 0 gpio_holdover[28]
port 393 nsew
flabel metal3 s -424 614149 56 614219 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[28]
port 261 nsew
flabel metal3 s -424 620957 56 621027 0 FreeSans 400 0 0 0 gpio_inp_dis[28]
port 217 nsew
flabel metal3 s -424 613505 56 613575 0 FreeSans 400 0 0 0 gpio_oeb[28]
port 173 nsew
flabel metal3 s -424 616633 56 616703 0 FreeSans 400 0 0 0 gpio_out[28]
port 129 nsew
flabel metal3 s -424 625833 56 625903 0 FreeSans 400 0 0 0 gpio_slow_sel[28]
port 349 nsew
flabel metal3 s -424 614793 56 614863 0 FreeSans 400 0 0 0 gpio_vtrip_sel[28]
port 305 nsew
flabel metal3 s -424 627673 56 627743 0 FreeSans 400 0 0 0 gpio_in[28]
port 701 nsew
flabel metal3 s -424 579597 56 579667 0 FreeSans 400 0 0 0 gpio_analog_en[29]
port 436 nsew
flabel metal3 s -424 578309 56 578379 0 FreeSans 400 0 0 0 gpio_analog_pol[29]
port 524 nsew
flabel metal3 s -424 575273 56 575343 0 FreeSans 400 0 0 0 gpio_analog_sel[29]
port 480 nsew
flabel metal3 s -424 578953 56 579023 0 FreeSans 400 0 0 0 gpio_dm0[29]
port 568 nsew
flabel metal3 s -424 580793 56 580863 0 FreeSans 400 0 0 0 gpio_dm1[29]
port 612 nsew
flabel metal3 s -424 574629 56 574699 0 FreeSans 400 0 0 0 gpio_dm2[29]
port 656 nsew
flabel metal3 s -424 573985 56 574055 0 FreeSans 400 0 0 0 gpio_holdover[29]
port 392 nsew
flabel metal3 s -424 570949 56 571019 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[29]
port 260 nsew
flabel metal3 s -424 577757 56 577827 0 FreeSans 400 0 0 0 gpio_inp_dis[29]
port 216 nsew
flabel metal3 s -424 570305 56 570375 0 FreeSans 400 0 0 0 gpio_oeb[29]
port 172 nsew
flabel metal3 s -424 573433 56 573503 0 FreeSans 400 0 0 0 gpio_out[29]
port 128 nsew
flabel metal3 s -424 582633 56 582703 0 FreeSans 400 0 0 0 gpio_slow_sel[29]
port 348 nsew
flabel metal3 s -424 571593 56 571663 0 FreeSans 400 0 0 0 gpio_vtrip_sel[29]
port 304 nsew
flabel metal3 s -424 584473 56 584543 0 FreeSans 400 0 0 0 gpio_in[29]
port 700 nsew
flabel metal3 s -424 536397 56 536467 0 FreeSans 400 0 0 0 gpio_analog_en[30]
port 435 nsew
flabel metal3 s -424 535109 56 535179 0 FreeSans 400 0 0 0 gpio_analog_pol[30]
port 523 nsew
flabel metal3 s -424 532073 56 532143 0 FreeSans 400 0 0 0 gpio_analog_sel[30]
port 479 nsew
flabel metal3 s -424 712877 56 712947 0 FreeSans 400 0 0 0 gpio_loopback_one[26]
port 835 nsew
flabel metal3 s -424 669677 56 669747 0 FreeSans 400 0 0 0 gpio_loopback_one[27]
port 834 nsew
flabel metal3 s -424 626477 56 626547 0 FreeSans 400 0 0 0 gpio_loopback_one[28]
port 833 nsew
flabel metal3 s -424 583277 56 583347 0 FreeSans 400 0 0 0 gpio_loopback_one[29]
port 832 nsew
flabel metal3 s -424 540077 56 540147 0 FreeSans 400 0 0 0 gpio_loopback_one[30]
port 831 nsew
flabel metal3 s -424 496877 56 496947 0 FreeSans 400 0 0 0 gpio_loopback_one[31]
port 830 nsew
flabel metal3 s -424 193993 56 194064 0 FreeSans 400 0 0 0 gpio_dm1[36]
port 605 nsew
flabel metal3 s -424 187829 56 187900 0 FreeSans 400 0 0 0 gpio_dm2[36]
port 649 nsew
flabel metal3 s -424 187185 56 187256 0 FreeSans 400 0 0 0 gpio_holdover[36]
port 385 nsew
flabel metal3 s -424 184149 56 184220 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[36]
port 253 nsew
flabel metal3 s -424 190957 56 191028 0 FreeSans 400 0 0 0 gpio_inp_dis[36]
port 209 nsew
flabel metal3 s -424 183505 56 183576 0 FreeSans 400 0 0 0 gpio_oeb[36]
port 165 nsew
flabel metal3 s -424 186633 56 186704 0 FreeSans 400 0 0 0 gpio_out[36]
port 121 nsew
flabel metal3 s -424 195833 56 195904 0 FreeSans 400 0 0 0 gpio_slow_sel[36]
port 341 nsew
flabel metal3 s -424 184793 56 184864 0 FreeSans 400 0 0 0 gpio_vtrip_sel[36]
port 297 nsew
flabel metal3 s -424 197673 56 197744 0 FreeSans 400 0 0 0 gpio_in[36]
port 693 nsew
flabel metal3 s -424 149597 56 149668 0 FreeSans 400 0 0 0 gpio_analog_en[37]
port 428 nsew
flabel metal3 s -424 148309 56 148380 0 FreeSans 400 0 0 0 gpio_analog_pol[37]
port 516 nsew
flabel metal3 s -424 145273 56 145344 0 FreeSans 400 0 0 0 gpio_analog_sel[37]
port 472 nsew
flabel metal3 s -424 148953 56 149024 0 FreeSans 400 0 0 0 gpio_dm0[37]
port 560 nsew
flabel metal3 s -424 150793 56 150864 0 FreeSans 400 0 0 0 gpio_dm1[37]
port 604 nsew
flabel metal3 s -424 144629 56 144700 0 FreeSans 400 0 0 0 gpio_dm2[37]
port 648 nsew
flabel metal3 s -424 143985 56 144056 0 FreeSans 400 0 0 0 gpio_holdover[37]
port 384 nsew
flabel metal3 s -424 140949 56 141020 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[37]
port 252 nsew
flabel metal3 s -424 140305 56 140376 0 FreeSans 400 0 0 0 gpio_oeb[37]
port 164 nsew
flabel metal3 s -424 143433 56 143504 0 FreeSans 400 0 0 0 gpio_out[37]
port 120 nsew
flabel metal3 s -424 152633 56 152704 0 FreeSans 400 0 0 0 gpio_slow_sel[37]
port 340 nsew
flabel metal3 s -424 154473 56 154544 0 FreeSans 400 0 0 0 gpio_in[37]
port 692 nsew
flabel metal3 s -424 365597 56 365667 0 FreeSans 400 0 0 0 gpio_analog_en[32]
port 433 nsew
flabel metal3 s -424 364309 56 364379 0 FreeSans 400 0 0 0 gpio_analog_pol[32]
port 521 nsew
flabel metal3 s -424 361273 56 361343 0 FreeSans 400 0 0 0 gpio_analog_sel[32]
port 477 nsew
flabel metal3 s -424 364953 56 365023 0 FreeSans 400 0 0 0 gpio_dm0[32]
port 565 nsew
flabel metal3 s -424 366793 56 366863 0 FreeSans 400 0 0 0 gpio_dm1[32]
port 609 nsew
flabel metal3 s -424 360629 56 360699 0 FreeSans 400 0 0 0 gpio_dm2[32]
port 653 nsew
flabel metal3 s -424 359985 56 360055 0 FreeSans 400 0 0 0 gpio_holdover[32]
port 389 nsew
flabel metal3 s -424 356949 56 357019 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[32]
port 257 nsew
flabel metal3 s -424 363757 56 363827 0 FreeSans 400 0 0 0 gpio_inp_dis[32]
port 213 nsew
flabel metal3 s -424 356305 56 356375 0 FreeSans 400 0 0 0 gpio_oeb[32]
port 169 nsew
flabel metal3 s -424 359433 56 359503 0 FreeSans 400 0 0 0 gpio_out[32]
port 125 nsew
flabel metal3 s -424 368633 56 368703 0 FreeSans 400 0 0 0 gpio_slow_sel[32]
port 345 nsew
flabel metal3 s -424 357593 56 357663 0 FreeSans 400 0 0 0 gpio_vtrip_sel[32]
port 301 nsew
flabel metal3 s -424 370473 56 370543 0 FreeSans 400 0 0 0 gpio_in[32]
port 697 nsew
flabel metal3 s -424 322397 56 322467 0 FreeSans 400 0 0 0 gpio_analog_en[33]
port 432 nsew
flabel metal3 s -424 318073 56 318143 0 FreeSans 400 0 0 0 gpio_analog_sel[33]
port 476 nsew
flabel metal3 s -424 323593 56 323663 0 FreeSans 400 0 0 0 gpio_dm1[33]
port 608 nsew
flabel metal3 s -424 317429 56 317499 0 FreeSans 400 0 0 0 gpio_dm2[33]
port 652 nsew
flabel metal3 s -424 321753 56 321823 0 FreeSans 400 0 0 0 gpio_dm0[33]
port 564 nsew
flabel metal3 s -424 316785 56 316855 0 FreeSans 400 0 0 0 gpio_holdover[33]
port 388 nsew
flabel metal3 s -424 313749 56 313819 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[33]
port 256 nsew
flabel metal3 s -424 320557 56 320627 0 FreeSans 400 0 0 0 gpio_inp_dis[33]
port 212 nsew
flabel metal3 s -424 313105 56 313175 0 FreeSans 400 0 0 0 gpio_oeb[33]
port 168 nsew
flabel metal3 s -424 316233 56 316303 0 FreeSans 400 0 0 0 gpio_out[33]
port 124 nsew
flabel metal3 s -424 325433 56 325503 0 FreeSans 400 0 0 0 gpio_slow_sel[33]
port 344 nsew
flabel metal3 s -424 314393 56 314463 0 FreeSans 400 0 0 0 gpio_vtrip_sel[33]
port 300 nsew
flabel metal3 s -424 327273 56 327343 0 FreeSans 400 0 0 0 gpio_in[33]
port 696 nsew
flabel metal3 s -424 279197 56 279267 0 FreeSans 400 0 0 0 gpio_analog_en[34]
port 431 nsew
flabel metal3 s -424 277909 56 277979 0 FreeSans 400 0 0 0 gpio_analog_pol[34]
port 519 nsew
flabel metal3 s -424 274873 56 274943 0 FreeSans 400 0 0 0 gpio_analog_sel[34]
port 475 nsew
flabel metal3 s -424 278553 56 278623 0 FreeSans 400 0 0 0 gpio_dm0[34]
port 563 nsew
flabel metal3 s -424 280393 56 280463 0 FreeSans 400 0 0 0 gpio_dm1[34]
port 607 nsew
flabel metal3 s -424 274229 56 274299 0 FreeSans 400 0 0 0 gpio_dm2[34]
port 651 nsew
flabel metal3 s -424 273585 56 273655 0 FreeSans 400 0 0 0 gpio_holdover[34]
port 387 nsew
flabel metal3 s -424 270549 56 270619 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[34]
port 255 nsew
flabel metal3 s -424 277357 56 277427 0 FreeSans 400 0 0 0 gpio_inp_dis[34]
port 211 nsew
flabel metal3 s -424 269905 56 269975 0 FreeSans 400 0 0 0 gpio_oeb[34]
port 167 nsew
flabel metal3 s -424 273033 56 273103 0 FreeSans 400 0 0 0 gpio_out[34]
port 123 nsew
flabel metal3 s -424 282233 56 282303 0 FreeSans 400 0 0 0 gpio_slow_sel[34]
port 343 nsew
flabel metal3 s -424 271193 56 271263 0 FreeSans 400 0 0 0 gpio_vtrip_sel[34]
port 299 nsew
flabel metal3 s -424 284073 56 284143 0 FreeSans 400 0 0 0 gpio_in[34]
port 695 nsew
flabel metal3 s -424 235997 56 236067 0 FreeSans 400 0 0 0 gpio_analog_en[35]
port 430 nsew
flabel metal3 s -424 234709 56 234779 0 FreeSans 400 0 0 0 gpio_analog_pol[35]
port 518 nsew
flabel metal3 s -424 231673 56 231743 0 FreeSans 400 0 0 0 gpio_analog_sel[35]
port 474 nsew
flabel metal3 s -424 235353 56 235423 0 FreeSans 400 0 0 0 gpio_dm0[35]
port 562 nsew
flabel metal3 s -424 237193 56 237263 0 FreeSans 400 0 0 0 gpio_dm1[35]
port 606 nsew
flabel metal3 s -424 231029 56 231099 0 FreeSans 400 0 0 0 gpio_dm2[35]
port 650 nsew
flabel metal3 s -424 230385 56 230455 0 FreeSans 400 0 0 0 gpio_holdover[35]
port 386 nsew
flabel metal3 s -424 227349 56 227419 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[35]
port 254 nsew
flabel metal3 s -424 234157 56 234227 0 FreeSans 400 0 0 0 gpio_inp_dis[35]
port 210 nsew
flabel metal3 s -424 226705 56 226775 0 FreeSans 400 0 0 0 gpio_oeb[35]
port 166 nsew
flabel metal3 s -424 229833 56 229903 0 FreeSans 400 0 0 0 gpio_out[35]
port 122 nsew
flabel metal3 s -424 239033 56 239103 0 FreeSans 400 0 0 0 gpio_slow_sel[35]
port 342 nsew
flabel metal3 s -424 227993 56 228063 0 FreeSans 400 0 0 0 gpio_vtrip_sel[35]
port 298 nsew
flabel metal3 s -424 240873 56 240943 0 FreeSans 400 0 0 0 gpio_in[35]
port 694 nsew
flabel metal3 s -424 192797 56 192868 0 FreeSans 400 0 0 0 gpio_analog_en[36]
port 429 nsew
flabel metal3 s -424 191509 56 191580 0 FreeSans 400 0 0 0 gpio_analog_pol[36]
port 517 nsew
flabel metal3 s -424 188473 56 188544 0 FreeSans 400 0 0 0 gpio_analog_sel[36]
port 473 nsew
flabel metal3 s -424 192153 56 192224 0 FreeSans 400 0 0 0 gpio_dm0[36]
port 561 nsew
flabel metal3 s -424 369277 56 369347 0 FreeSans 400 0 0 0 gpio_loopback_one[32]
port 829 nsew
flabel metal3 s -424 326077 56 326147 0 FreeSans 400 0 0 0 gpio_loopback_one[33]
port 828 nsew
flabel metal3 s -424 282877 56 282947 0 FreeSans 400 0 0 0 gpio_loopback_one[34]
port 827 nsew
flabel metal3 s -424 239677 56 239747 0 FreeSans 400 0 0 0 gpio_loopback_one[35]
port 826 nsew
flabel metal3 s -424 196477 56 196548 0 FreeSans 400 0 0 0 gpio_loopback_one[36]
port 825 nsew
flabel metal3 s -424 153277 56 153348 0 FreeSans 400 0 0 0 gpio_loopback_one[37]
port 824 nsew
flabel metal3 s -424 147757 56 147828 0 FreeSans 400 0 0 0 gpio_inp_dis[37]
port 208 nsew
flabel metal3 s -424 742553 56 742623 0 FreeSans 400 0 0 0 gpio_in_h[25]
port 748 nsew
flabel metal3 s -424 699353 56 699423 0 FreeSans 400 0 0 0 gpio_in_h[26]
port 747 nsew
flabel metal3 s -424 656153 56 656223 0 FreeSans 400 0 0 0 gpio_in_h[27]
port 746 nsew
flabel metal3 s -424 612953 56 613023 0 FreeSans 400 0 0 0 gpio_in_h[28]
port 745 nsew
flabel metal3 s -424 569753 56 569823 0 FreeSans 400 0 0 0 gpio_in_h[29]
port 744 nsew
flabel metal3 s -424 526553 56 526623 0 FreeSans 400 0 0 0 gpio_in_h[30]
port 743 nsew
flabel metal3 s -424 483353 56 483423 0 FreeSans 400 0 0 0 gpio_in_h[31]
port 742 nsew
flabel metal3 s -424 355753 56 355823 0 FreeSans 400 0 0 0 gpio_in_h[32]
port 741 nsew
flabel metal3 s -424 312553 56 312623 0 FreeSans 400 0 0 0 gpio_in_h[33]
port 740 nsew
flabel metal3 s -424 269353 56 269423 0 FreeSans 400 0 0 0 gpio_in_h[34]
port 739 nsew
flabel metal3 s -424 226153 56 226223 0 FreeSans 400 0 0 0 gpio_in_h[35]
port 738 nsew
flabel metal3 s -424 182953 56 183024 0 FreeSans 400 0 0 0 gpio_in_h[36]
port 737 nsew
flabel metal3 s -424 139753 56 139824 0 FreeSans 400 0 0 0 gpio_in_h[37]
port 736 nsew
flabel metal3 s -424 754789 56 754859 0 FreeSans 400 0 0 0 analog_io[25]
port 880 nsew
flabel metal3 s -424 711589 56 711659 0 FreeSans 400 0 0 0 analog_io[26]
port 879 nsew
flabel metal3 s -424 668389 56 668459 0 FreeSans 400 0 0 0 analog_io[27]
port 878 nsew
flabel metal3 s -424 625189 56 625259 0 FreeSans 400 0 0 0 analog_io[28]
port 877 nsew
flabel metal3 s -424 581989 56 582059 0 FreeSans 400 0 0 0 analog_io[29]
port 876 nsew
flabel metal3 s -424 538789 56 538859 0 FreeSans 400 0 0 0 analog_io[30]
port 875 nsew
flabel metal3 s -424 495589 56 495659 0 FreeSans 400 0 0 0 analog_io[31]
port 874 nsew
flabel metal3 s -424 367989 56 368059 0 FreeSans 400 0 0 0 analog_io[32]
port 873 nsew
flabel metal3 s -424 324789 56 324859 0 FreeSans 400 0 0 0 analog_io[33]
port 872 nsew
flabel metal3 s -424 281589 56 281659 0 FreeSans 400 0 0 0 analog_io[34]
port 871 nsew
flabel metal3 s -424 238389 56 238459 0 FreeSans 400 0 0 0 analog_io[35]
port 870 nsew
flabel metal3 s -424 195189 56 195260 0 FreeSans 400 0 0 0 analog_io[36]
port 869 nsew
flabel metal3 s -424 151989 56 152060 0 FreeSans 400 0 0 0 analog_io[37]
port 868 nsew
flabel metal3 s -424 752949 56 753019 0 FreeSans 400 0 0 0 analog_noesd_io[25]
port 924 nsew
flabel metal3 s -424 709749 56 709819 0 FreeSans 400 0 0 0 analog_noesd_io[26]
port 923 nsew
flabel metal3 s -424 666549 56 666619 0 FreeSans 400 0 0 0 analog_noesd_io[27]
port 922 nsew
flabel metal3 s -424 623349 56 623419 0 FreeSans 400 0 0 0 analog_noesd_io[28]
port 921 nsew
flabel metal3 s -424 580149 56 580219 0 FreeSans 400 0 0 0 analog_noesd_io[29]
port 920 nsew
flabel metal3 s -424 536949 56 537019 0 FreeSans 400 0 0 0 analog_noesd_io[30]
port 919 nsew
flabel metal3 s -424 493749 56 493819 0 FreeSans 400 0 0 0 analog_noesd_io[31]
port 918 nsew
flabel metal3 s -424 366149 56 366219 0 FreeSans 400 0 0 0 analog_noesd_io[32]
port 917 nsew
flabel metal3 s -424 322949 56 323019 0 FreeSans 400 0 0 0 analog_noesd_io[33]
port 916 nsew
flabel metal3 s -424 279749 56 279819 0 FreeSans 400 0 0 0 analog_noesd_io[34]
port 915 nsew
flabel metal3 s -424 236549 56 236619 0 FreeSans 400 0 0 0 analog_noesd_io[35]
port 914 nsew
flabel metal3 s -424 193349 56 193420 0 FreeSans 400 0 0 0 analog_noesd_io[36]
port 913 nsew
flabel metal3 s -424 150149 56 150220 0 FreeSans 400 0 0 0 analog_noesd_io[37]
port 912 nsew
flabel metal3 s -424 744393 56 744463 0 FreeSans 400 0 0 0 gpio_vtrip_sel[25]
port 308 nsew
flabel metal3 s -424 321116 56 321172 0 FreeSans 400 0 0 0 gpio_analog_pol[33]
port 520 nsew
<< properties >>
string FIXED_BBOX 0 0 633326 953326
<< end >>
