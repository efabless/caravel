magic
tech sky130A
magscale 1 2
timestamp 1675864079
<< obsli1 >>
rect 1104 2159 74888 107729
<< obsm1 >>
rect 106 1504 75978 107840
<< metal2 >>
rect 2870 109390 2926 110190
rect 3422 109390 3478 110190
rect 3974 109390 4030 110190
rect 4526 109390 4582 110190
rect 5078 109390 5134 110190
rect 5630 109390 5686 110190
rect 6182 109390 6238 110190
rect 6734 109390 6790 110190
rect 7286 109390 7342 110190
rect 7838 109390 7894 110190
rect 8390 109390 8446 110190
rect 8942 109390 8998 110190
rect 9494 109390 9550 110190
rect 10046 109390 10102 110190
rect 10598 109390 10654 110190
rect 11150 109390 11206 110190
rect 11702 109390 11758 110190
rect 12254 109390 12310 110190
rect 12806 109390 12862 110190
rect 13358 109390 13414 110190
rect 13910 109390 13966 110190
rect 14462 109390 14518 110190
rect 15014 109390 15070 110190
rect 15566 109390 15622 110190
rect 16118 109390 16174 110190
rect 16670 109390 16726 110190
rect 17222 109390 17278 110190
rect 17774 109390 17830 110190
rect 18326 109390 18382 110190
rect 18878 109390 18934 110190
rect 19430 109390 19486 110190
rect 19982 109390 20038 110190
rect 20534 109390 20590 110190
rect 21086 109390 21142 110190
rect 21638 109390 21694 110190
rect 22190 109390 22246 110190
rect 22742 109390 22798 110190
rect 23294 109390 23350 110190
rect 23846 109390 23902 110190
rect 24398 109390 24454 110190
rect 24950 109390 25006 110190
rect 25502 109390 25558 110190
rect 26054 109390 26110 110190
rect 26606 109390 26662 110190
rect 27158 109390 27214 110190
rect 27710 109390 27766 110190
rect 28262 109390 28318 110190
rect 28814 109390 28870 110190
rect 29366 109390 29422 110190
rect 29918 109390 29974 110190
rect 30470 109390 30526 110190
rect 31022 109390 31078 110190
rect 31574 109390 31630 110190
rect 32126 109390 32182 110190
rect 32678 109390 32734 110190
rect 33230 109390 33286 110190
rect 33782 109390 33838 110190
rect 34334 109390 34390 110190
rect 34886 109390 34942 110190
rect 35438 109390 35494 110190
rect 35990 109390 36046 110190
rect 36542 109390 36598 110190
rect 37094 109390 37150 110190
rect 37646 109390 37702 110190
rect 38198 109390 38254 110190
rect 38750 109390 38806 110190
rect 39302 109390 39358 110190
rect 39854 109390 39910 110190
rect 40406 109390 40462 110190
rect 40958 109390 41014 110190
rect 41510 109390 41566 110190
rect 42062 109390 42118 110190
rect 42614 109390 42670 110190
rect 43166 109390 43222 110190
rect 43718 109390 43774 110190
rect 44270 109390 44326 110190
rect 44822 109390 44878 110190
rect 45374 109390 45430 110190
rect 45926 109390 45982 110190
rect 46478 109390 46534 110190
rect 47030 109390 47086 110190
rect 47582 109390 47638 110190
rect 48134 109390 48190 110190
rect 48686 109390 48742 110190
rect 49238 109390 49294 110190
rect 49790 109390 49846 110190
rect 50342 109390 50398 110190
rect 50894 109390 50950 110190
rect 51446 109390 51502 110190
rect 51998 109390 52054 110190
rect 52550 109390 52606 110190
rect 53102 109390 53158 110190
rect 53654 109390 53710 110190
rect 54206 109390 54262 110190
rect 54758 109390 54814 110190
rect 55310 109390 55366 110190
rect 55862 109390 55918 110190
rect 56414 109390 56470 110190
rect 56966 109390 57022 110190
rect 57518 109390 57574 110190
rect 58070 109390 58126 110190
rect 58622 109390 58678 110190
rect 59174 109390 59230 110190
rect 59726 109390 59782 110190
rect 60278 109390 60334 110190
rect 60830 109390 60886 110190
rect 61382 109390 61438 110190
rect 61934 109390 61990 110190
rect 62486 109390 62542 110190
rect 63038 109390 63094 110190
rect 63590 109390 63646 110190
rect 64142 109390 64198 110190
rect 64694 109390 64750 110190
rect 65246 109390 65302 110190
rect 65798 109390 65854 110190
rect 66350 109390 66406 110190
rect 66902 109390 66958 110190
rect 67454 109390 67510 110190
rect 68006 109390 68062 110190
rect 68558 109390 68614 110190
rect 69110 109390 69166 110190
rect 69662 109390 69718 110190
rect 70214 109390 70270 110190
rect 70766 109390 70822 110190
rect 71318 109390 71374 110190
rect 71870 109390 71926 110190
rect 72422 109390 72478 110190
rect 72974 109390 73030 110190
rect 4066 0 4122 800
rect 4802 0 4858 800
rect 5538 0 5594 800
rect 6274 0 6330 800
rect 7010 0 7066 800
rect 7746 0 7802 800
rect 8482 0 8538 800
rect 9218 0 9274 800
rect 9954 0 10010 800
rect 10690 0 10746 800
rect 11426 0 11482 800
rect 12162 0 12218 800
rect 12898 0 12954 800
rect 13634 0 13690 800
rect 14370 0 14426 800
rect 15106 0 15162 800
rect 15842 0 15898 800
rect 16578 0 16634 800
rect 17314 0 17370 800
rect 18050 0 18106 800
rect 18786 0 18842 800
rect 19522 0 19578 800
rect 20258 0 20314 800
rect 20994 0 21050 800
rect 21730 0 21786 800
rect 22466 0 22522 800
rect 23202 0 23258 800
rect 23938 0 23994 800
rect 24674 0 24730 800
rect 25410 0 25466 800
rect 26146 0 26202 800
rect 26882 0 26938 800
rect 27618 0 27674 800
rect 28354 0 28410 800
rect 29090 0 29146 800
rect 29826 0 29882 800
rect 30562 0 30618 800
rect 31298 0 31354 800
rect 32034 0 32090 800
rect 32770 0 32826 800
rect 33506 0 33562 800
rect 34242 0 34298 800
rect 34978 0 35034 800
rect 35714 0 35770 800
rect 36450 0 36506 800
rect 37186 0 37242 800
rect 37922 0 37978 800
rect 38658 0 38714 800
rect 39394 0 39450 800
rect 40130 0 40186 800
rect 40866 0 40922 800
rect 41602 0 41658 800
rect 42338 0 42394 800
rect 43074 0 43130 800
rect 43810 0 43866 800
rect 44546 0 44602 800
rect 45282 0 45338 800
rect 46018 0 46074 800
rect 46754 0 46810 800
rect 47490 0 47546 800
rect 48226 0 48282 800
rect 48962 0 49018 800
rect 49698 0 49754 800
rect 50434 0 50490 800
rect 51170 0 51226 800
rect 51906 0 51962 800
rect 52642 0 52698 800
rect 53378 0 53434 800
rect 54114 0 54170 800
rect 54850 0 54906 800
rect 55586 0 55642 800
rect 56322 0 56378 800
rect 57058 0 57114 800
rect 57794 0 57850 800
rect 58530 0 58586 800
rect 59266 0 59322 800
rect 60002 0 60058 800
rect 60738 0 60794 800
rect 61474 0 61530 800
rect 62210 0 62266 800
rect 62946 0 63002 800
rect 63682 0 63738 800
rect 64418 0 64474 800
rect 65154 0 65210 800
rect 65890 0 65946 800
rect 66626 0 66682 800
rect 67362 0 67418 800
rect 68098 0 68154 800
rect 68834 0 68890 800
rect 69570 0 69626 800
rect 70306 0 70362 800
rect 71042 0 71098 800
rect 71778 0 71834 800
<< obsm2 >>
rect 110 109334 2814 109426
rect 2982 109334 3366 109426
rect 3534 109334 3918 109426
rect 4086 109334 4470 109426
rect 4638 109334 5022 109426
rect 5190 109334 5574 109426
rect 5742 109334 6126 109426
rect 6294 109334 6678 109426
rect 6846 109334 7230 109426
rect 7398 109334 7782 109426
rect 7950 109334 8334 109426
rect 8502 109334 8886 109426
rect 9054 109334 9438 109426
rect 9606 109334 9990 109426
rect 10158 109334 10542 109426
rect 10710 109334 11094 109426
rect 11262 109334 11646 109426
rect 11814 109334 12198 109426
rect 12366 109334 12750 109426
rect 12918 109334 13302 109426
rect 13470 109334 13854 109426
rect 14022 109334 14406 109426
rect 14574 109334 14958 109426
rect 15126 109334 15510 109426
rect 15678 109334 16062 109426
rect 16230 109334 16614 109426
rect 16782 109334 17166 109426
rect 17334 109334 17718 109426
rect 17886 109334 18270 109426
rect 18438 109334 18822 109426
rect 18990 109334 19374 109426
rect 19542 109334 19926 109426
rect 20094 109334 20478 109426
rect 20646 109334 21030 109426
rect 21198 109334 21582 109426
rect 21750 109334 22134 109426
rect 22302 109334 22686 109426
rect 22854 109334 23238 109426
rect 23406 109334 23790 109426
rect 23958 109334 24342 109426
rect 24510 109334 24894 109426
rect 25062 109334 25446 109426
rect 25614 109334 25998 109426
rect 26166 109334 26550 109426
rect 26718 109334 27102 109426
rect 27270 109334 27654 109426
rect 27822 109334 28206 109426
rect 28374 109334 28758 109426
rect 28926 109334 29310 109426
rect 29478 109334 29862 109426
rect 30030 109334 30414 109426
rect 30582 109334 30966 109426
rect 31134 109334 31518 109426
rect 31686 109334 32070 109426
rect 32238 109334 32622 109426
rect 32790 109334 33174 109426
rect 33342 109334 33726 109426
rect 33894 109334 34278 109426
rect 34446 109334 34830 109426
rect 34998 109334 35382 109426
rect 35550 109334 35934 109426
rect 36102 109334 36486 109426
rect 36654 109334 37038 109426
rect 37206 109334 37590 109426
rect 37758 109334 38142 109426
rect 38310 109334 38694 109426
rect 38862 109334 39246 109426
rect 39414 109334 39798 109426
rect 39966 109334 40350 109426
rect 40518 109334 40902 109426
rect 41070 109334 41454 109426
rect 41622 109334 42006 109426
rect 42174 109334 42558 109426
rect 42726 109334 43110 109426
rect 43278 109334 43662 109426
rect 43830 109334 44214 109426
rect 44382 109334 44766 109426
rect 44934 109334 45318 109426
rect 45486 109334 45870 109426
rect 46038 109334 46422 109426
rect 46590 109334 46974 109426
rect 47142 109334 47526 109426
rect 47694 109334 48078 109426
rect 48246 109334 48630 109426
rect 48798 109334 49182 109426
rect 49350 109334 49734 109426
rect 49902 109334 50286 109426
rect 50454 109334 50838 109426
rect 51006 109334 51390 109426
rect 51558 109334 51942 109426
rect 52110 109334 52494 109426
rect 52662 109334 53046 109426
rect 53214 109334 53598 109426
rect 53766 109334 54150 109426
rect 54318 109334 54702 109426
rect 54870 109334 55254 109426
rect 55422 109334 55806 109426
rect 55974 109334 56358 109426
rect 56526 109334 56910 109426
rect 57078 109334 57462 109426
rect 57630 109334 58014 109426
rect 58182 109334 58566 109426
rect 58734 109334 59118 109426
rect 59286 109334 59670 109426
rect 59838 109334 60222 109426
rect 60390 109334 60774 109426
rect 60942 109334 61326 109426
rect 61494 109334 61878 109426
rect 62046 109334 62430 109426
rect 62598 109334 62982 109426
rect 63150 109334 63534 109426
rect 63702 109334 64086 109426
rect 64254 109334 64638 109426
rect 64806 109334 65190 109426
rect 65358 109334 65742 109426
rect 65910 109334 66294 109426
rect 66462 109334 66846 109426
rect 67014 109334 67398 109426
rect 67566 109334 67950 109426
rect 68118 109334 68502 109426
rect 68670 109334 69054 109426
rect 69222 109334 69606 109426
rect 69774 109334 70158 109426
rect 70326 109334 70710 109426
rect 70878 109334 71262 109426
rect 71430 109334 71814 109426
rect 71982 109334 72366 109426
rect 72534 109334 72918 109426
rect 73086 109334 75974 109426
rect 110 856 75974 109334
rect 110 734 4010 856
rect 4178 734 4746 856
rect 4914 734 5482 856
rect 5650 734 6218 856
rect 6386 734 6954 856
rect 7122 734 7690 856
rect 7858 734 8426 856
rect 8594 734 9162 856
rect 9330 734 9898 856
rect 10066 734 10634 856
rect 10802 734 11370 856
rect 11538 734 12106 856
rect 12274 734 12842 856
rect 13010 734 13578 856
rect 13746 734 14314 856
rect 14482 734 15050 856
rect 15218 734 15786 856
rect 15954 734 16522 856
rect 16690 734 17258 856
rect 17426 734 17994 856
rect 18162 734 18730 856
rect 18898 734 19466 856
rect 19634 734 20202 856
rect 20370 734 20938 856
rect 21106 734 21674 856
rect 21842 734 22410 856
rect 22578 734 23146 856
rect 23314 734 23882 856
rect 24050 734 24618 856
rect 24786 734 25354 856
rect 25522 734 26090 856
rect 26258 734 26826 856
rect 26994 734 27562 856
rect 27730 734 28298 856
rect 28466 734 29034 856
rect 29202 734 29770 856
rect 29938 734 30506 856
rect 30674 734 31242 856
rect 31410 734 31978 856
rect 32146 734 32714 856
rect 32882 734 33450 856
rect 33618 734 34186 856
rect 34354 734 34922 856
rect 35090 734 35658 856
rect 35826 734 36394 856
rect 36562 734 37130 856
rect 37298 734 37866 856
rect 38034 734 38602 856
rect 38770 734 39338 856
rect 39506 734 40074 856
rect 40242 734 40810 856
rect 40978 734 41546 856
rect 41714 734 42282 856
rect 42450 734 43018 856
rect 43186 734 43754 856
rect 43922 734 44490 856
rect 44658 734 45226 856
rect 45394 734 45962 856
rect 46130 734 46698 856
rect 46866 734 47434 856
rect 47602 734 48170 856
rect 48338 734 48906 856
rect 49074 734 49642 856
rect 49810 734 50378 856
rect 50546 734 51114 856
rect 51282 734 51850 856
rect 52018 734 52586 856
rect 52754 734 53322 856
rect 53490 734 54058 856
rect 54226 734 54794 856
rect 54962 734 55530 856
rect 55698 734 56266 856
rect 56434 734 57002 856
rect 57170 734 57738 856
rect 57906 734 58474 856
rect 58642 734 59210 856
rect 59378 734 59946 856
rect 60114 734 60682 856
rect 60850 734 61418 856
rect 61586 734 62154 856
rect 62322 734 62890 856
rect 63058 734 63626 856
rect 63794 734 64362 856
rect 64530 734 65098 856
rect 65266 734 65834 856
rect 66002 734 66570 856
rect 66738 734 67306 856
rect 67474 734 68042 856
rect 68210 734 68778 856
rect 68946 734 69514 856
rect 69682 734 70250 856
rect 70418 734 70986 856
rect 71154 734 71722 856
rect 71890 734 75974 856
<< metal3 >>
rect 0 107992 800 108112
rect 75246 107176 76046 107296
rect 0 106360 800 106480
rect 75246 105544 76046 105664
rect 0 104728 800 104848
rect 75246 103912 76046 104032
rect 0 103096 800 103216
rect 75246 102280 76046 102400
rect 0 101464 800 101584
rect 75246 100648 76046 100768
rect 0 99832 800 99952
rect 75246 99016 76046 99136
rect 0 98200 800 98320
rect 75246 97384 76046 97504
rect 0 96568 800 96688
rect 75246 95752 76046 95872
rect 0 94936 800 95056
rect 75246 94120 76046 94240
rect 0 93304 800 93424
rect 75246 92488 76046 92608
rect 0 91672 800 91792
rect 75246 90856 76046 90976
rect 0 90040 800 90160
rect 75246 89224 76046 89344
rect 0 88408 800 88528
rect 75246 87592 76046 87712
rect 0 86776 800 86896
rect 75246 85960 76046 86080
rect 0 85144 800 85264
rect 75246 84328 76046 84448
rect 0 83512 800 83632
rect 75246 82696 76046 82816
rect 0 81880 800 82000
rect 75246 81064 76046 81184
rect 0 80248 800 80368
rect 75246 79432 76046 79552
rect 0 78616 800 78736
rect 75246 77800 76046 77920
rect 0 76984 800 77104
rect 75246 76168 76046 76288
rect 0 75352 800 75472
rect 75246 74536 76046 74656
rect 0 73720 800 73840
rect 75246 72904 76046 73024
rect 0 72088 800 72208
rect 75246 71272 76046 71392
rect 0 70456 800 70576
rect 75246 69640 76046 69760
rect 0 68824 800 68944
rect 75246 68008 76046 68128
rect 0 67192 800 67312
rect 75246 66376 76046 66496
rect 0 65560 800 65680
rect 75246 64744 76046 64864
rect 0 63928 800 64048
rect 75246 63112 76046 63232
rect 0 62296 800 62416
rect 75246 61480 76046 61600
rect 0 60664 800 60784
rect 75246 59848 76046 59968
rect 0 59032 800 59152
rect 75246 58216 76046 58336
rect 0 57400 800 57520
rect 75246 56584 76046 56704
rect 0 55768 800 55888
rect 75246 54952 76046 55072
rect 0 54136 800 54256
rect 75246 53320 76046 53440
rect 0 52504 800 52624
rect 75246 51688 76046 51808
rect 0 50872 800 50992
rect 75246 50056 76046 50176
rect 0 49240 800 49360
rect 75246 48424 76046 48544
rect 0 47608 800 47728
rect 75246 46792 76046 46912
rect 0 45976 800 46096
rect 75246 45160 76046 45280
rect 0 44344 800 44464
rect 75246 43528 76046 43648
rect 0 42712 800 42832
rect 75246 41896 76046 42016
rect 0 41080 800 41200
rect 75246 40264 76046 40384
rect 0 39448 800 39568
rect 75246 38632 76046 38752
rect 0 37816 800 37936
rect 75246 37000 76046 37120
rect 0 36184 800 36304
rect 75246 35368 76046 35488
rect 0 34552 800 34672
rect 75246 33736 76046 33856
rect 0 32920 800 33040
rect 75246 32104 76046 32224
rect 0 31288 800 31408
rect 75246 30472 76046 30592
rect 0 29656 800 29776
rect 75246 28840 76046 28960
rect 0 28024 800 28144
rect 75246 27208 76046 27328
rect 0 26392 800 26512
rect 75246 25576 76046 25696
rect 0 24760 800 24880
rect 75246 23944 76046 24064
rect 0 23128 800 23248
rect 75246 22312 76046 22432
rect 0 21496 800 21616
rect 75246 20680 76046 20800
rect 0 19864 800 19984
rect 75246 19048 76046 19168
rect 0 18232 800 18352
rect 75246 17416 76046 17536
rect 0 16600 800 16720
rect 75246 15784 76046 15904
rect 0 14968 800 15088
rect 75246 14152 76046 14272
rect 0 13336 800 13456
rect 75246 12520 76046 12640
rect 0 11704 800 11824
rect 75246 10888 76046 11008
rect 0 10072 800 10192
rect 75246 9256 76046 9376
rect 0 8440 800 8560
rect 75246 7624 76046 7744
rect 0 6808 800 6928
rect 75246 5992 76046 6112
rect 0 5176 800 5296
rect 75246 4360 76046 4480
rect 0 3544 800 3664
rect 75246 2728 76046 2848
rect 0 1912 800 2032
<< obsm3 >>
rect 880 107912 75979 108085
rect 54 107376 75979 107912
rect 54 107096 75166 107376
rect 54 106560 75979 107096
rect 880 106280 75979 106560
rect 54 105744 75979 106280
rect 54 105464 75166 105744
rect 54 104928 75979 105464
rect 880 104648 75979 104928
rect 54 104112 75979 104648
rect 54 103832 75166 104112
rect 54 103296 75979 103832
rect 880 103016 75979 103296
rect 54 102480 75979 103016
rect 54 102200 75166 102480
rect 54 101664 75979 102200
rect 880 101384 75979 101664
rect 54 100848 75979 101384
rect 54 100568 75166 100848
rect 54 100032 75979 100568
rect 880 99752 75979 100032
rect 54 99216 75979 99752
rect 54 98936 75166 99216
rect 54 98400 75979 98936
rect 880 98120 75979 98400
rect 54 97584 75979 98120
rect 54 97304 75166 97584
rect 54 96768 75979 97304
rect 880 96488 75979 96768
rect 54 95952 75979 96488
rect 54 95672 75166 95952
rect 54 95136 75979 95672
rect 880 94856 75979 95136
rect 54 94320 75979 94856
rect 54 94040 75166 94320
rect 54 93504 75979 94040
rect 880 93224 75979 93504
rect 54 92688 75979 93224
rect 54 92408 75166 92688
rect 54 91872 75979 92408
rect 880 91592 75979 91872
rect 54 91056 75979 91592
rect 54 90776 75166 91056
rect 54 90240 75979 90776
rect 880 89960 75979 90240
rect 54 89424 75979 89960
rect 54 89144 75166 89424
rect 54 88608 75979 89144
rect 880 88328 75979 88608
rect 54 87792 75979 88328
rect 54 87512 75166 87792
rect 54 86976 75979 87512
rect 880 86696 75979 86976
rect 54 86160 75979 86696
rect 54 85880 75166 86160
rect 54 85344 75979 85880
rect 880 85064 75979 85344
rect 54 84528 75979 85064
rect 54 84248 75166 84528
rect 54 83712 75979 84248
rect 880 83432 75979 83712
rect 54 82896 75979 83432
rect 54 82616 75166 82896
rect 54 82080 75979 82616
rect 880 81800 75979 82080
rect 54 81264 75979 81800
rect 54 80984 75166 81264
rect 54 80448 75979 80984
rect 880 80168 75979 80448
rect 54 79632 75979 80168
rect 54 79352 75166 79632
rect 54 78816 75979 79352
rect 880 78536 75979 78816
rect 54 78000 75979 78536
rect 54 77720 75166 78000
rect 54 77184 75979 77720
rect 880 76904 75979 77184
rect 54 76368 75979 76904
rect 54 76088 75166 76368
rect 54 75552 75979 76088
rect 880 75272 75979 75552
rect 54 74736 75979 75272
rect 54 74456 75166 74736
rect 54 73920 75979 74456
rect 880 73640 75979 73920
rect 54 73104 75979 73640
rect 54 72824 75166 73104
rect 54 72288 75979 72824
rect 880 72008 75979 72288
rect 54 71472 75979 72008
rect 54 71192 75166 71472
rect 54 70656 75979 71192
rect 880 70376 75979 70656
rect 54 69840 75979 70376
rect 54 69560 75166 69840
rect 54 69024 75979 69560
rect 880 68744 75979 69024
rect 54 68208 75979 68744
rect 54 67928 75166 68208
rect 54 67392 75979 67928
rect 880 67112 75979 67392
rect 54 66576 75979 67112
rect 54 66296 75166 66576
rect 54 65760 75979 66296
rect 880 65480 75979 65760
rect 54 64944 75979 65480
rect 54 64664 75166 64944
rect 54 64128 75979 64664
rect 880 63848 75979 64128
rect 54 63312 75979 63848
rect 54 63032 75166 63312
rect 54 62496 75979 63032
rect 880 62216 75979 62496
rect 54 61680 75979 62216
rect 54 61400 75166 61680
rect 54 60864 75979 61400
rect 880 60584 75979 60864
rect 54 60048 75979 60584
rect 54 59768 75166 60048
rect 54 59232 75979 59768
rect 880 58952 75979 59232
rect 54 58416 75979 58952
rect 54 58136 75166 58416
rect 54 57600 75979 58136
rect 880 57320 75979 57600
rect 54 56784 75979 57320
rect 54 56504 75166 56784
rect 54 55968 75979 56504
rect 880 55688 75979 55968
rect 54 55152 75979 55688
rect 54 54872 75166 55152
rect 54 54336 75979 54872
rect 880 54056 75979 54336
rect 54 53520 75979 54056
rect 54 53240 75166 53520
rect 54 52704 75979 53240
rect 880 52424 75979 52704
rect 54 51888 75979 52424
rect 54 51608 75166 51888
rect 54 51072 75979 51608
rect 880 50792 75979 51072
rect 54 50256 75979 50792
rect 54 49976 75166 50256
rect 54 49440 75979 49976
rect 880 49160 75979 49440
rect 54 48624 75979 49160
rect 54 48344 75166 48624
rect 54 47808 75979 48344
rect 880 47528 75979 47808
rect 54 46992 75979 47528
rect 54 46712 75166 46992
rect 54 46176 75979 46712
rect 880 45896 75979 46176
rect 54 45360 75979 45896
rect 54 45080 75166 45360
rect 54 44544 75979 45080
rect 880 44264 75979 44544
rect 54 43728 75979 44264
rect 54 43448 75166 43728
rect 54 42912 75979 43448
rect 880 42632 75979 42912
rect 54 42096 75979 42632
rect 54 41816 75166 42096
rect 54 41280 75979 41816
rect 880 41000 75979 41280
rect 54 40464 75979 41000
rect 54 40184 75166 40464
rect 54 39648 75979 40184
rect 880 39368 75979 39648
rect 54 38832 75979 39368
rect 54 38552 75166 38832
rect 54 38016 75979 38552
rect 880 37736 75979 38016
rect 54 37200 75979 37736
rect 54 36920 75166 37200
rect 54 36384 75979 36920
rect 880 36104 75979 36384
rect 54 35568 75979 36104
rect 54 35288 75166 35568
rect 54 34752 75979 35288
rect 880 34472 75979 34752
rect 54 33936 75979 34472
rect 54 33656 75166 33936
rect 54 33120 75979 33656
rect 880 32840 75979 33120
rect 54 32304 75979 32840
rect 54 32024 75166 32304
rect 54 31488 75979 32024
rect 880 31208 75979 31488
rect 54 30672 75979 31208
rect 54 30392 75166 30672
rect 54 29856 75979 30392
rect 880 29576 75979 29856
rect 54 29040 75979 29576
rect 54 28760 75166 29040
rect 54 28224 75979 28760
rect 880 27944 75979 28224
rect 54 27408 75979 27944
rect 54 27128 75166 27408
rect 54 26592 75979 27128
rect 880 26312 75979 26592
rect 54 25776 75979 26312
rect 54 25496 75166 25776
rect 54 24960 75979 25496
rect 880 24680 75979 24960
rect 54 24144 75979 24680
rect 54 23864 75166 24144
rect 54 23328 75979 23864
rect 880 23048 75979 23328
rect 54 22512 75979 23048
rect 54 22232 75166 22512
rect 54 21696 75979 22232
rect 880 21416 75979 21696
rect 54 20880 75979 21416
rect 54 20600 75166 20880
rect 54 20064 75979 20600
rect 880 19784 75979 20064
rect 54 19248 75979 19784
rect 54 18968 75166 19248
rect 54 18432 75979 18968
rect 880 18152 75979 18432
rect 54 17616 75979 18152
rect 54 17336 75166 17616
rect 54 16800 75979 17336
rect 880 16520 75979 16800
rect 54 15984 75979 16520
rect 54 15704 75166 15984
rect 54 15168 75979 15704
rect 880 14888 75979 15168
rect 54 14352 75979 14888
rect 54 14072 75166 14352
rect 54 13536 75979 14072
rect 880 13256 75979 13536
rect 54 12720 75979 13256
rect 54 12440 75166 12720
rect 54 11904 75979 12440
rect 880 11624 75979 11904
rect 54 11088 75979 11624
rect 54 10808 75166 11088
rect 54 10272 75979 10808
rect 880 9992 75979 10272
rect 54 9456 75979 9992
rect 54 9176 75166 9456
rect 54 8640 75979 9176
rect 880 8360 75979 8640
rect 54 7824 75979 8360
rect 54 7544 75166 7824
rect 54 7008 75979 7544
rect 880 6728 75979 7008
rect 54 6192 75979 6728
rect 54 5912 75166 6192
rect 54 5376 75979 5912
rect 880 5096 75979 5376
rect 54 4560 75979 5096
rect 54 4280 75166 4560
rect 54 3744 75979 4280
rect 880 3464 75979 3744
rect 54 2928 75979 3464
rect 54 2648 75166 2928
rect 54 2112 75979 2648
rect 880 1832 75979 2112
rect 54 1803 75979 1832
<< metal4 >>
rect 4208 2128 4528 107760
rect 11888 2128 12208 107760
rect 19568 2128 19888 107760
rect 27248 2128 27568 107760
rect 34928 2128 35248 107760
rect 42608 2128 42928 107760
rect 50288 2128 50608 107760
rect 57968 2128 58288 107760
rect 65648 2128 65968 107760
rect 73328 2128 73648 107760
<< obsm4 >>
rect 59 2048 4128 107405
rect 4608 2048 11808 107405
rect 12288 2048 19488 107405
rect 19968 2048 27168 107405
rect 27648 2048 34848 107405
rect 35328 2048 42528 107405
rect 43008 2048 50208 107405
rect 50688 2048 57888 107405
rect 58368 2048 65568 107405
rect 66048 2048 73248 107405
rect 73728 2048 75749 107405
rect 59 1803 75749 2048
<< labels >>
rlabel metal4 s 11888 2128 12208 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27248 2128 27568 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 42608 2128 42928 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 57968 2128 58288 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 73328 2128 73648 107760 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 107760 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 1912 800 2032 6 debug_in
port 3 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 debug_mode
port 4 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 debug_oeb
port 5 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 debug_out
port 6 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 irq[0]
port 7 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 irq[1]
port 8 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 irq[2]
port 9 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 mask_rev_in[0]
port 10 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 mask_rev_in[10]
port 11 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 mask_rev_in[11]
port 12 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 mask_rev_in[12]
port 13 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 mask_rev_in[13]
port 14 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 mask_rev_in[14]
port 15 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 mask_rev_in[15]
port 16 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 mask_rev_in[16]
port 17 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 mask_rev_in[17]
port 18 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 mask_rev_in[18]
port 19 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 mask_rev_in[19]
port 20 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 mask_rev_in[1]
port 21 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 mask_rev_in[20]
port 22 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 mask_rev_in[21]
port 23 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 mask_rev_in[22]
port 24 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 mask_rev_in[23]
port 25 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 mask_rev_in[24]
port 26 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 mask_rev_in[25]
port 27 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 mask_rev_in[26]
port 28 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 mask_rev_in[27]
port 29 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 mask_rev_in[28]
port 30 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 mask_rev_in[29]
port 31 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 mask_rev_in[2]
port 32 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 mask_rev_in[30]
port 33 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 mask_rev_in[31]
port 34 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 mask_rev_in[3]
port 35 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 mask_rev_in[4]
port 36 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 mask_rev_in[5]
port 37 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 mask_rev_in[6]
port 38 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 mask_rev_in[7]
port 39 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 mask_rev_in[8]
port 40 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 mask_rev_in[9]
port 41 nsew signal input
rlabel metal3 s 75246 10888 76046 11008 6 mgmt_gpio_in[0]
port 42 nsew signal input
rlabel metal3 s 75246 59848 76046 59968 6 mgmt_gpio_in[10]
port 43 nsew signal input
rlabel metal3 s 75246 64744 76046 64864 6 mgmt_gpio_in[11]
port 44 nsew signal input
rlabel metal3 s 75246 69640 76046 69760 6 mgmt_gpio_in[12]
port 45 nsew signal input
rlabel metal3 s 75246 74536 76046 74656 6 mgmt_gpio_in[13]
port 46 nsew signal input
rlabel metal3 s 75246 79432 76046 79552 6 mgmt_gpio_in[14]
port 47 nsew signal input
rlabel metal3 s 75246 84328 76046 84448 6 mgmt_gpio_in[15]
port 48 nsew signal input
rlabel metal3 s 75246 89224 76046 89344 6 mgmt_gpio_in[16]
port 49 nsew signal input
rlabel metal3 s 75246 94120 76046 94240 6 mgmt_gpio_in[17]
port 50 nsew signal input
rlabel metal3 s 75246 99016 76046 99136 6 mgmt_gpio_in[18]
port 51 nsew signal input
rlabel metal3 s 75246 103912 76046 104032 6 mgmt_gpio_in[19]
port 52 nsew signal input
rlabel metal3 s 75246 15784 76046 15904 6 mgmt_gpio_in[1]
port 53 nsew signal input
rlabel metal2 s 43718 109390 43774 110190 6 mgmt_gpio_in[20]
port 54 nsew signal input
rlabel metal2 s 45374 109390 45430 110190 6 mgmt_gpio_in[21]
port 55 nsew signal input
rlabel metal2 s 47030 109390 47086 110190 6 mgmt_gpio_in[22]
port 56 nsew signal input
rlabel metal2 s 48686 109390 48742 110190 6 mgmt_gpio_in[23]
port 57 nsew signal input
rlabel metal2 s 50342 109390 50398 110190 6 mgmt_gpio_in[24]
port 58 nsew signal input
rlabel metal2 s 51998 109390 52054 110190 6 mgmt_gpio_in[25]
port 59 nsew signal input
rlabel metal2 s 53654 109390 53710 110190 6 mgmt_gpio_in[26]
port 60 nsew signal input
rlabel metal2 s 55310 109390 55366 110190 6 mgmt_gpio_in[27]
port 61 nsew signal input
rlabel metal2 s 56966 109390 57022 110190 6 mgmt_gpio_in[28]
port 62 nsew signal input
rlabel metal2 s 58622 109390 58678 110190 6 mgmt_gpio_in[29]
port 63 nsew signal input
rlabel metal3 s 75246 20680 76046 20800 6 mgmt_gpio_in[2]
port 64 nsew signal input
rlabel metal2 s 60278 109390 60334 110190 6 mgmt_gpio_in[30]
port 65 nsew signal input
rlabel metal2 s 61934 109390 61990 110190 6 mgmt_gpio_in[31]
port 66 nsew signal input
rlabel metal2 s 63590 109390 63646 110190 6 mgmt_gpio_in[32]
port 67 nsew signal input
rlabel metal2 s 65246 109390 65302 110190 6 mgmt_gpio_in[33]
port 68 nsew signal input
rlabel metal2 s 66902 109390 66958 110190 6 mgmt_gpio_in[34]
port 69 nsew signal input
rlabel metal2 s 68558 109390 68614 110190 6 mgmt_gpio_in[35]
port 70 nsew signal input
rlabel metal2 s 70214 109390 70270 110190 6 mgmt_gpio_in[36]
port 71 nsew signal input
rlabel metal2 s 71870 109390 71926 110190 6 mgmt_gpio_in[37]
port 72 nsew signal input
rlabel metal3 s 75246 25576 76046 25696 6 mgmt_gpio_in[3]
port 73 nsew signal input
rlabel metal3 s 75246 30472 76046 30592 6 mgmt_gpio_in[4]
port 74 nsew signal input
rlabel metal3 s 75246 35368 76046 35488 6 mgmt_gpio_in[5]
port 75 nsew signal input
rlabel metal3 s 75246 40264 76046 40384 6 mgmt_gpio_in[6]
port 76 nsew signal input
rlabel metal3 s 75246 45160 76046 45280 6 mgmt_gpio_in[7]
port 77 nsew signal input
rlabel metal3 s 75246 50056 76046 50176 6 mgmt_gpio_in[8]
port 78 nsew signal input
rlabel metal3 s 75246 54952 76046 55072 6 mgmt_gpio_in[9]
port 79 nsew signal input
rlabel metal3 s 75246 12520 76046 12640 6 mgmt_gpio_oeb[0]
port 80 nsew signal output
rlabel metal3 s 75246 61480 76046 61600 6 mgmt_gpio_oeb[10]
port 81 nsew signal output
rlabel metal3 s 75246 66376 76046 66496 6 mgmt_gpio_oeb[11]
port 82 nsew signal output
rlabel metal3 s 75246 71272 76046 71392 6 mgmt_gpio_oeb[12]
port 83 nsew signal output
rlabel metal3 s 75246 76168 76046 76288 6 mgmt_gpio_oeb[13]
port 84 nsew signal output
rlabel metal3 s 75246 81064 76046 81184 6 mgmt_gpio_oeb[14]
port 85 nsew signal output
rlabel metal3 s 75246 85960 76046 86080 6 mgmt_gpio_oeb[15]
port 86 nsew signal output
rlabel metal3 s 75246 90856 76046 90976 6 mgmt_gpio_oeb[16]
port 87 nsew signal output
rlabel metal3 s 75246 95752 76046 95872 6 mgmt_gpio_oeb[17]
port 88 nsew signal output
rlabel metal3 s 75246 100648 76046 100768 6 mgmt_gpio_oeb[18]
port 89 nsew signal output
rlabel metal3 s 75246 105544 76046 105664 6 mgmt_gpio_oeb[19]
port 90 nsew signal output
rlabel metal3 s 75246 17416 76046 17536 6 mgmt_gpio_oeb[1]
port 91 nsew signal output
rlabel metal2 s 44270 109390 44326 110190 6 mgmt_gpio_oeb[20]
port 92 nsew signal output
rlabel metal2 s 45926 109390 45982 110190 6 mgmt_gpio_oeb[21]
port 93 nsew signal output
rlabel metal2 s 47582 109390 47638 110190 6 mgmt_gpio_oeb[22]
port 94 nsew signal output
rlabel metal2 s 49238 109390 49294 110190 6 mgmt_gpio_oeb[23]
port 95 nsew signal output
rlabel metal2 s 50894 109390 50950 110190 6 mgmt_gpio_oeb[24]
port 96 nsew signal output
rlabel metal2 s 52550 109390 52606 110190 6 mgmt_gpio_oeb[25]
port 97 nsew signal output
rlabel metal2 s 54206 109390 54262 110190 6 mgmt_gpio_oeb[26]
port 98 nsew signal output
rlabel metal2 s 55862 109390 55918 110190 6 mgmt_gpio_oeb[27]
port 99 nsew signal output
rlabel metal2 s 57518 109390 57574 110190 6 mgmt_gpio_oeb[28]
port 100 nsew signal output
rlabel metal2 s 59174 109390 59230 110190 6 mgmt_gpio_oeb[29]
port 101 nsew signal output
rlabel metal3 s 75246 22312 76046 22432 6 mgmt_gpio_oeb[2]
port 102 nsew signal output
rlabel metal2 s 60830 109390 60886 110190 6 mgmt_gpio_oeb[30]
port 103 nsew signal output
rlabel metal2 s 62486 109390 62542 110190 6 mgmt_gpio_oeb[31]
port 104 nsew signal output
rlabel metal2 s 64142 109390 64198 110190 6 mgmt_gpio_oeb[32]
port 105 nsew signal output
rlabel metal2 s 65798 109390 65854 110190 6 mgmt_gpio_oeb[33]
port 106 nsew signal output
rlabel metal2 s 67454 109390 67510 110190 6 mgmt_gpio_oeb[34]
port 107 nsew signal output
rlabel metal2 s 69110 109390 69166 110190 6 mgmt_gpio_oeb[35]
port 108 nsew signal output
rlabel metal2 s 70766 109390 70822 110190 6 mgmt_gpio_oeb[36]
port 109 nsew signal output
rlabel metal2 s 72422 109390 72478 110190 6 mgmt_gpio_oeb[37]
port 110 nsew signal output
rlabel metal3 s 75246 27208 76046 27328 6 mgmt_gpio_oeb[3]
port 111 nsew signal output
rlabel metal3 s 75246 32104 76046 32224 6 mgmt_gpio_oeb[4]
port 112 nsew signal output
rlabel metal3 s 75246 37000 76046 37120 6 mgmt_gpio_oeb[5]
port 113 nsew signal output
rlabel metal3 s 75246 41896 76046 42016 6 mgmt_gpio_oeb[6]
port 114 nsew signal output
rlabel metal3 s 75246 46792 76046 46912 6 mgmt_gpio_oeb[7]
port 115 nsew signal output
rlabel metal3 s 75246 51688 76046 51808 6 mgmt_gpio_oeb[8]
port 116 nsew signal output
rlabel metal3 s 75246 56584 76046 56704 6 mgmt_gpio_oeb[9]
port 117 nsew signal output
rlabel metal3 s 75246 14152 76046 14272 6 mgmt_gpio_out[0]
port 118 nsew signal output
rlabel metal3 s 75246 63112 76046 63232 6 mgmt_gpio_out[10]
port 119 nsew signal output
rlabel metal3 s 75246 68008 76046 68128 6 mgmt_gpio_out[11]
port 120 nsew signal output
rlabel metal3 s 75246 72904 76046 73024 6 mgmt_gpio_out[12]
port 121 nsew signal output
rlabel metal3 s 75246 77800 76046 77920 6 mgmt_gpio_out[13]
port 122 nsew signal output
rlabel metal3 s 75246 82696 76046 82816 6 mgmt_gpio_out[14]
port 123 nsew signal output
rlabel metal3 s 75246 87592 76046 87712 6 mgmt_gpio_out[15]
port 124 nsew signal output
rlabel metal3 s 75246 92488 76046 92608 6 mgmt_gpio_out[16]
port 125 nsew signal output
rlabel metal3 s 75246 97384 76046 97504 6 mgmt_gpio_out[17]
port 126 nsew signal output
rlabel metal3 s 75246 102280 76046 102400 6 mgmt_gpio_out[18]
port 127 nsew signal output
rlabel metal3 s 75246 107176 76046 107296 6 mgmt_gpio_out[19]
port 128 nsew signal output
rlabel metal3 s 75246 19048 76046 19168 6 mgmt_gpio_out[1]
port 129 nsew signal output
rlabel metal2 s 44822 109390 44878 110190 6 mgmt_gpio_out[20]
port 130 nsew signal output
rlabel metal2 s 46478 109390 46534 110190 6 mgmt_gpio_out[21]
port 131 nsew signal output
rlabel metal2 s 48134 109390 48190 110190 6 mgmt_gpio_out[22]
port 132 nsew signal output
rlabel metal2 s 49790 109390 49846 110190 6 mgmt_gpio_out[23]
port 133 nsew signal output
rlabel metal2 s 51446 109390 51502 110190 6 mgmt_gpio_out[24]
port 134 nsew signal output
rlabel metal2 s 53102 109390 53158 110190 6 mgmt_gpio_out[25]
port 135 nsew signal output
rlabel metal2 s 54758 109390 54814 110190 6 mgmt_gpio_out[26]
port 136 nsew signal output
rlabel metal2 s 56414 109390 56470 110190 6 mgmt_gpio_out[27]
port 137 nsew signal output
rlabel metal2 s 58070 109390 58126 110190 6 mgmt_gpio_out[28]
port 138 nsew signal output
rlabel metal2 s 59726 109390 59782 110190 6 mgmt_gpio_out[29]
port 139 nsew signal output
rlabel metal3 s 75246 23944 76046 24064 6 mgmt_gpio_out[2]
port 140 nsew signal output
rlabel metal2 s 61382 109390 61438 110190 6 mgmt_gpio_out[30]
port 141 nsew signal output
rlabel metal2 s 63038 109390 63094 110190 6 mgmt_gpio_out[31]
port 142 nsew signal output
rlabel metal2 s 64694 109390 64750 110190 6 mgmt_gpio_out[32]
port 143 nsew signal output
rlabel metal2 s 66350 109390 66406 110190 6 mgmt_gpio_out[33]
port 144 nsew signal output
rlabel metal2 s 68006 109390 68062 110190 6 mgmt_gpio_out[34]
port 145 nsew signal output
rlabel metal2 s 69662 109390 69718 110190 6 mgmt_gpio_out[35]
port 146 nsew signal output
rlabel metal2 s 71318 109390 71374 110190 6 mgmt_gpio_out[36]
port 147 nsew signal output
rlabel metal2 s 72974 109390 73030 110190 6 mgmt_gpio_out[37]
port 148 nsew signal output
rlabel metal3 s 75246 28840 76046 28960 6 mgmt_gpio_out[3]
port 149 nsew signal output
rlabel metal3 s 75246 33736 76046 33856 6 mgmt_gpio_out[4]
port 150 nsew signal output
rlabel metal3 s 75246 38632 76046 38752 6 mgmt_gpio_out[5]
port 151 nsew signal output
rlabel metal3 s 75246 43528 76046 43648 6 mgmt_gpio_out[6]
port 152 nsew signal output
rlabel metal3 s 75246 48424 76046 48544 6 mgmt_gpio_out[7]
port 153 nsew signal output
rlabel metal3 s 75246 53320 76046 53440 6 mgmt_gpio_out[8]
port 154 nsew signal output
rlabel metal3 s 75246 58216 76046 58336 6 mgmt_gpio_out[9]
port 155 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 pad_flash_clk
port 156 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 pad_flash_clk_oeb
port 157 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 pad_flash_csb
port 158 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 pad_flash_csb_oeb
port 159 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 pad_flash_io0_di
port 160 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 pad_flash_io0_do
port 161 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 pad_flash_io0_ieb
port 162 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 pad_flash_io0_oeb
port 163 nsew signal output
rlabel metal2 s 10690 0 10746 800 6 pad_flash_io1_di
port 164 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 pad_flash_io1_do
port 165 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 pad_flash_io1_ieb
port 166 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 pad_flash_io1_oeb
port 167 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 pll90_sel[0]
port 168 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 pll90_sel[1]
port 169 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 pll90_sel[2]
port 170 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 pll_bypass
port 171 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 pll_dco_ena
port 172 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 pll_div[0]
port 173 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 pll_div[1]
port 174 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 pll_div[2]
port 175 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 pll_div[3]
port 176 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 pll_div[4]
port 177 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 pll_ena
port 178 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 pll_sel[0]
port 179 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 pll_sel[1]
port 180 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 pll_sel[2]
port 181 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 pll_trim[0]
port 182 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 pll_trim[10]
port 183 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 pll_trim[11]
port 184 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 pll_trim[12]
port 185 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 pll_trim[13]
port 186 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 pll_trim[14]
port 187 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 pll_trim[15]
port 188 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 pll_trim[16]
port 189 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 pll_trim[17]
port 190 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 pll_trim[18]
port 191 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 pll_trim[19]
port 192 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 pll_trim[1]
port 193 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 pll_trim[20]
port 194 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 pll_trim[21]
port 195 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 pll_trim[22]
port 196 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 pll_trim[23]
port 197 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 pll_trim[24]
port 198 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 pll_trim[25]
port 199 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 pll_trim[2]
port 200 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 pll_trim[3]
port 201 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 pll_trim[4]
port 202 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 pll_trim[5]
port 203 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 pll_trim[6]
port 204 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 pll_trim[7]
port 205 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 pll_trim[8]
port 206 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 pll_trim[9]
port 207 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 porb
port 208 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 pwr_ctrl_out[0]
port 209 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 pwr_ctrl_out[1]
port 210 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 pwr_ctrl_out[2]
port 211 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 pwr_ctrl_out[3]
port 212 nsew signal output
rlabel metal3 s 0 26392 800 26512 6 qspi_enabled
port 213 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 reset
port 214 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 ser_rx
port 215 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 ser_tx
port 216 nsew signal input
rlabel metal3 s 75246 2728 76046 2848 6 serial_clock
port 217 nsew signal output
rlabel metal3 s 75246 7624 76046 7744 6 serial_data_1
port 218 nsew signal output
rlabel metal3 s 75246 9256 76046 9376 6 serial_data_2
port 219 nsew signal output
rlabel metal3 s 75246 5992 76046 6112 6 serial_load
port 220 nsew signal output
rlabel metal3 s 75246 4360 76046 4480 6 serial_resetn
port 221 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 spi_csb
port 222 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 spi_enabled
port 223 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 spi_sck
port 224 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 spi_sdi
port 225 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 spi_sdo
port 226 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 spi_sdoenb
port 227 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 spimemio_flash_clk
port 228 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 spimemio_flash_csb
port 229 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 spimemio_flash_io0_di
port 230 nsew signal output
rlabel metal3 s 0 91672 800 91792 6 spimemio_flash_io0_do
port 231 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 spimemio_flash_io0_oeb
port 232 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 spimemio_flash_io1_di
port 233 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 spimemio_flash_io1_do
port 234 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 spimemio_flash_io1_oeb
port 235 nsew signal input
rlabel metal3 s 0 99832 800 99952 6 spimemio_flash_io2_di
port 236 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 spimemio_flash_io2_do
port 237 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 spimemio_flash_io2_oeb
port 238 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 spimemio_flash_io3_di
port 239 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 spimemio_flash_io3_do
port 240 nsew signal input
rlabel metal3 s 0 107992 800 108112 6 spimemio_flash_io3_oeb
port 241 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 trap
port 242 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 uart_enabled
port 243 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 user_clock
port 244 nsew signal input
rlabel metal2 s 41510 109390 41566 110190 6 usr1_vcc_pwrgood
port 245 nsew signal input
rlabel metal2 s 42614 109390 42670 110190 6 usr1_vdd_pwrgood
port 246 nsew signal input
rlabel metal2 s 42062 109390 42118 110190 6 usr2_vcc_pwrgood
port 247 nsew signal input
rlabel metal2 s 43166 109390 43222 110190 6 usr2_vdd_pwrgood
port 248 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 wb_ack_o
port 249 nsew signal output
rlabel metal2 s 2870 109390 2926 110190 6 wb_adr_i[0]
port 250 nsew signal input
rlabel metal2 s 8390 109390 8446 110190 6 wb_adr_i[10]
port 251 nsew signal input
rlabel metal2 s 8942 109390 8998 110190 6 wb_adr_i[11]
port 252 nsew signal input
rlabel metal2 s 9494 109390 9550 110190 6 wb_adr_i[12]
port 253 nsew signal input
rlabel metal2 s 10046 109390 10102 110190 6 wb_adr_i[13]
port 254 nsew signal input
rlabel metal2 s 10598 109390 10654 110190 6 wb_adr_i[14]
port 255 nsew signal input
rlabel metal2 s 11150 109390 11206 110190 6 wb_adr_i[15]
port 256 nsew signal input
rlabel metal2 s 11702 109390 11758 110190 6 wb_adr_i[16]
port 257 nsew signal input
rlabel metal2 s 12254 109390 12310 110190 6 wb_adr_i[17]
port 258 nsew signal input
rlabel metal2 s 12806 109390 12862 110190 6 wb_adr_i[18]
port 259 nsew signal input
rlabel metal2 s 13358 109390 13414 110190 6 wb_adr_i[19]
port 260 nsew signal input
rlabel metal2 s 3422 109390 3478 110190 6 wb_adr_i[1]
port 261 nsew signal input
rlabel metal2 s 13910 109390 13966 110190 6 wb_adr_i[20]
port 262 nsew signal input
rlabel metal2 s 14462 109390 14518 110190 6 wb_adr_i[21]
port 263 nsew signal input
rlabel metal2 s 15014 109390 15070 110190 6 wb_adr_i[22]
port 264 nsew signal input
rlabel metal2 s 15566 109390 15622 110190 6 wb_adr_i[23]
port 265 nsew signal input
rlabel metal2 s 16118 109390 16174 110190 6 wb_adr_i[24]
port 266 nsew signal input
rlabel metal2 s 16670 109390 16726 110190 6 wb_adr_i[25]
port 267 nsew signal input
rlabel metal2 s 17222 109390 17278 110190 6 wb_adr_i[26]
port 268 nsew signal input
rlabel metal2 s 17774 109390 17830 110190 6 wb_adr_i[27]
port 269 nsew signal input
rlabel metal2 s 18326 109390 18382 110190 6 wb_adr_i[28]
port 270 nsew signal input
rlabel metal2 s 18878 109390 18934 110190 6 wb_adr_i[29]
port 271 nsew signal input
rlabel metal2 s 3974 109390 4030 110190 6 wb_adr_i[2]
port 272 nsew signal input
rlabel metal2 s 19430 109390 19486 110190 6 wb_adr_i[30]
port 273 nsew signal input
rlabel metal2 s 19982 109390 20038 110190 6 wb_adr_i[31]
port 274 nsew signal input
rlabel metal2 s 4526 109390 4582 110190 6 wb_adr_i[3]
port 275 nsew signal input
rlabel metal2 s 5078 109390 5134 110190 6 wb_adr_i[4]
port 276 nsew signal input
rlabel metal2 s 5630 109390 5686 110190 6 wb_adr_i[5]
port 277 nsew signal input
rlabel metal2 s 6182 109390 6238 110190 6 wb_adr_i[6]
port 278 nsew signal input
rlabel metal2 s 6734 109390 6790 110190 6 wb_adr_i[7]
port 279 nsew signal input
rlabel metal2 s 7286 109390 7342 110190 6 wb_adr_i[8]
port 280 nsew signal input
rlabel metal2 s 7838 109390 7894 110190 6 wb_adr_i[9]
port 281 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wb_clk_i
port 282 nsew signal input
rlabel metal2 s 40958 109390 41014 110190 6 wb_cyc_i
port 283 nsew signal input
rlabel metal2 s 20534 109390 20590 110190 6 wb_dat_i[0]
port 284 nsew signal input
rlabel metal2 s 26054 109390 26110 110190 6 wb_dat_i[10]
port 285 nsew signal input
rlabel metal2 s 26606 109390 26662 110190 6 wb_dat_i[11]
port 286 nsew signal input
rlabel metal2 s 27158 109390 27214 110190 6 wb_dat_i[12]
port 287 nsew signal input
rlabel metal2 s 27710 109390 27766 110190 6 wb_dat_i[13]
port 288 nsew signal input
rlabel metal2 s 28262 109390 28318 110190 6 wb_dat_i[14]
port 289 nsew signal input
rlabel metal2 s 28814 109390 28870 110190 6 wb_dat_i[15]
port 290 nsew signal input
rlabel metal2 s 29366 109390 29422 110190 6 wb_dat_i[16]
port 291 nsew signal input
rlabel metal2 s 29918 109390 29974 110190 6 wb_dat_i[17]
port 292 nsew signal input
rlabel metal2 s 30470 109390 30526 110190 6 wb_dat_i[18]
port 293 nsew signal input
rlabel metal2 s 31022 109390 31078 110190 6 wb_dat_i[19]
port 294 nsew signal input
rlabel metal2 s 21086 109390 21142 110190 6 wb_dat_i[1]
port 295 nsew signal input
rlabel metal2 s 31574 109390 31630 110190 6 wb_dat_i[20]
port 296 nsew signal input
rlabel metal2 s 32126 109390 32182 110190 6 wb_dat_i[21]
port 297 nsew signal input
rlabel metal2 s 32678 109390 32734 110190 6 wb_dat_i[22]
port 298 nsew signal input
rlabel metal2 s 33230 109390 33286 110190 6 wb_dat_i[23]
port 299 nsew signal input
rlabel metal2 s 33782 109390 33838 110190 6 wb_dat_i[24]
port 300 nsew signal input
rlabel metal2 s 34334 109390 34390 110190 6 wb_dat_i[25]
port 301 nsew signal input
rlabel metal2 s 34886 109390 34942 110190 6 wb_dat_i[26]
port 302 nsew signal input
rlabel metal2 s 35438 109390 35494 110190 6 wb_dat_i[27]
port 303 nsew signal input
rlabel metal2 s 35990 109390 36046 110190 6 wb_dat_i[28]
port 304 nsew signal input
rlabel metal2 s 36542 109390 36598 110190 6 wb_dat_i[29]
port 305 nsew signal input
rlabel metal2 s 21638 109390 21694 110190 6 wb_dat_i[2]
port 306 nsew signal input
rlabel metal2 s 37094 109390 37150 110190 6 wb_dat_i[30]
port 307 nsew signal input
rlabel metal2 s 37646 109390 37702 110190 6 wb_dat_i[31]
port 308 nsew signal input
rlabel metal2 s 22190 109390 22246 110190 6 wb_dat_i[3]
port 309 nsew signal input
rlabel metal2 s 22742 109390 22798 110190 6 wb_dat_i[4]
port 310 nsew signal input
rlabel metal2 s 23294 109390 23350 110190 6 wb_dat_i[5]
port 311 nsew signal input
rlabel metal2 s 23846 109390 23902 110190 6 wb_dat_i[6]
port 312 nsew signal input
rlabel metal2 s 24398 109390 24454 110190 6 wb_dat_i[7]
port 313 nsew signal input
rlabel metal2 s 24950 109390 25006 110190 6 wb_dat_i[8]
port 314 nsew signal input
rlabel metal2 s 25502 109390 25558 110190 6 wb_dat_i[9]
port 315 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 wb_dat_o[0]
port 316 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 wb_dat_o[10]
port 317 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 wb_dat_o[11]
port 318 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 wb_dat_o[12]
port 319 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 wb_dat_o[13]
port 320 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 wb_dat_o[14]
port 321 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 wb_dat_o[15]
port 322 nsew signal output
rlabel metal3 s 0 60664 800 60784 6 wb_dat_o[16]
port 323 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 wb_dat_o[17]
port 324 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 wb_dat_o[18]
port 325 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 wb_dat_o[19]
port 326 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 wb_dat_o[1]
port 327 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 wb_dat_o[20]
port 328 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 wb_dat_o[21]
port 329 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 wb_dat_o[22]
port 330 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 wb_dat_o[23]
port 331 nsew signal output
rlabel metal3 s 0 73720 800 73840 6 wb_dat_o[24]
port 332 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 wb_dat_o[25]
port 333 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 wb_dat_o[26]
port 334 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 wb_dat_o[27]
port 335 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 wb_dat_o[28]
port 336 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 wb_dat_o[29]
port 337 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 wb_dat_o[2]
port 338 nsew signal output
rlabel metal3 s 0 83512 800 83632 6 wb_dat_o[30]
port 339 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 wb_dat_o[31]
port 340 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 wb_dat_o[3]
port 341 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 wb_dat_o[4]
port 342 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 wb_dat_o[5]
port 343 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 wb_dat_o[6]
port 344 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 wb_dat_o[7]
port 345 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 wb_dat_o[8]
port 346 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 wb_dat_o[9]
port 347 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 wb_rstn_i
port 348 nsew signal input
rlabel metal2 s 38198 109390 38254 110190 6 wb_sel_i[0]
port 349 nsew signal input
rlabel metal2 s 38750 109390 38806 110190 6 wb_sel_i[1]
port 350 nsew signal input
rlabel metal2 s 39302 109390 39358 110190 6 wb_sel_i[2]
port 351 nsew signal input
rlabel metal2 s 39854 109390 39910 110190 6 wb_sel_i[3]
port 352 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 wb_stb_i
port 353 nsew signal input
rlabel metal2 s 40406 109390 40462 110190 6 wb_we_i
port 354 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 76046 110190
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27242318
string GDS_FILE /home/hosni/caravel_sky130/caravel/openlane/housekeeping/runs/23_02_08_05_38/results/signoff/housekeeping.magic.gds
string GDS_START 1528686
<< end >>

