* trimmed fd_pr

.subckt  sky130_fd_pr__cap_mim_m3_1 c0 c1 w=1 l=1 mf=1
.ends

.subckt  sky130_fd_pr__cap_mim_m3_2 c0 c1 w=1 l=1 mf=1
.ends

.subckt  sky130_fd_pr__cap_var_hvt c0 c1 b w=5 l=0.5 vm=1
.ends

.subckt  sky130_fd_pr__cap_var_lvt c0 c1 b w=5 l=0.5 vm=1
.ends

.subckt  sky130_fd_pr__cap_vpp_01p8x01p8_m1m2_noshield c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_02p4x04p6_m1m2_noshield c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_02p7x06p1_m1m2m3m4_shieldl1_fingercap c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_02p7x11p1_m1m2m3m4_shieldl1_fingercap c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_02p7x21p1_m1m2m3m4_shieldl1_fingercap c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_02p7x41p1_m1m2m3m4_shieldl1_fingercap c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_02p9x06p1_m1m2m3m4_shieldl1_fingercap2 c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3 c0 c1 b m3
.ends

.subckt  sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield_o1 c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3 c0 c1 b m3
.ends

.subckt  sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o1nhv c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o1phv c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o2 c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1 c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1 c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1m5_floatm4 c0 c1 b m5
.ends

.subckt sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1m5_floatm4_top C0 C1 M5 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_05p9x05p9_m1m2m3m4_shieldl1_wafflecap c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4 c0 c1 b m4
.ends

.subckt sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4_top C0 C1 M4 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_06p8x06p1_m1m2m3_shieldl1m4 c0 c1 b m4
.ends

.subckt sky130_fd_pr__cap_vpp_06p8x06p1_m1m2m3_shieldl1m4_top C0 C1 M4 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o1 c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3 c0 c1 b m3
.ends

.subckt  sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_shieldl1 c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1 c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4 c0 c1 b m5
.ends

.subckt sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4_top C0 C1 M5 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_11p3x11p3_m1m2m3m4_shieldl1_wafflecap c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhv c0 c1 b m5
.ends

.subckt  sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhv__base d g s b
.ends

.subckt sky130_fd_pr__cap_vpp_11p3x11p8_l1m1m2m3m4_shieldm5_nhvtop C0 M5 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_noshield c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3 c0 c1 b m3
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4 c0 c1 b m4
.ends

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4_top C0 C1 M4 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4 c0 c1 b m4
.ends

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top C0 C1 M4 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5 c0 c1 b m5
.ends

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5_top C0 C1 M5 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5 c0 c1 b m5
.ends

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_top C0 C1 M5 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x c0 c1 b m5
.ends

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x6 C0 C1 M5A SUB
.ends

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x7 C0 C1 M5A SUB
.ends

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x8 C0 C1 M5A SUB
.ends

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_x9 C0 C1 M5A SUB
.ends

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5_xtop C0 C1 M5 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1 c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1 c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4 c0 c1 b m5
.ends

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1m5_floatm4_top C0 C1 M5 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5 c0 c1 b m5
.ends

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_top C0 C1 M5 SUB
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldm5 c0 c1 b m5
.ends

.subckt  sky130_fd_pr__cap_vpp_11p5x11p7_m1m4_noshield c0 c1 b
.ends

.subckt  sky130_fd_pr__cap_vpp_44p7x23p1_pol1m1m2m3m4m5_noshield c0 c1 b mf=1
.ends

.subckt  sky130_fd_pr__esd_nfet_01v8 d g s b
.ends

.subckt  sky130_fd_pr__esd_nfet_05v0_nvt d g s b
.ends

.subckt  sky130_fd_pr__esd_nfet_g5v0d10v5 d g s b
.ends

.subckt  sky130_fd_pr__esd_pfet_g5v0d10v5 d g s b
.ends

.subckt  sky130_fd_pr__esd_rf_diode_pd2nw_11v0_100 c0 c1
.ends

.subckt  sky130_fd_pr__esd_rf_diode_pd2nw_11v0_200 c0 c1
.ends

.subckt  sky130_fd_pr__esd_rf_diode_pd2nw_11v0_300 c0 c1
.ends

.subckt  sky130_fd_pr__esd_rf_diode_pw2nd_11v0_100 c0 c1
.ends

.subckt  sky130_fd_pr__esd_rf_diode_pw2nd_11v0_100__parasitic__diode_pw2dn c0 c1
.ends

.subckt  sky130_fd_pr__esd_rf_diode_pw2nd_11v0_200 c0 c1
.ends

.subckt  sky130_fd_pr__esd_rf_diode_pw2nd_11v0_200__parasitic__diode_pw2dn c0 c1
.ends

.subckt  sky130_fd_pr__esd_rf_diode_pw2nd_11v0_300 c0 c1
.ends

.subckt  sky130_fd_pr__esd_rf_diode_pw2nd_11v0_300__parasitic__diode_pw2dn c0 c1
.ends

.subckt  sky130_fd_pr__ind_03_90 a b ct sub
.ends

.subckt  sky130_fd_pr__ind_05_125 a b ct sub
.ends

.subckt  sky130_fd_pr__ind_05_220 a b ct sub
.ends

.subckt  sky130_fd_pr__nfet_01v8 d g s b
.ends

.subckt  sky130_fd_pr__nfet_01v8_lvt d g s b
.ends

.subckt  sky130_fd_pr__nfet_03v3_nvt d g s b
.ends

.subckt  sky130_fd_pr__nfet_05v0_nvt d g s b
.ends

.subckt  sky130_fd_pr__nfet_20v0 d g s b  w=60u l=2u m=1 t=30
.ends

.subckt  sky130_fd_pr__nfet_20v0_iso d g s b sub  w=60u l=2u m=1 t=30
.ends

.subckt  sky130_fd_pr__nfet_20v0_nvt d g s b  w=60u l=2u m=1 t=30
.ends

.subckt  sky130_fd_pr__nfet_20v0_nvt_iso d g s b sub  w=60u l=2u m=1 t=30
.ends

.subckt  sky130_fd_pr__nfet_20v0_reverse_iso d g s b sub w=60u l=2u m=1 t=30
.ends

.subckt  sky130_fd_pr__nfet_20v0_zvt d g s b  w=60u l=2u m=1 t=30
.ends

.subckt  sky130_fd_pr__nfet_g5v0d10v5 d g s b
.ends

.subckt  sky130_fd_pr__nfet_g5v0d16v0__base d g s b
.ends

.subckt  sky130_fd_pr__nfet_g5v0d16v0 d g s b  w=5.0 l=0.7 nf=1 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0 delvto=0 m=1 sa=0.28 sb=2.41 sd=0 mult=1
.ends

.subckt  sky130_fd_pr__npn_05v5_W1p00L1p00 c b e s
.ends

.subckt  sky130_fd_pr__npn_05v5_W1p00L2p00 c b e s
.ends

.subckt  sky130_fd_pr__npn_11v0_W1p00L1p00 c b e s
.ends

.subckt  sky130_fd_pr__pfet_01v8 d g s b
.ends

.subckt  sky130_fd_pr__pfet_01v8_hvt d g s b
.ends

.subckt  sky130_fd_pr__pfet_01v8_lvt d g s b
.ends

.subckt  sky130_fd_pr__pfet_01v8_mvt d g s b
.ends

.subckt  sky130_fd_pr__pfet_20v0 d g s b  w=50u l=2u m=1 t=30 ad=0 as=0 pd=0 ps=0 nrd=0 nrs=0
.ends

.subckt  sky130_fd_pr__pfet_g5v0d10v5 d g s b
.ends

.subckt  sky130_fd_pr__pfet_g5v0d16v0__base d g s b
.ends

.subckt  sky130_fd_pr__pfet_g5v0d16v0 d g s b  w=5.0 l=0.66 nf=1 ad=0 as=0 pd=0 ps=0.0 m=1 nrd=0 nrs=0 sa=0.28 sb=1.19 sd=0 mult=1
.ends

.subckt  sky130_fd_pr__pnp_05v5_W0p68L0p68 Collector Base Emitter
.ends

.subckt  sky130_fd_pr__pnp_05v5_W3p40L3p40 Collector Base Emitter
.ends

.subckt  sky130_fd_pr__res_generic_nd t1 t2 b
.ends

.subckt  sky130_fd_pr__res_generic_pd t1 t2 b
.ends

.subckt  sky130_fd_pr__res_high_po r0 r1 b
.ends

.subckt  sky130_fd_pr__res_high_po_0p35 r0 r1 b
.ends

.subckt  sky130_fd_pr__res_high_po_0p69 r0 r1 b
.ends

.subckt  sky130_fd_pr__res_high_po_1p41 r0 r1 b
.ends

.subckt  sky130_fd_pr__res_high_po_2p85 r0 r1 b
.ends

.subckt  sky130_fd_pr__res_high_po_5p73 r0 r1 b
.ends

.subckt  sky130_fd_pr__res_iso_pw r0 r1 b
.ends

.subckt  sky130_fd_pr__res_xhigh_po r0 r1 sub
.ends

.subckt  sky130_fd_pr__res_xhigh_po_0p35 r0 r1 b
.ends

.subckt  sky130_fd_pr__res_xhigh_po_0p69 r0 r1 b
.ends

.subckt  sky130_fd_pr__res_xhigh_po_1p41 r0 r1 b
.ends

.subckt  sky130_fd_pr__res_xhigh_po_2p85 r0 r1 b
.ends

.subckt  sky130_fd_pr__res_xhigh_po_5p73 r0 r1 b
.ends

.subckt  sky130_fd_pr__res_xhigh_po__base r1 r2 b
.ends

.subckt sky130_fd_pr__rf_aura_blocking B_P D_N2 D_P D_P2 G G_N2 G_P G_P2 NWELL S S_N2
.ends

.subckt sky130_fd_pr__rf_aura_drc_flag_check B_P NWELL VGND
.ends

.subckt sky130_fd_pr__rf_aura_lvs_drc B_P D_P G G_P NWELL S S_P VGND VPWR
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02W1p65L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04W1p65L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02W3p00L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04W3p00L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02W5p00L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p25 d g s b
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM02W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM04W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM04W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02W3p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM02W5p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04W3p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_bM04W5p00 d g s b
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_hcM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_hcM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p84L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_aF04W3p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_aF02W3p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_aF08W0p84L0p15 d g s b
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aF02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p42L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aF04W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aF06W0p42L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aF06W0p84L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aF06W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aF06W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aF08W0p42L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aF08W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM02W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM02W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM02W5p00L0p25 GATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM04W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM04W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_aM04W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_bM02 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_bM04 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p25 d g s b
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM02W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM04W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM04W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_bM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM02W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM02W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM02W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM02W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM02W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM02W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM02W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM04W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM04W1p65L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM04W1p65L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM04W3p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM04W3p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM04W5p00L0p18 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cM04W5p00L0p25 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_mcM04W3p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_mcM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_20v0_nvt_aup D PSUB S
.ends

.subckt sky130_fd_pr__rf_nfet_20v0_nvt_withptap D G PSUB S
.ends

.subckt sky130_fd_pr__rf_nfet_20v0_zvt_withptap D PSUB S
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W3p00L0p50 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W3p00L0p50 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00L0p50 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00L0p50 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00L0p50 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00L0p50 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00L0p50 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W3p00L0p50 d g s b
.ends

.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W3p00L0p50 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W5p00L0p50 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_aM04W7p00L0p50 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W3p00L0p50 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W5p00L0p50 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_aM10W7p00L0p50 DRAIN GATE SOURCE SUBSTRATE
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM02W5p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W5p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM04W7p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W5p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_nfet_g5v0d10v5_bM10W7p00 d g s b
.ends

.subckt sky130_fd_pr__rf_npn_11v0_W1p00L1p00 E B C
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15 d g s b
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aF02W2p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aF04W0p84L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aF04W2p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aF04W3p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aF06W0p84L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aF06W1p68L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aF06W2p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aF06W3p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aF08W0p84L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aF08W1p68L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p18 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM02W1p65L0p25 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p18 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM02W3p00L0p25 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p18 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM02W5p00L0p25 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p18 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM04W1p65L0p25 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p18 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM04W3p00L0p25 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p18 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p25 BULK DRAIN GATE SOURCE
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W3p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W5p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W3p00 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W5p00 d g s b
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_hcM04W3p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_hcM04W5p00L0p15 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_lvt_aM02W3p00L0p35 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_lvt_aM02W3p00L0p50 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_lvt_aM02W5p00L0p35 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_lvt_aM02W5p00L0p50 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_lvt_aM04W3p00L0p35 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_lvt_aM04W3p00L0p50 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p35 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_lvt_aM04W5p00L0p50 BULK DRAIN GATE SOURCE
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_mcM04W3p00L0p15 DRAIN GATE SOURCE BULK
.ends

.subckt sky130_fd_pr__rf_pfet_01v8_mcM04W5p00L0p15 DRAIN GATE SOURCE Bulk
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_mvt_aF02W1p68L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_mvt_aF02W0p84L0p15 d g s b
.ends

.subckt  sky130_fd_pr__rf_pfet_01v8_mvt_aF04W1p68L0p15 d g s b
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W0p68L0p68 Base Collector Emitter
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base
.ends

.subckt  sky130_fd_pr__special_nfet_latch d g s b
.ends

.subckt  sky130_fd_pr__special_nfet_pass d g s b
.ends

.subckt  sky130_fd_pr__special_nfet_pass_flash d g s b
.ends

.subckt  sky130_fd_pr__special_nfet_pass_lvt d g s b
.ends

.subckt  sky130_fd_pr__special_pfet_pass d g s b
.ends

