magic
tech sky130A
magscale 1 2
timestamp 1539367940
<< checkpaint >>
rect -4476 -9457 636864 956856
<< metal3 >>
rect 533387 954354 538193 955596
rect 533387 952770 533467 954354
rect 538091 952770 538193 954354
rect 533387 952680 538193 952770
rect 543368 954354 548174 955596
rect 543368 952770 543448 954354
rect 548072 952770 548174 954354
rect 543368 952680 548174 952770
rect -3216 884758 1182 884840
rect -3216 880134 -1777 884758
rect 1087 880134 1182 884758
rect -3216 880051 1182 880134
rect 631206 880318 635604 880400
rect -2200 879648 1182 879730
rect -2200 875184 -1777 879648
rect 1087 875184 1182 879648
rect 631206 875694 631301 880318
rect 634165 875694 635604 880318
rect 631206 875611 635604 875694
rect -2200 875120 1182 875184
rect 631206 875208 635204 875290
rect -3216 874718 1182 874800
rect -3216 870094 -1777 874718
rect 1087 870094 1182 874718
rect 631206 870744 631301 875208
rect 634165 870744 635204 875208
rect 631206 870669 635204 870744
rect -3216 870011 1182 870094
rect 631206 870267 635604 870349
rect 631206 865643 631301 870267
rect 634165 865643 635604 870267
rect 631206 865560 635604 865643
rect -3216 800276 1182 800358
rect -3216 795652 -1777 800276
rect 1087 795652 1182 800276
rect -3216 795569 1182 795652
rect 631206 791119 635604 791201
rect -3216 790297 1182 790379
rect -3216 785673 -1777 790297
rect 1087 785673 1182 790297
rect 631206 786495 631301 791119
rect 634165 786495 635604 791119
rect 631206 786412 635604 786495
rect -3216 785590 1182 785673
rect 631206 781136 635604 781218
rect 631206 776512 631301 781136
rect 634165 776512 635604 781136
rect 631206 776429 635604 776512
rect 631206 476519 635604 476601
rect 631206 471895 631301 476519
rect 634165 471895 635604 476519
rect 631206 471812 635604 471895
rect 631206 466536 635604 466618
rect 631206 461912 631301 466536
rect 634165 461912 635604 466536
rect 631206 461829 635604 461912
rect -3216 455676 1182 455758
rect -3216 451052 -1777 455676
rect 1087 451052 1182 455676
rect -3216 450969 1182 451052
rect -3216 445697 1182 445779
rect -3216 441073 -1777 445697
rect 1087 441073 1182 445697
rect -3216 440990 1182 441073
rect 631206 432518 635604 432600
rect 631206 427894 631301 432518
rect 634165 427894 635604 432518
rect 631206 427811 635604 427894
rect 631206 427408 635204 427490
rect 631206 422944 631301 427408
rect 634165 422944 635204 427408
rect 631206 422869 635204 422944
rect 631206 422467 635604 422549
rect 631206 417843 631301 422467
rect 634165 417843 635604 422467
rect 631206 417760 635604 417843
rect -3216 413558 1182 413640
rect -3216 408934 -1777 413558
rect 1087 408934 1182 413558
rect -3216 408851 1182 408934
rect -2216 408448 1182 408530
rect -2216 403984 -1777 408448
rect 1087 403984 1182 408448
rect -2216 403920 1182 403984
rect -3216 403518 1182 403600
rect -3216 398894 -1777 403518
rect 1087 398894 1182 403518
rect -3216 398811 1182 398894
rect 631206 388327 635604 388409
rect 631206 383703 631301 388327
rect 634165 383703 635604 388327
rect 631206 383620 635604 383703
rect 631206 378344 635604 378426
rect 631206 373720 631301 378344
rect 634165 373720 635604 378344
rect 631206 373637 635604 373720
rect -3216 40758 1182 40840
rect -3216 36134 -1777 40758
rect 1087 36134 1182 40758
rect -3216 36051 1182 36134
rect 546304 30917 547584 30925
rect 546304 30885 546312 30917
rect -3216 30718 1182 30800
rect -3216 26094 -1777 30718
rect 1087 26094 1182 30718
rect 543584 30638 546312 30885
rect 546304 30613 546312 30638
rect 547576 30613 547584 30917
rect 546304 30605 547584 30613
rect 529744 30433 532658 30483
rect 529744 30209 529796 30433
rect 530660 30209 532658 30433
rect 529744 30164 532658 30209
rect -3216 26011 1182 26094
rect 134544 7832 139976 7881
rect 134544 7608 134595 7832
rect 135459 7738 139976 7832
rect 135459 7608 139772 7738
rect 134544 7594 139772 7608
rect 139916 7594 139976 7738
rect 134544 7560 139976 7594
rect 135904 7168 138678 7214
rect 135904 6944 135947 7168
rect 136811 7164 138678 7168
rect 136811 7020 138472 7164
rect 138616 7020 138678 7164
rect 136811 6944 138678 7020
rect 135904 6894 138678 6944
rect 198943 -112 203749 -22
rect 175700 -225 179302 -135
rect 175700 -1809 175798 -225
rect 179222 -1809 179302 -225
rect 175700 -6251 179302 -1809
rect 198943 -1696 199023 -112
rect 203647 -1696 203749 -112
rect 198943 -2938 203749 -1696
rect 208994 -112 213800 -22
rect 208994 -1696 209074 -112
rect 213698 -1696 213800 -112
rect 208994 -2938 213800 -1696
rect 215005 -225 217749 -135
rect 215005 -1809 215103 -225
rect 217647 -1809 217749 -225
rect 215005 -7342 217749 -1809
rect 215005 -8126 215108 -7342
rect 217572 -8126 217749 -7342
rect 215005 -8197 217749 -8126
<< via3 >>
rect 533467 952770 538091 954354
rect 543448 952770 548072 954354
rect -1777 880134 1087 884758
rect -1777 875184 1087 879648
rect 631301 875694 634165 880318
rect -1777 870094 1087 874718
rect 631301 870744 634165 875208
rect 631301 865643 634165 870267
rect -1777 795652 1087 800276
rect -1777 785673 1087 790297
rect 631301 786495 634165 791119
rect 631301 776512 634165 781136
rect 631301 471895 634165 476519
rect 631301 461912 634165 466536
rect -1777 451052 1087 455676
rect -1777 441073 1087 445697
rect 631301 427894 634165 432518
rect 631301 422944 634165 427408
rect 631301 417843 634165 422467
rect -1777 408934 1087 413558
rect -1777 403984 1087 408448
rect -1777 398894 1087 403518
rect 631301 383703 634165 388327
rect 631301 373720 634165 378344
rect -1777 36134 1087 40758
rect -1777 26094 1087 30718
rect 546312 30613 547576 30917
rect 529796 30209 530660 30433
rect 134595 7608 135459 7832
rect 139772 7594 139916 7738
rect 135947 6944 136811 7168
rect 138472 7020 138616 7164
rect 175798 -1809 179222 -225
rect 199023 -1696 203647 -112
rect 209074 -1696 213698 -112
rect 215103 -1809 217647 -225
rect 215108 -8126 217572 -7342
<< metal4 >>
rect 533387 954354 538193 954482
rect 533387 952770 533467 954354
rect 538091 952770 538193 954354
rect 533387 935910 538193 952770
rect 533387 934074 533550 935910
rect 537946 934074 538193 935910
rect 533387 933992 538193 934074
rect 543368 954354 548174 954482
rect 543368 952770 543448 954354
rect 548072 952770 548174 954354
rect 543368 935910 548174 952770
rect 543368 934074 543531 935910
rect 547927 934074 548174 935910
rect 543368 933992 548174 934074
rect -1858 884758 1182 884840
rect -1858 880134 -1777 884758
rect 1087 880134 1182 884758
rect 631206 880318 634246 880400
rect -1858 880051 1182 880134
rect -1858 879648 1182 879730
rect -1858 875184 -1777 879648
rect 1087 875184 1182 879648
rect 631206 875694 631301 880318
rect 634165 875694 634246 880318
rect 631206 875611 634246 875694
rect -1858 875120 1182 875184
rect 631206 875208 634246 875290
rect -1858 874718 1182 874800
rect -1858 870094 -1777 874718
rect 1087 870094 1182 874718
rect 631206 870744 631301 875208
rect 634165 870744 634246 875208
rect 631206 870669 634246 870744
rect 631206 870267 634246 870349
rect -1858 870011 1182 870094
rect 631206 865643 631301 870267
rect 634165 865643 634246 870267
rect 631206 865560 634246 865643
rect -1858 800276 1182 800358
rect -1858 795652 -1777 800276
rect 1087 795652 1182 800276
rect -1858 795569 1182 795652
rect 631206 791119 634246 791201
rect -1858 790297 1182 790318
rect -1858 785673 -1777 790297
rect 1087 785673 1182 790297
rect 631206 786495 631301 791119
rect 634165 786495 634246 791119
rect 631206 786412 634246 786495
rect -1858 785589 1182 785673
rect 631206 781136 634246 781218
rect 631206 776512 631301 781136
rect 634165 776512 634246 781136
rect 631206 776429 634246 776512
rect 631206 476519 634246 476601
rect 631206 471895 631301 476519
rect 634165 471895 634246 476519
rect 631206 471812 634246 471895
rect 631206 466536 634246 466618
rect 631206 461912 631301 466536
rect 634165 461912 634246 466536
rect 631206 461829 634246 461912
rect -1858 455676 1182 455758
rect -1858 451052 -1777 455676
rect 1087 451052 1182 455676
rect -1858 450969 1182 451052
rect -1858 445697 1182 445718
rect -1858 441073 -1777 445697
rect 1087 441073 1182 445697
rect -1858 440989 1182 441073
rect 631206 432518 634246 432600
rect 631206 427894 631301 432518
rect 634165 427894 634246 432518
rect 631206 427811 634246 427894
rect 631206 427408 634246 427490
rect 631206 422944 631301 427408
rect 634165 422944 634246 427408
rect 631206 422869 634246 422944
rect 631206 422467 634246 422549
rect 631206 417843 631301 422467
rect 634165 417843 634246 422467
rect 631206 417760 634246 417843
rect -1858 413558 1182 413640
rect -1858 408934 -1777 413558
rect 1087 408934 1182 413558
rect -1858 408851 1182 408934
rect -1858 408448 1182 408530
rect -1858 403984 -1777 408448
rect 1087 403984 1182 408448
rect -1858 403920 1182 403984
rect -1858 403518 1182 403600
rect -1858 398894 -1777 403518
rect 1087 398894 1182 403518
rect -1858 398811 1182 398894
rect 631206 388327 634246 388409
rect 631206 383703 631301 388327
rect 634165 383703 634246 388327
rect 631206 383620 634246 383703
rect 631206 378344 634246 378426
rect 631206 373720 631301 378344
rect 634165 373720 634246 378344
rect 631206 373637 634246 373720
rect -1858 40758 1182 40840
rect -1858 36134 -1777 40758
rect 1087 36134 1182 40758
rect -1858 36051 1182 36134
rect -1858 30718 1182 30800
rect -1858 26094 -1777 30718
rect 1087 26094 1182 30718
rect 543604 30162 546064 30491
rect 531104 29454 532817 29855
rect 135904 26314 136864 26476
rect -1858 26011 1182 26094
rect 135904 25438 135946 26314
rect 136822 25438 136864 26314
rect 134544 24714 135504 24876
rect 134544 23838 134586 24714
rect 135462 23838 135504 24714
rect 134544 7832 135504 23838
rect 134544 7608 134595 7832
rect 135459 7608 135504 7832
rect 134544 7560 135504 7608
rect 135904 7168 136864 25438
rect 215005 26314 217749 26476
rect 215005 25438 215151 26314
rect 217627 25438 217749 26314
rect 175700 24714 179302 24876
rect 175700 23838 175946 24714
rect 179062 23838 179302 24714
rect 135904 6944 135947 7168
rect 136811 6944 136864 7168
rect 135904 6894 136864 6944
rect 137400 5713 137791 5896
rect 137400 5477 137476 5713
rect 137712 5477 137791 5713
rect 137400 5393 137791 5477
rect 137400 5157 137476 5393
rect 137712 5157 137791 5393
rect 137400 5073 137791 5157
rect 137400 4837 137476 5073
rect 137712 4837 137791 5073
rect 137400 4753 137791 4837
rect 137400 4517 137476 4753
rect 137712 4517 137791 4753
rect 137400 4296 137791 4517
rect 138800 3774 139282 5896
rect 138800 3538 138932 3774
rect 139168 3538 139282 3774
rect 138800 3454 139282 3538
rect 138800 3218 138932 3454
rect 139168 3218 139282 3454
rect 138800 3134 139282 3218
rect 138800 2898 138932 3134
rect 139168 2898 139282 3134
rect 138800 2814 139282 2898
rect 138800 2578 138932 2814
rect 139168 2578 139282 2814
rect 138800 2376 139282 2578
rect 175700 -225 179302 23838
rect 175700 -1809 175798 -225
rect 179222 -1809 179302 -225
rect 175700 -1937 179302 -1809
rect 198943 5854 203749 5896
rect 198943 4338 199106 5854
rect 203502 4338 203749 5854
rect 198943 -112 203749 4338
rect 198943 -1696 199023 -112
rect 203647 -1696 203749 -112
rect 198943 -1824 203749 -1696
rect 208994 5854 213800 5896
rect 208994 4338 209157 5854
rect 213553 4338 213800 5854
rect 208994 -112 213800 4338
rect 208994 -1696 209074 -112
rect 213698 -1696 213800 -112
rect 208994 -1824 213800 -1696
rect 215005 -225 217749 25438
rect 215005 -1809 215103 -225
rect 217647 -1809 217749 -225
rect 215005 -1937 217749 -1809
rect 215005 -7342 217749 -7285
rect 215005 -8126 215108 -7342
rect 217572 -8126 217749 -7342
rect 215005 -8197 217749 -8126
<< via4 >>
rect 533550 934074 537946 935910
rect 543531 934074 547927 935910
rect -1736 880322 1060 884718
rect 13046 880322 13922 884718
rect -1736 875212 1060 879608
rect 11846 875212 12722 879608
rect 627098 875882 627974 880278
rect 631328 875882 634124 880278
rect -1736 870282 1060 874678
rect 13046 870282 13922 874678
rect 625898 870772 626774 875168
rect 631328 870772 634124 875168
rect 627098 865831 627974 870227
rect 631328 865831 634124 870227
rect -1736 795840 1060 800236
rect 7046 795840 7922 800236
rect -1736 785861 1060 790257
rect 7046 785861 7922 790257
rect 621098 786683 621974 791079
rect 631328 786683 634124 791079
rect 621098 776700 621974 781096
rect 631328 776700 634124 781096
rect 621098 472083 621974 476479
rect 631328 472083 634124 476479
rect 621098 462100 621974 466496
rect 631328 462100 634124 466496
rect -1736 451240 1060 455636
rect 8246 451240 9122 455636
rect -1736 441261 1060 445657
rect 8246 441261 9122 445657
rect 625898 428082 626774 432478
rect 631328 428082 634124 432478
rect 627098 422972 627974 427368
rect 631328 422972 634124 427368
rect 625898 418031 626774 422427
rect 631328 418031 634124 422427
rect -1736 409122 1060 413518
rect 11846 409122 12722 413518
rect -1736 404012 1060 408408
rect 13046 404012 13922 408408
rect -1736 399082 1060 403478
rect 11846 399082 12722 403478
rect 622298 383891 623174 388287
rect 631328 383891 634124 388287
rect 622298 373908 623174 378304
rect 631328 373908 634124 378304
rect -1736 36322 1060 40718
rect 2246 36322 3122 40718
rect -1736 26282 1060 30678
rect 2246 26282 3122 30678
rect 135946 25438 136822 26314
rect 134586 23838 135462 24714
rect 215151 25438 217627 26314
rect 175946 23838 179062 24714
rect 137476 5477 137712 5713
rect 137476 5157 137712 5393
rect 137476 4837 137712 5073
rect 137476 4517 137712 4753
rect 138932 3538 139168 3774
rect 138932 3218 139168 3454
rect 138932 2898 139168 3134
rect 138932 2578 139168 2814
rect 199106 4338 203502 5854
rect 209157 4338 213553 5854
<< metal5 >>
rect -1858 884718 13984 884840
rect -1858 880322 -1736 884718
rect 1060 880322 13046 884718
rect 13922 880322 13984 884718
rect -1858 880050 13984 880322
rect 627036 880278 634246 880400
rect -1858 879608 12784 879730
rect -1858 875212 -1736 879608
rect 1060 875212 11846 879608
rect 12722 875212 12784 879608
rect 627036 875882 627098 880278
rect 627974 875882 631328 880278
rect 634124 875882 634246 880278
rect 627036 875610 634246 875882
rect -1858 875120 12784 875212
rect 625836 875168 634246 875290
rect -1858 874678 13984 874800
rect -1858 870282 -1736 874678
rect 1060 870282 13046 874678
rect 13922 870282 13984 874678
rect 625836 870772 625898 875168
rect 626774 870772 631328 875168
rect 634124 870772 634246 875168
rect 625836 870669 634246 870772
rect -1858 870010 13984 870282
rect 627036 870227 634246 870349
rect 627036 865831 627098 870227
rect 627974 865831 631328 870227
rect 634124 865831 634246 870227
rect 627036 865559 634246 865831
rect -1858 800236 7984 800358
rect -1858 795840 -1736 800236
rect 1060 795840 7046 800236
rect 7922 795840 7984 800236
rect -1858 795568 7984 795840
rect 621036 791079 634246 791201
rect -1858 790257 7984 790379
rect -1858 785861 -1736 790257
rect 1060 785861 7046 790257
rect 7922 785861 7984 790257
rect 621036 786683 621098 791079
rect 621974 786683 631328 791079
rect 634124 786683 634246 791079
rect 621036 786411 634246 786683
rect -1858 785589 7984 785861
rect 621036 781096 634246 781218
rect 621036 776700 621098 781096
rect 621974 776700 631328 781096
rect 634124 776700 634246 781096
rect 621036 776428 634246 776700
rect 621036 476479 634246 476601
rect 621036 472083 621098 476479
rect 621974 472083 631328 476479
rect 634124 472083 634246 476479
rect 621036 471811 634246 472083
rect 621036 466496 634246 466618
rect 621036 462100 621098 466496
rect 621974 462100 631328 466496
rect 634124 462100 634246 466496
rect 621036 461828 634246 462100
rect -1858 455636 9184 455758
rect -1858 451240 -1736 455636
rect 1060 451240 8246 455636
rect 9122 451240 9184 455636
rect -1858 450968 9184 451240
rect -1858 445657 9184 445779
rect -1858 441261 -1736 445657
rect 1060 441261 8246 445657
rect 9122 441261 9184 445657
rect -1858 440989 9184 441261
rect 625836 432478 634246 432600
rect 625836 428082 625898 432478
rect 626774 428082 631328 432478
rect 634124 428082 634246 432478
rect 625836 427810 634246 428082
rect 627036 427368 634246 427490
rect 627036 422972 627098 427368
rect 627974 422972 631328 427368
rect 634124 422972 634246 427368
rect 627036 422869 634246 422972
rect 625836 422427 634246 422549
rect 625836 418031 625898 422427
rect 626774 418031 631328 422427
rect 634124 418031 634246 422427
rect 625836 417759 634246 418031
rect -1858 413518 12784 413640
rect -1858 409122 -1736 413518
rect 1060 409122 11846 413518
rect 12722 409122 12784 413518
rect -1858 408850 12784 409122
rect -1858 408408 13984 408530
rect -1858 404012 -1736 408408
rect 1060 404012 13046 408408
rect 13922 404012 13984 408408
rect -1858 403920 13984 404012
rect -1858 403478 12784 403600
rect -1858 399082 -1736 403478
rect 1060 399082 11846 403478
rect 12722 399082 12784 403478
rect -1858 398810 12784 399082
rect 622236 388287 634246 388409
rect 622236 383891 622298 388287
rect 623174 383891 631328 388287
rect 634124 383891 634246 388287
rect 622236 383619 634246 383891
rect 622236 378304 634246 378426
rect 622236 373908 622298 378304
rect 623174 373908 631328 378304
rect 634124 373908 634246 378304
rect 622236 373636 634246 373908
rect -1858 40718 3184 40840
rect -1858 36322 -1736 40718
rect 1060 36322 2246 40718
rect 3122 36322 3184 40718
rect -1858 36050 3184 36322
rect -1858 30678 3184 30800
rect -1858 26282 -1736 30678
rect 1060 26282 2246 30678
rect 3122 26282 3184 30678
rect -1858 26010 3184 26282
<< properties >>
string FIXED_BBOX 0 0 200 200
<< end >>
