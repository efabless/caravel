VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_protect
  CLASS BLOCK ;
  FOREIGN mgmt_protect ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 120.000 ;
  PIN caravel_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 19.760 4.000 20.360 ;
    END
  END caravel_clk
  PIN caravel_clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 59.200 4.000 59.800 ;
    END
  END caravel_clk2
  PIN caravel_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 99.320 4.000 99.920 ;
    END
  END caravel_rstn
  PIN la_data_in_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 116.000 237.270 122.000 ;
    END
  END la_data_in_core[0]
  PIN la_data_in_core[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 116.000 905.190 122.000 ;
    END
  END la_data_in_core[100]
  PIN la_data_in_core[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 116.000 911.630 122.000 ;
    END
  END la_data_in_core[101]
  PIN la_data_in_core[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 116.000 918.530 122.000 ;
    END
  END la_data_in_core[102]
  PIN la_data_in_core[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 116.000 924.970 122.000 ;
    END
  END la_data_in_core[103]
  PIN la_data_in_core[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 116.000 931.870 122.000 ;
    END
  END la_data_in_core[104]
  PIN la_data_in_core[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 116.000 938.310 122.000 ;
    END
  END la_data_in_core[105]
  PIN la_data_in_core[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 116.000 945.210 122.000 ;
    END
  END la_data_in_core[106]
  PIN la_data_in_core[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 116.000 951.650 122.000 ;
    END
  END la_data_in_core[107]
  PIN la_data_in_core[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.270 116.000 958.550 122.000 ;
    END
  END la_data_in_core[108]
  PIN la_data_in_core[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 116.000 964.990 122.000 ;
    END
  END la_data_in_core[109]
  PIN la_data_in_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 116.000 303.970 122.000 ;
    END
  END la_data_in_core[10]
  PIN la_data_in_core[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.610 116.000 971.890 122.000 ;
    END
  END la_data_in_core[110]
  PIN la_data_in_core[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.050 116.000 978.330 122.000 ;
    END
  END la_data_in_core[111]
  PIN la_data_in_core[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 116.000 985.230 122.000 ;
    END
  END la_data_in_core[112]
  PIN la_data_in_core[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 116.000 991.670 122.000 ;
    END
  END la_data_in_core[113]
  PIN la_data_in_core[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 116.000 998.570 122.000 ;
    END
  END la_data_in_core[114]
  PIN la_data_in_core[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 116.000 1005.010 122.000 ;
    END
  END la_data_in_core[115]
  PIN la_data_in_core[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.630 116.000 1011.910 122.000 ;
    END
  END la_data_in_core[116]
  PIN la_data_in_core[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.070 116.000 1018.350 122.000 ;
    END
  END la_data_in_core[117]
  PIN la_data_in_core[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.970 116.000 1025.250 122.000 ;
    END
  END la_data_in_core[118]
  PIN la_data_in_core[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.410 116.000 1031.690 122.000 ;
    END
  END la_data_in_core[119]
  PIN la_data_in_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 116.000 310.410 122.000 ;
    END
  END la_data_in_core[11]
  PIN la_data_in_core[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.310 116.000 1038.590 122.000 ;
    END
  END la_data_in_core[120]
  PIN la_data_in_core[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 116.000 1045.030 122.000 ;
    END
  END la_data_in_core[121]
  PIN la_data_in_core[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 116.000 1051.930 122.000 ;
    END
  END la_data_in_core[122]
  PIN la_data_in_core[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 116.000 1058.830 122.000 ;
    END
  END la_data_in_core[123]
  PIN la_data_in_core[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.990 116.000 1065.270 122.000 ;
    END
  END la_data_in_core[124]
  PIN la_data_in_core[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 116.000 1072.170 122.000 ;
    END
  END la_data_in_core[125]
  PIN la_data_in_core[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.330 116.000 1078.610 122.000 ;
    END
  END la_data_in_core[126]
  PIN la_data_in_core[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 116.000 1085.510 122.000 ;
    END
  END la_data_in_core[127]
  PIN la_data_in_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 116.000 317.310 122.000 ;
    END
  END la_data_in_core[12]
  PIN la_data_in_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 116.000 323.750 122.000 ;
    END
  END la_data_in_core[13]
  PIN la_data_in_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 116.000 330.650 122.000 ;
    END
  END la_data_in_core[14]
  PIN la_data_in_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 116.000 337.090 122.000 ;
    END
  END la_data_in_core[15]
  PIN la_data_in_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 116.000 343.990 122.000 ;
    END
  END la_data_in_core[16]
  PIN la_data_in_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 116.000 350.430 122.000 ;
    END
  END la_data_in_core[17]
  PIN la_data_in_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 116.000 357.330 122.000 ;
    END
  END la_data_in_core[18]
  PIN la_data_in_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 116.000 363.770 122.000 ;
    END
  END la_data_in_core[19]
  PIN la_data_in_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 116.000 243.710 122.000 ;
    END
  END la_data_in_core[1]
  PIN la_data_in_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 116.000 370.670 122.000 ;
    END
  END la_data_in_core[20]
  PIN la_data_in_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 116.000 377.110 122.000 ;
    END
  END la_data_in_core[21]
  PIN la_data_in_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 116.000 384.010 122.000 ;
    END
  END la_data_in_core[22]
  PIN la_data_in_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 116.000 390.910 122.000 ;
    END
  END la_data_in_core[23]
  PIN la_data_in_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 116.000 397.350 122.000 ;
    END
  END la_data_in_core[24]
  PIN la_data_in_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 116.000 404.250 122.000 ;
    END
  END la_data_in_core[25]
  PIN la_data_in_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 116.000 410.690 122.000 ;
    END
  END la_data_in_core[26]
  PIN la_data_in_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 116.000 417.590 122.000 ;
    END
  END la_data_in_core[27]
  PIN la_data_in_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 116.000 424.030 122.000 ;
    END
  END la_data_in_core[28]
  PIN la_data_in_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 116.000 430.930 122.000 ;
    END
  END la_data_in_core[29]
  PIN la_data_in_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 116.000 250.610 122.000 ;
    END
  END la_data_in_core[2]
  PIN la_data_in_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 116.000 437.370 122.000 ;
    END
  END la_data_in_core[30]
  PIN la_data_in_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 116.000 444.270 122.000 ;
    END
  END la_data_in_core[31]
  PIN la_data_in_core[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 116.000 450.710 122.000 ;
    END
  END la_data_in_core[32]
  PIN la_data_in_core[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 116.000 457.610 122.000 ;
    END
  END la_data_in_core[33]
  PIN la_data_in_core[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 116.000 464.050 122.000 ;
    END
  END la_data_in_core[34]
  PIN la_data_in_core[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 116.000 470.950 122.000 ;
    END
  END la_data_in_core[35]
  PIN la_data_in_core[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 116.000 477.390 122.000 ;
    END
  END la_data_in_core[36]
  PIN la_data_in_core[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 116.000 484.290 122.000 ;
    END
  END la_data_in_core[37]
  PIN la_data_in_core[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 116.000 490.730 122.000 ;
    END
  END la_data_in_core[38]
  PIN la_data_in_core[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 116.000 497.630 122.000 ;
    END
  END la_data_in_core[39]
  PIN la_data_in_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 116.000 257.050 122.000 ;
    END
  END la_data_in_core[3]
  PIN la_data_in_core[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 116.000 504.070 122.000 ;
    END
  END la_data_in_core[40]
  PIN la_data_in_core[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 116.000 510.970 122.000 ;
    END
  END la_data_in_core[41]
  PIN la_data_in_core[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 116.000 517.410 122.000 ;
    END
  END la_data_in_core[42]
  PIN la_data_in_core[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 116.000 524.310 122.000 ;
    END
  END la_data_in_core[43]
  PIN la_data_in_core[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 116.000 530.750 122.000 ;
    END
  END la_data_in_core[44]
  PIN la_data_in_core[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 116.000 537.650 122.000 ;
    END
  END la_data_in_core[45]
  PIN la_data_in_core[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 116.000 544.090 122.000 ;
    END
  END la_data_in_core[46]
  PIN la_data_in_core[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 116.000 550.990 122.000 ;
    END
  END la_data_in_core[47]
  PIN la_data_in_core[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 116.000 557.890 122.000 ;
    END
  END la_data_in_core[48]
  PIN la_data_in_core[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 116.000 564.330 122.000 ;
    END
  END la_data_in_core[49]
  PIN la_data_in_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 116.000 263.950 122.000 ;
    END
  END la_data_in_core[4]
  PIN la_data_in_core[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 116.000 571.230 122.000 ;
    END
  END la_data_in_core[50]
  PIN la_data_in_core[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 116.000 577.670 122.000 ;
    END
  END la_data_in_core[51]
  PIN la_data_in_core[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 116.000 584.570 122.000 ;
    END
  END la_data_in_core[52]
  PIN la_data_in_core[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 116.000 591.010 122.000 ;
    END
  END la_data_in_core[53]
  PIN la_data_in_core[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 116.000 597.910 122.000 ;
    END
  END la_data_in_core[54]
  PIN la_data_in_core[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 116.000 604.350 122.000 ;
    END
  END la_data_in_core[55]
  PIN la_data_in_core[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 116.000 611.250 122.000 ;
    END
  END la_data_in_core[56]
  PIN la_data_in_core[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 116.000 617.690 122.000 ;
    END
  END la_data_in_core[57]
  PIN la_data_in_core[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 116.000 624.590 122.000 ;
    END
  END la_data_in_core[58]
  PIN la_data_in_core[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 116.000 631.030 122.000 ;
    END
  END la_data_in_core[59]
  PIN la_data_in_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 116.000 270.390 122.000 ;
    END
  END la_data_in_core[5]
  PIN la_data_in_core[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 116.000 637.930 122.000 ;
    END
  END la_data_in_core[60]
  PIN la_data_in_core[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 116.000 644.370 122.000 ;
    END
  END la_data_in_core[61]
  PIN la_data_in_core[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 116.000 651.270 122.000 ;
    END
  END la_data_in_core[62]
  PIN la_data_in_core[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 116.000 657.710 122.000 ;
    END
  END la_data_in_core[63]
  PIN la_data_in_core[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 116.000 664.610 122.000 ;
    END
  END la_data_in_core[64]
  PIN la_data_in_core[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 116.000 671.050 122.000 ;
    END
  END la_data_in_core[65]
  PIN la_data_in_core[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 116.000 677.950 122.000 ;
    END
  END la_data_in_core[66]
  PIN la_data_in_core[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 116.000 684.390 122.000 ;
    END
  END la_data_in_core[67]
  PIN la_data_in_core[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 116.000 691.290 122.000 ;
    END
  END la_data_in_core[68]
  PIN la_data_in_core[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 116.000 697.730 122.000 ;
    END
  END la_data_in_core[69]
  PIN la_data_in_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 116.000 277.290 122.000 ;
    END
  END la_data_in_core[6]
  PIN la_data_in_core[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 116.000 704.630 122.000 ;
    END
  END la_data_in_core[70]
  PIN la_data_in_core[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 116.000 711.070 122.000 ;
    END
  END la_data_in_core[71]
  PIN la_data_in_core[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 116.000 717.970 122.000 ;
    END
  END la_data_in_core[72]
  PIN la_data_in_core[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 116.000 724.870 122.000 ;
    END
  END la_data_in_core[73]
  PIN la_data_in_core[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 116.000 731.310 122.000 ;
    END
  END la_data_in_core[74]
  PIN la_data_in_core[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 116.000 738.210 122.000 ;
    END
  END la_data_in_core[75]
  PIN la_data_in_core[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 116.000 744.650 122.000 ;
    END
  END la_data_in_core[76]
  PIN la_data_in_core[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 116.000 751.550 122.000 ;
    END
  END la_data_in_core[77]
  PIN la_data_in_core[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 116.000 757.990 122.000 ;
    END
  END la_data_in_core[78]
  PIN la_data_in_core[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 116.000 764.890 122.000 ;
    END
  END la_data_in_core[79]
  PIN la_data_in_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 116.000 283.730 122.000 ;
    END
  END la_data_in_core[7]
  PIN la_data_in_core[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 116.000 771.330 122.000 ;
    END
  END la_data_in_core[80]
  PIN la_data_in_core[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 116.000 778.230 122.000 ;
    END
  END la_data_in_core[81]
  PIN la_data_in_core[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 116.000 784.670 122.000 ;
    END
  END la_data_in_core[82]
  PIN la_data_in_core[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 116.000 791.570 122.000 ;
    END
  END la_data_in_core[83]
  PIN la_data_in_core[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 116.000 798.010 122.000 ;
    END
  END la_data_in_core[84]
  PIN la_data_in_core[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 116.000 804.910 122.000 ;
    END
  END la_data_in_core[85]
  PIN la_data_in_core[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 116.000 811.350 122.000 ;
    END
  END la_data_in_core[86]
  PIN la_data_in_core[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 116.000 818.250 122.000 ;
    END
  END la_data_in_core[87]
  PIN la_data_in_core[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 116.000 824.690 122.000 ;
    END
  END la_data_in_core[88]
  PIN la_data_in_core[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 116.000 831.590 122.000 ;
    END
  END la_data_in_core[89]
  PIN la_data_in_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 116.000 290.630 122.000 ;
    END
  END la_data_in_core[8]
  PIN la_data_in_core[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 116.000 838.030 122.000 ;
    END
  END la_data_in_core[90]
  PIN la_data_in_core[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 116.000 844.930 122.000 ;
    END
  END la_data_in_core[91]
  PIN la_data_in_core[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 116.000 851.370 122.000 ;
    END
  END la_data_in_core[92]
  PIN la_data_in_core[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 116.000 858.270 122.000 ;
    END
  END la_data_in_core[93]
  PIN la_data_in_core[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430 116.000 864.710 122.000 ;
    END
  END la_data_in_core[94]
  PIN la_data_in_core[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.330 116.000 871.610 122.000 ;
    END
  END la_data_in_core[95]
  PIN la_data_in_core[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 116.000 878.050 122.000 ;
    END
  END la_data_in_core[96]
  PIN la_data_in_core[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 116.000 884.950 122.000 ;
    END
  END la_data_in_core[97]
  PIN la_data_in_core[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 116.000 891.850 122.000 ;
    END
  END la_data_in_core[98]
  PIN la_data_in_core[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.010 116.000 898.290 122.000 ;
    END
  END la_data_in_core[99]
  PIN la_data_in_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 116.000 297.070 122.000 ;
    END
  END la_data_in_core[9]
  PIN la_data_in_mprj[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 -2.000 0.830 4.000 ;
    END
  END la_data_in_mprj[0]
  PIN la_data_in_mprj[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 -2.000 713.830 4.000 ;
    END
  END la_data_in_mprj[100]
  PIN la_data_in_mprj[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 -2.000 720.730 4.000 ;
    END
  END la_data_in_mprj[101]
  PIN la_data_in_mprj[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 -2.000 728.090 4.000 ;
    END
  END la_data_in_mprj[102]
  PIN la_data_in_mprj[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 -2.000 734.990 4.000 ;
    END
  END la_data_in_mprj[103]
  PIN la_data_in_mprj[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 -2.000 742.350 4.000 ;
    END
  END la_data_in_mprj[104]
  PIN la_data_in_mprj[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 -2.000 749.250 4.000 ;
    END
  END la_data_in_mprj[105]
  PIN la_data_in_mprj[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 -2.000 756.610 4.000 ;
    END
  END la_data_in_mprj[106]
  PIN la_data_in_mprj[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 -2.000 763.510 4.000 ;
    END
  END la_data_in_mprj[107]
  PIN la_data_in_mprj[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 -2.000 770.870 4.000 ;
    END
  END la_data_in_mprj[108]
  PIN la_data_in_mprj[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 -2.000 777.770 4.000 ;
    END
  END la_data_in_mprj[109]
  PIN la_data_in_mprj[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 -2.000 72.130 4.000 ;
    END
  END la_data_in_mprj[10]
  PIN la_data_in_mprj[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 -2.000 785.130 4.000 ;
    END
  END la_data_in_mprj[110]
  PIN la_data_in_mprj[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.750 -2.000 792.030 4.000 ;
    END
  END la_data_in_mprj[111]
  PIN la_data_in_mprj[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 -2.000 799.390 4.000 ;
    END
  END la_data_in_mprj[112]
  PIN la_data_in_mprj[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 -2.000 806.290 4.000 ;
    END
  END la_data_in_mprj[113]
  PIN la_data_in_mprj[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 -2.000 813.650 4.000 ;
    END
  END la_data_in_mprj[114]
  PIN la_data_in_mprj[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 -2.000 820.550 4.000 ;
    END
  END la_data_in_mprj[115]
  PIN la_data_in_mprj[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 -2.000 827.910 4.000 ;
    END
  END la_data_in_mprj[116]
  PIN la_data_in_mprj[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 -2.000 834.810 4.000 ;
    END
  END la_data_in_mprj[117]
  PIN la_data_in_mprj[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 -2.000 842.170 4.000 ;
    END
  END la_data_in_mprj[118]
  PIN la_data_in_mprj[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 -2.000 849.070 4.000 ;
    END
  END la_data_in_mprj[119]
  PIN la_data_in_mprj[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 -2.000 79.030 4.000 ;
    END
  END la_data_in_mprj[11]
  PIN la_data_in_mprj[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 -2.000 856.430 4.000 ;
    END
  END la_data_in_mprj[120]
  PIN la_data_in_mprj[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 -2.000 863.330 4.000 ;
    END
  END la_data_in_mprj[121]
  PIN la_data_in_mprj[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 -2.000 870.690 4.000 ;
    END
  END la_data_in_mprj[122]
  PIN la_data_in_mprj[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 -2.000 877.590 4.000 ;
    END
  END la_data_in_mprj[123]
  PIN la_data_in_mprj[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 -2.000 884.950 4.000 ;
    END
  END la_data_in_mprj[124]
  PIN la_data_in_mprj[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 -2.000 891.850 4.000 ;
    END
  END la_data_in_mprj[125]
  PIN la_data_in_mprj[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.930 -2.000 899.210 4.000 ;
    END
  END la_data_in_mprj[126]
  PIN la_data_in_mprj[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.830 -2.000 906.110 4.000 ;
    END
  END la_data_in_mprj[127]
  PIN la_data_in_mprj[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 -2.000 86.390 4.000 ;
    END
  END la_data_in_mprj[12]
  PIN la_data_in_mprj[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 -2.000 93.290 4.000 ;
    END
  END la_data_in_mprj[13]
  PIN la_data_in_mprj[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 -2.000 100.650 4.000 ;
    END
  END la_data_in_mprj[14]
  PIN la_data_in_mprj[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 -2.000 107.550 4.000 ;
    END
  END la_data_in_mprj[15]
  PIN la_data_in_mprj[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 -2.000 114.910 4.000 ;
    END
  END la_data_in_mprj[16]
  PIN la_data_in_mprj[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 -2.000 121.810 4.000 ;
    END
  END la_data_in_mprj[17]
  PIN la_data_in_mprj[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 -2.000 129.170 4.000 ;
    END
  END la_data_in_mprj[18]
  PIN la_data_in_mprj[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 -2.000 136.070 4.000 ;
    END
  END la_data_in_mprj[19]
  PIN la_data_in_mprj[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 -2.000 7.730 4.000 ;
    END
  END la_data_in_mprj[1]
  PIN la_data_in_mprj[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 -2.000 143.430 4.000 ;
    END
  END la_data_in_mprj[20]
  PIN la_data_in_mprj[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 -2.000 150.330 4.000 ;
    END
  END la_data_in_mprj[21]
  PIN la_data_in_mprj[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 -2.000 157.690 4.000 ;
    END
  END la_data_in_mprj[22]
  PIN la_data_in_mprj[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 -2.000 164.590 4.000 ;
    END
  END la_data_in_mprj[23]
  PIN la_data_in_mprj[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 -2.000 171.950 4.000 ;
    END
  END la_data_in_mprj[24]
  PIN la_data_in_mprj[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 -2.000 178.850 4.000 ;
    END
  END la_data_in_mprj[25]
  PIN la_data_in_mprj[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 -2.000 186.210 4.000 ;
    END
  END la_data_in_mprj[26]
  PIN la_data_in_mprj[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 -2.000 193.110 4.000 ;
    END
  END la_data_in_mprj[27]
  PIN la_data_in_mprj[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 -2.000 200.470 4.000 ;
    END
  END la_data_in_mprj[28]
  PIN la_data_in_mprj[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 -2.000 207.370 4.000 ;
    END
  END la_data_in_mprj[29]
  PIN la_data_in_mprj[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 -2.000 15.090 4.000 ;
    END
  END la_data_in_mprj[2]
  PIN la_data_in_mprj[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 -2.000 214.730 4.000 ;
    END
  END la_data_in_mprj[30]
  PIN la_data_in_mprj[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 -2.000 221.630 4.000 ;
    END
  END la_data_in_mprj[31]
  PIN la_data_in_mprj[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 -2.000 228.990 4.000 ;
    END
  END la_data_in_mprj[32]
  PIN la_data_in_mprj[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 -2.000 235.890 4.000 ;
    END
  END la_data_in_mprj[33]
  PIN la_data_in_mprj[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 -2.000 243.250 4.000 ;
    END
  END la_data_in_mprj[34]
  PIN la_data_in_mprj[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 -2.000 250.150 4.000 ;
    END
  END la_data_in_mprj[35]
  PIN la_data_in_mprj[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 -2.000 257.510 4.000 ;
    END
  END la_data_in_mprj[36]
  PIN la_data_in_mprj[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 -2.000 264.410 4.000 ;
    END
  END la_data_in_mprj[37]
  PIN la_data_in_mprj[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 -2.000 271.770 4.000 ;
    END
  END la_data_in_mprj[38]
  PIN la_data_in_mprj[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 -2.000 278.670 4.000 ;
    END
  END la_data_in_mprj[39]
  PIN la_data_in_mprj[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 -2.000 21.990 4.000 ;
    END
  END la_data_in_mprj[3]
  PIN la_data_in_mprj[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 -2.000 286.030 4.000 ;
    END
  END la_data_in_mprj[40]
  PIN la_data_in_mprj[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 -2.000 292.930 4.000 ;
    END
  END la_data_in_mprj[41]
  PIN la_data_in_mprj[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 -2.000 300.290 4.000 ;
    END
  END la_data_in_mprj[42]
  PIN la_data_in_mprj[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 -2.000 307.190 4.000 ;
    END
  END la_data_in_mprj[43]
  PIN la_data_in_mprj[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 -2.000 314.550 4.000 ;
    END
  END la_data_in_mprj[44]
  PIN la_data_in_mprj[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 -2.000 321.450 4.000 ;
    END
  END la_data_in_mprj[45]
  PIN la_data_in_mprj[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 -2.000 328.810 4.000 ;
    END
  END la_data_in_mprj[46]
  PIN la_data_in_mprj[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 -2.000 335.710 4.000 ;
    END
  END la_data_in_mprj[47]
  PIN la_data_in_mprj[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 -2.000 343.070 4.000 ;
    END
  END la_data_in_mprj[48]
  PIN la_data_in_mprj[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 -2.000 349.970 4.000 ;
    END
  END la_data_in_mprj[49]
  PIN la_data_in_mprj[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 -2.000 29.350 4.000 ;
    END
  END la_data_in_mprj[4]
  PIN la_data_in_mprj[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 -2.000 357.330 4.000 ;
    END
  END la_data_in_mprj[50]
  PIN la_data_in_mprj[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 -2.000 364.230 4.000 ;
    END
  END la_data_in_mprj[51]
  PIN la_data_in_mprj[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 -2.000 371.590 4.000 ;
    END
  END la_data_in_mprj[52]
  PIN la_data_in_mprj[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 -2.000 378.490 4.000 ;
    END
  END la_data_in_mprj[53]
  PIN la_data_in_mprj[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 -2.000 385.850 4.000 ;
    END
  END la_data_in_mprj[54]
  PIN la_data_in_mprj[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 -2.000 392.750 4.000 ;
    END
  END la_data_in_mprj[55]
  PIN la_data_in_mprj[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 -2.000 400.110 4.000 ;
    END
  END la_data_in_mprj[56]
  PIN la_data_in_mprj[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 -2.000 407.010 4.000 ;
    END
  END la_data_in_mprj[57]
  PIN la_data_in_mprj[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 -2.000 414.370 4.000 ;
    END
  END la_data_in_mprj[58]
  PIN la_data_in_mprj[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 -2.000 421.270 4.000 ;
    END
  END la_data_in_mprj[59]
  PIN la_data_in_mprj[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 -2.000 36.250 4.000 ;
    END
  END la_data_in_mprj[5]
  PIN la_data_in_mprj[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 -2.000 428.630 4.000 ;
    END
  END la_data_in_mprj[60]
  PIN la_data_in_mprj[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 -2.000 435.530 4.000 ;
    END
  END la_data_in_mprj[61]
  PIN la_data_in_mprj[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 -2.000 442.890 4.000 ;
    END
  END la_data_in_mprj[62]
  PIN la_data_in_mprj[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 -2.000 449.790 4.000 ;
    END
  END la_data_in_mprj[63]
  PIN la_data_in_mprj[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 -2.000 457.150 4.000 ;
    END
  END la_data_in_mprj[64]
  PIN la_data_in_mprj[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 -2.000 464.050 4.000 ;
    END
  END la_data_in_mprj[65]
  PIN la_data_in_mprj[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 -2.000 471.410 4.000 ;
    END
  END la_data_in_mprj[66]
  PIN la_data_in_mprj[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 -2.000 478.310 4.000 ;
    END
  END la_data_in_mprj[67]
  PIN la_data_in_mprj[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 -2.000 485.670 4.000 ;
    END
  END la_data_in_mprj[68]
  PIN la_data_in_mprj[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 -2.000 492.570 4.000 ;
    END
  END la_data_in_mprj[69]
  PIN la_data_in_mprj[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 -2.000 43.610 4.000 ;
    END
  END la_data_in_mprj[6]
  PIN la_data_in_mprj[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 -2.000 499.930 4.000 ;
    END
  END la_data_in_mprj[70]
  PIN la_data_in_mprj[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 -2.000 506.830 4.000 ;
    END
  END la_data_in_mprj[71]
  PIN la_data_in_mprj[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 -2.000 514.190 4.000 ;
    END
  END la_data_in_mprj[72]
  PIN la_data_in_mprj[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 -2.000 521.090 4.000 ;
    END
  END la_data_in_mprj[73]
  PIN la_data_in_mprj[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 -2.000 528.450 4.000 ;
    END
  END la_data_in_mprj[74]
  PIN la_data_in_mprj[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 -2.000 535.350 4.000 ;
    END
  END la_data_in_mprj[75]
  PIN la_data_in_mprj[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 -2.000 542.710 4.000 ;
    END
  END la_data_in_mprj[76]
  PIN la_data_in_mprj[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 -2.000 549.610 4.000 ;
    END
  END la_data_in_mprj[77]
  PIN la_data_in_mprj[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 -2.000 556.970 4.000 ;
    END
  END la_data_in_mprj[78]
  PIN la_data_in_mprj[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 -2.000 563.870 4.000 ;
    END
  END la_data_in_mprj[79]
  PIN la_data_in_mprj[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 -2.000 50.510 4.000 ;
    END
  END la_data_in_mprj[7]
  PIN la_data_in_mprj[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 -2.000 571.230 4.000 ;
    END
  END la_data_in_mprj[80]
  PIN la_data_in_mprj[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 -2.000 578.130 4.000 ;
    END
  END la_data_in_mprj[81]
  PIN la_data_in_mprj[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 -2.000 585.490 4.000 ;
    END
  END la_data_in_mprj[82]
  PIN la_data_in_mprj[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 -2.000 592.390 4.000 ;
    END
  END la_data_in_mprj[83]
  PIN la_data_in_mprj[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 -2.000 599.750 4.000 ;
    END
  END la_data_in_mprj[84]
  PIN la_data_in_mprj[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 -2.000 606.650 4.000 ;
    END
  END la_data_in_mprj[85]
  PIN la_data_in_mprj[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.730 -2.000 614.010 4.000 ;
    END
  END la_data_in_mprj[86]
  PIN la_data_in_mprj[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 -2.000 620.910 4.000 ;
    END
  END la_data_in_mprj[87]
  PIN la_data_in_mprj[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 -2.000 628.270 4.000 ;
    END
  END la_data_in_mprj[88]
  PIN la_data_in_mprj[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 -2.000 635.170 4.000 ;
    END
  END la_data_in_mprj[89]
  PIN la_data_in_mprj[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 -2.000 57.870 4.000 ;
    END
  END la_data_in_mprj[8]
  PIN la_data_in_mprj[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 -2.000 642.530 4.000 ;
    END
  END la_data_in_mprj[90]
  PIN la_data_in_mprj[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 -2.000 649.430 4.000 ;
    END
  END la_data_in_mprj[91]
  PIN la_data_in_mprj[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 -2.000 656.790 4.000 ;
    END
  END la_data_in_mprj[92]
  PIN la_data_in_mprj[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 -2.000 663.690 4.000 ;
    END
  END la_data_in_mprj[93]
  PIN la_data_in_mprj[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 -2.000 671.050 4.000 ;
    END
  END la_data_in_mprj[94]
  PIN la_data_in_mprj[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 -2.000 677.950 4.000 ;
    END
  END la_data_in_mprj[95]
  PIN la_data_in_mprj[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 -2.000 685.310 4.000 ;
    END
  END la_data_in_mprj[96]
  PIN la_data_in_mprj[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.930 -2.000 692.210 4.000 ;
    END
  END la_data_in_mprj[97]
  PIN la_data_in_mprj[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 -2.000 699.570 4.000 ;
    END
  END la_data_in_mprj[98]
  PIN la_data_in_mprj[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 -2.000 706.470 4.000 ;
    END
  END la_data_in_mprj[99]
  PIN la_data_in_mprj[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 -2.000 64.770 4.000 ;
    END
  END la_data_in_mprj[9]
  PIN la_data_out_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 116.000 239.110 122.000 ;
    END
  END la_data_out_core[0]
  PIN la_data_out_core[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 116.000 907.030 122.000 ;
    END
  END la_data_out_core[100]
  PIN la_data_out_core[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 116.000 913.930 122.000 ;
    END
  END la_data_out_core[101]
  PIN la_data_out_core[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 116.000 920.370 122.000 ;
    END
  END la_data_out_core[102]
  PIN la_data_out_core[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 116.000 927.270 122.000 ;
    END
  END la_data_out_core[103]
  PIN la_data_out_core[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 116.000 933.710 122.000 ;
    END
  END la_data_out_core[104]
  PIN la_data_out_core[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 116.000 940.610 122.000 ;
    END
  END la_data_out_core[105]
  PIN la_data_out_core[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 116.000 947.510 122.000 ;
    END
  END la_data_out_core[106]
  PIN la_data_out_core[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 116.000 953.950 122.000 ;
    END
  END la_data_out_core[107]
  PIN la_data_out_core[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.570 116.000 960.850 122.000 ;
    END
  END la_data_out_core[108]
  PIN la_data_out_core[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.010 116.000 967.290 122.000 ;
    END
  END la_data_out_core[109]
  PIN la_data_out_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 116.000 306.270 122.000 ;
    END
  END la_data_out_core[10]
  PIN la_data_out_core[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.910 116.000 974.190 122.000 ;
    END
  END la_data_out_core[110]
  PIN la_data_out_core[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 116.000 980.630 122.000 ;
    END
  END la_data_out_core[111]
  PIN la_data_out_core[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 116.000 987.530 122.000 ;
    END
  END la_data_out_core[112]
  PIN la_data_out_core[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 116.000 993.970 122.000 ;
    END
  END la_data_out_core[113]
  PIN la_data_out_core[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 116.000 1000.870 122.000 ;
    END
  END la_data_out_core[114]
  PIN la_data_out_core[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.030 116.000 1007.310 122.000 ;
    END
  END la_data_out_core[115]
  PIN la_data_out_core[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.930 116.000 1014.210 122.000 ;
    END
  END la_data_out_core[116]
  PIN la_data_out_core[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.370 116.000 1020.650 122.000 ;
    END
  END la_data_out_core[117]
  PIN la_data_out_core[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 116.000 1027.550 122.000 ;
    END
  END la_data_out_core[118]
  PIN la_data_out_core[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 116.000 1033.990 122.000 ;
    END
  END la_data_out_core[119]
  PIN la_data_out_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 116.000 312.710 122.000 ;
    END
  END la_data_out_core[11]
  PIN la_data_out_core[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.610 116.000 1040.890 122.000 ;
    END
  END la_data_out_core[120]
  PIN la_data_out_core[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.050 116.000 1047.330 122.000 ;
    END
  END la_data_out_core[121]
  PIN la_data_out_core[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.950 116.000 1054.230 122.000 ;
    END
  END la_data_out_core[122]
  PIN la_data_out_core[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.390 116.000 1060.670 122.000 ;
    END
  END la_data_out_core[123]
  PIN la_data_out_core[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.290 116.000 1067.570 122.000 ;
    END
  END la_data_out_core[124]
  PIN la_data_out_core[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.730 116.000 1074.010 122.000 ;
    END
  END la_data_out_core[125]
  PIN la_data_out_core[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630 116.000 1080.910 122.000 ;
    END
  END la_data_out_core[126]
  PIN la_data_out_core[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.070 116.000 1087.350 122.000 ;
    END
  END la_data_out_core[127]
  PIN la_data_out_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 116.000 319.610 122.000 ;
    END
  END la_data_out_core[12]
  PIN la_data_out_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 116.000 326.050 122.000 ;
    END
  END la_data_out_core[13]
  PIN la_data_out_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 116.000 332.950 122.000 ;
    END
  END la_data_out_core[14]
  PIN la_data_out_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 116.000 339.390 122.000 ;
    END
  END la_data_out_core[15]
  PIN la_data_out_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 116.000 346.290 122.000 ;
    END
  END la_data_out_core[16]
  PIN la_data_out_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 116.000 352.730 122.000 ;
    END
  END la_data_out_core[17]
  PIN la_data_out_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 116.000 359.630 122.000 ;
    END
  END la_data_out_core[18]
  PIN la_data_out_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 116.000 366.070 122.000 ;
    END
  END la_data_out_core[19]
  PIN la_data_out_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 116.000 246.010 122.000 ;
    END
  END la_data_out_core[1]
  PIN la_data_out_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 116.000 372.970 122.000 ;
    END
  END la_data_out_core[20]
  PIN la_data_out_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 116.000 379.410 122.000 ;
    END
  END la_data_out_core[21]
  PIN la_data_out_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 116.000 386.310 122.000 ;
    END
  END la_data_out_core[22]
  PIN la_data_out_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 116.000 392.750 122.000 ;
    END
  END la_data_out_core[23]
  PIN la_data_out_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 116.000 399.650 122.000 ;
    END
  END la_data_out_core[24]
  PIN la_data_out_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 116.000 406.090 122.000 ;
    END
  END la_data_out_core[25]
  PIN la_data_out_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 116.000 412.990 122.000 ;
    END
  END la_data_out_core[26]
  PIN la_data_out_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 116.000 419.430 122.000 ;
    END
  END la_data_out_core[27]
  PIN la_data_out_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 116.000 426.330 122.000 ;
    END
  END la_data_out_core[28]
  PIN la_data_out_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 116.000 432.770 122.000 ;
    END
  END la_data_out_core[29]
  PIN la_data_out_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 116.000 252.450 122.000 ;
    END
  END la_data_out_core[2]
  PIN la_data_out_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 116.000 439.670 122.000 ;
    END
  END la_data_out_core[30]
  PIN la_data_out_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 116.000 446.570 122.000 ;
    END
  END la_data_out_core[31]
  PIN la_data_out_core[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 116.000 453.010 122.000 ;
    END
  END la_data_out_core[32]
  PIN la_data_out_core[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 116.000 459.910 122.000 ;
    END
  END la_data_out_core[33]
  PIN la_data_out_core[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 116.000 466.350 122.000 ;
    END
  END la_data_out_core[34]
  PIN la_data_out_core[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 116.000 473.250 122.000 ;
    END
  END la_data_out_core[35]
  PIN la_data_out_core[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 116.000 479.690 122.000 ;
    END
  END la_data_out_core[36]
  PIN la_data_out_core[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 116.000 486.590 122.000 ;
    END
  END la_data_out_core[37]
  PIN la_data_out_core[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 116.000 493.030 122.000 ;
    END
  END la_data_out_core[38]
  PIN la_data_out_core[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 116.000 499.930 122.000 ;
    END
  END la_data_out_core[39]
  PIN la_data_out_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 116.000 259.350 122.000 ;
    END
  END la_data_out_core[3]
  PIN la_data_out_core[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 116.000 506.370 122.000 ;
    END
  END la_data_out_core[40]
  PIN la_data_out_core[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 116.000 513.270 122.000 ;
    END
  END la_data_out_core[41]
  PIN la_data_out_core[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 116.000 519.710 122.000 ;
    END
  END la_data_out_core[42]
  PIN la_data_out_core[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 116.000 526.610 122.000 ;
    END
  END la_data_out_core[43]
  PIN la_data_out_core[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 116.000 533.050 122.000 ;
    END
  END la_data_out_core[44]
  PIN la_data_out_core[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 116.000 539.950 122.000 ;
    END
  END la_data_out_core[45]
  PIN la_data_out_core[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 116.000 546.390 122.000 ;
    END
  END la_data_out_core[46]
  PIN la_data_out_core[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 116.000 553.290 122.000 ;
    END
  END la_data_out_core[47]
  PIN la_data_out_core[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 116.000 559.730 122.000 ;
    END
  END la_data_out_core[48]
  PIN la_data_out_core[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 116.000 566.630 122.000 ;
    END
  END la_data_out_core[49]
  PIN la_data_out_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 116.000 265.790 122.000 ;
    END
  END la_data_out_core[4]
  PIN la_data_out_core[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 116.000 573.070 122.000 ;
    END
  END la_data_out_core[50]
  PIN la_data_out_core[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 116.000 579.970 122.000 ;
    END
  END la_data_out_core[51]
  PIN la_data_out_core[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 116.000 586.410 122.000 ;
    END
  END la_data_out_core[52]
  PIN la_data_out_core[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 116.000 593.310 122.000 ;
    END
  END la_data_out_core[53]
  PIN la_data_out_core[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 116.000 599.750 122.000 ;
    END
  END la_data_out_core[54]
  PIN la_data_out_core[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 116.000 606.650 122.000 ;
    END
  END la_data_out_core[55]
  PIN la_data_out_core[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 116.000 613.550 122.000 ;
    END
  END la_data_out_core[56]
  PIN la_data_out_core[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 116.000 619.990 122.000 ;
    END
  END la_data_out_core[57]
  PIN la_data_out_core[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 116.000 626.890 122.000 ;
    END
  END la_data_out_core[58]
  PIN la_data_out_core[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 116.000 633.330 122.000 ;
    END
  END la_data_out_core[59]
  PIN la_data_out_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 116.000 272.690 122.000 ;
    END
  END la_data_out_core[5]
  PIN la_data_out_core[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 116.000 640.230 122.000 ;
    END
  END la_data_out_core[60]
  PIN la_data_out_core[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 116.000 646.670 122.000 ;
    END
  END la_data_out_core[61]
  PIN la_data_out_core[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 116.000 653.570 122.000 ;
    END
  END la_data_out_core[62]
  PIN la_data_out_core[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 116.000 660.010 122.000 ;
    END
  END la_data_out_core[63]
  PIN la_data_out_core[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 116.000 666.910 122.000 ;
    END
  END la_data_out_core[64]
  PIN la_data_out_core[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 116.000 673.350 122.000 ;
    END
  END la_data_out_core[65]
  PIN la_data_out_core[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 116.000 680.250 122.000 ;
    END
  END la_data_out_core[66]
  PIN la_data_out_core[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 116.000 686.690 122.000 ;
    END
  END la_data_out_core[67]
  PIN la_data_out_core[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 116.000 693.590 122.000 ;
    END
  END la_data_out_core[68]
  PIN la_data_out_core[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 116.000 700.030 122.000 ;
    END
  END la_data_out_core[69]
  PIN la_data_out_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 116.000 279.590 122.000 ;
    END
  END la_data_out_core[6]
  PIN la_data_out_core[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 116.000 706.930 122.000 ;
    END
  END la_data_out_core[70]
  PIN la_data_out_core[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 116.000 713.370 122.000 ;
    END
  END la_data_out_core[71]
  PIN la_data_out_core[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 116.000 720.270 122.000 ;
    END
  END la_data_out_core[72]
  PIN la_data_out_core[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 116.000 726.710 122.000 ;
    END
  END la_data_out_core[73]
  PIN la_data_out_core[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 116.000 733.610 122.000 ;
    END
  END la_data_out_core[74]
  PIN la_data_out_core[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 116.000 740.050 122.000 ;
    END
  END la_data_out_core[75]
  PIN la_data_out_core[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 116.000 746.950 122.000 ;
    END
  END la_data_out_core[76]
  PIN la_data_out_core[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 116.000 753.390 122.000 ;
    END
  END la_data_out_core[77]
  PIN la_data_out_core[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 116.000 760.290 122.000 ;
    END
  END la_data_out_core[78]
  PIN la_data_out_core[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 116.000 766.730 122.000 ;
    END
  END la_data_out_core[79]
  PIN la_data_out_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 116.000 286.030 122.000 ;
    END
  END la_data_out_core[7]
  PIN la_data_out_core[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 116.000 773.630 122.000 ;
    END
  END la_data_out_core[80]
  PIN la_data_out_core[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 116.000 780.530 122.000 ;
    END
  END la_data_out_core[81]
  PIN la_data_out_core[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 116.000 786.970 122.000 ;
    END
  END la_data_out_core[82]
  PIN la_data_out_core[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 116.000 793.870 122.000 ;
    END
  END la_data_out_core[83]
  PIN la_data_out_core[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 116.000 800.310 122.000 ;
    END
  END la_data_out_core[84]
  PIN la_data_out_core[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.930 116.000 807.210 122.000 ;
    END
  END la_data_out_core[85]
  PIN la_data_out_core[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 116.000 813.650 122.000 ;
    END
  END la_data_out_core[86]
  PIN la_data_out_core[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 116.000 820.550 122.000 ;
    END
  END la_data_out_core[87]
  PIN la_data_out_core[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 116.000 826.990 122.000 ;
    END
  END la_data_out_core[88]
  PIN la_data_out_core[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 116.000 833.890 122.000 ;
    END
  END la_data_out_core[89]
  PIN la_data_out_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 116.000 292.930 122.000 ;
    END
  END la_data_out_core[8]
  PIN la_data_out_core[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 116.000 840.330 122.000 ;
    END
  END la_data_out_core[90]
  PIN la_data_out_core[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 116.000 847.230 122.000 ;
    END
  END la_data_out_core[91]
  PIN la_data_out_core[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 116.000 853.670 122.000 ;
    END
  END la_data_out_core[92]
  PIN la_data_out_core[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 116.000 860.570 122.000 ;
    END
  END la_data_out_core[93]
  PIN la_data_out_core[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 116.000 867.010 122.000 ;
    END
  END la_data_out_core[94]
  PIN la_data_out_core[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 116.000 873.910 122.000 ;
    END
  END la_data_out_core[95]
  PIN la_data_out_core[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.070 116.000 880.350 122.000 ;
    END
  END la_data_out_core[96]
  PIN la_data_out_core[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.970 116.000 887.250 122.000 ;
    END
  END la_data_out_core[97]
  PIN la_data_out_core[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 116.000 893.690 122.000 ;
    END
  END la_data_out_core[98]
  PIN la_data_out_core[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 116.000 900.590 122.000 ;
    END
  END la_data_out_core[99]
  PIN la_data_out_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 116.000 299.370 122.000 ;
    END
  END la_data_out_core[9]
  PIN la_data_out_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 -2.000 2.210 4.000 ;
    END
  END la_data_out_mprj[0]
  PIN la_data_out_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 -2.000 715.210 4.000 ;
    END
  END la_data_out_mprj[100]
  PIN la_data_out_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 -2.000 722.570 4.000 ;
    END
  END la_data_out_mprj[101]
  PIN la_data_out_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 -2.000 729.470 4.000 ;
    END
  END la_data_out_mprj[102]
  PIN la_data_out_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 -2.000 736.830 4.000 ;
    END
  END la_data_out_mprj[103]
  PIN la_data_out_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 -2.000 743.730 4.000 ;
    END
  END la_data_out_mprj[104]
  PIN la_data_out_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 -2.000 751.090 4.000 ;
    END
  END la_data_out_mprj[105]
  PIN la_data_out_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 -2.000 757.990 4.000 ;
    END
  END la_data_out_mprj[106]
  PIN la_data_out_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.070 -2.000 765.350 4.000 ;
    END
  END la_data_out_mprj[107]
  PIN la_data_out_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 -2.000 772.250 4.000 ;
    END
  END la_data_out_mprj[108]
  PIN la_data_out_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 -2.000 779.610 4.000 ;
    END
  END la_data_out_mprj[109]
  PIN la_data_out_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 -2.000 73.510 4.000 ;
    END
  END la_data_out_mprj[10]
  PIN la_data_out_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 -2.000 786.510 4.000 ;
    END
  END la_data_out_mprj[110]
  PIN la_data_out_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 -2.000 793.870 4.000 ;
    END
  END la_data_out_mprj[111]
  PIN la_data_out_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 -2.000 800.770 4.000 ;
    END
  END la_data_out_mprj[112]
  PIN la_data_out_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 -2.000 808.130 4.000 ;
    END
  END la_data_out_mprj[113]
  PIN la_data_out_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 -2.000 815.030 4.000 ;
    END
  END la_data_out_mprj[114]
  PIN la_data_out_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 -2.000 822.390 4.000 ;
    END
  END la_data_out_mprj[115]
  PIN la_data_out_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 -2.000 829.290 4.000 ;
    END
  END la_data_out_mprj[116]
  PIN la_data_out_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 -2.000 836.650 4.000 ;
    END
  END la_data_out_mprj[117]
  PIN la_data_out_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 -2.000 843.550 4.000 ;
    END
  END la_data_out_mprj[118]
  PIN la_data_out_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 -2.000 850.910 4.000 ;
    END
  END la_data_out_mprj[119]
  PIN la_data_out_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 -2.000 80.870 4.000 ;
    END
  END la_data_out_mprj[11]
  PIN la_data_out_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.530 -2.000 857.810 4.000 ;
    END
  END la_data_out_mprj[120]
  PIN la_data_out_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 -2.000 865.170 4.000 ;
    END
  END la_data_out_mprj[121]
  PIN la_data_out_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 -2.000 872.070 4.000 ;
    END
  END la_data_out_mprj[122]
  PIN la_data_out_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 -2.000 879.430 4.000 ;
    END
  END la_data_out_mprj[123]
  PIN la_data_out_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 -2.000 886.330 4.000 ;
    END
  END la_data_out_mprj[124]
  PIN la_data_out_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 -2.000 893.690 4.000 ;
    END
  END la_data_out_mprj[125]
  PIN la_data_out_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 -2.000 900.590 4.000 ;
    END
  END la_data_out_mprj[126]
  PIN la_data_out_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.670 -2.000 907.950 4.000 ;
    END
  END la_data_out_mprj[127]
  PIN la_data_out_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 -2.000 87.770 4.000 ;
    END
  END la_data_out_mprj[12]
  PIN la_data_out_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 -2.000 95.130 4.000 ;
    END
  END la_data_out_mprj[13]
  PIN la_data_out_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 -2.000 102.030 4.000 ;
    END
  END la_data_out_mprj[14]
  PIN la_data_out_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 -2.000 109.390 4.000 ;
    END
  END la_data_out_mprj[15]
  PIN la_data_out_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 -2.000 116.290 4.000 ;
    END
  END la_data_out_mprj[16]
  PIN la_data_out_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 -2.000 123.650 4.000 ;
    END
  END la_data_out_mprj[17]
  PIN la_data_out_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 -2.000 130.550 4.000 ;
    END
  END la_data_out_mprj[18]
  PIN la_data_out_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 -2.000 137.910 4.000 ;
    END
  END la_data_out_mprj[19]
  PIN la_data_out_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 -2.000 9.570 4.000 ;
    END
  END la_data_out_mprj[1]
  PIN la_data_out_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 -2.000 144.810 4.000 ;
    END
  END la_data_out_mprj[20]
  PIN la_data_out_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 -2.000 152.170 4.000 ;
    END
  END la_data_out_mprj[21]
  PIN la_data_out_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 -2.000 159.070 4.000 ;
    END
  END la_data_out_mprj[22]
  PIN la_data_out_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 -2.000 166.430 4.000 ;
    END
  END la_data_out_mprj[23]
  PIN la_data_out_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 -2.000 173.330 4.000 ;
    END
  END la_data_out_mprj[24]
  PIN la_data_out_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 -2.000 180.690 4.000 ;
    END
  END la_data_out_mprj[25]
  PIN la_data_out_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 -2.000 187.590 4.000 ;
    END
  END la_data_out_mprj[26]
  PIN la_data_out_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 -2.000 194.950 4.000 ;
    END
  END la_data_out_mprj[27]
  PIN la_data_out_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 -2.000 201.850 4.000 ;
    END
  END la_data_out_mprj[28]
  PIN la_data_out_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 -2.000 209.210 4.000 ;
    END
  END la_data_out_mprj[29]
  PIN la_data_out_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 -2.000 16.470 4.000 ;
    END
  END la_data_out_mprj[2]
  PIN la_data_out_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 -2.000 216.110 4.000 ;
    END
  END la_data_out_mprj[30]
  PIN la_data_out_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 -2.000 223.470 4.000 ;
    END
  END la_data_out_mprj[31]
  PIN la_data_out_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 -2.000 230.370 4.000 ;
    END
  END la_data_out_mprj[32]
  PIN la_data_out_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 -2.000 237.730 4.000 ;
    END
  END la_data_out_mprj[33]
  PIN la_data_out_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 -2.000 244.630 4.000 ;
    END
  END la_data_out_mprj[34]
  PIN la_data_out_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 -2.000 251.990 4.000 ;
    END
  END la_data_out_mprj[35]
  PIN la_data_out_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 -2.000 258.890 4.000 ;
    END
  END la_data_out_mprj[36]
  PIN la_data_out_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 -2.000 266.250 4.000 ;
    END
  END la_data_out_mprj[37]
  PIN la_data_out_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 -2.000 273.150 4.000 ;
    END
  END la_data_out_mprj[38]
  PIN la_data_out_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 -2.000 280.510 4.000 ;
    END
  END la_data_out_mprj[39]
  PIN la_data_out_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 -2.000 23.830 4.000 ;
    END
  END la_data_out_mprj[3]
  PIN la_data_out_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 -2.000 287.410 4.000 ;
    END
  END la_data_out_mprj[40]
  PIN la_data_out_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 -2.000 294.770 4.000 ;
    END
  END la_data_out_mprj[41]
  PIN la_data_out_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 -2.000 301.670 4.000 ;
    END
  END la_data_out_mprj[42]
  PIN la_data_out_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 -2.000 309.030 4.000 ;
    END
  END la_data_out_mprj[43]
  PIN la_data_out_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 -2.000 315.930 4.000 ;
    END
  END la_data_out_mprj[44]
  PIN la_data_out_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 -2.000 323.290 4.000 ;
    END
  END la_data_out_mprj[45]
  PIN la_data_out_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 -2.000 330.190 4.000 ;
    END
  END la_data_out_mprj[46]
  PIN la_data_out_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 -2.000 337.550 4.000 ;
    END
  END la_data_out_mprj[47]
  PIN la_data_out_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 -2.000 344.450 4.000 ;
    END
  END la_data_out_mprj[48]
  PIN la_data_out_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 -2.000 351.810 4.000 ;
    END
  END la_data_out_mprj[49]
  PIN la_data_out_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 -2.000 30.730 4.000 ;
    END
  END la_data_out_mprj[4]
  PIN la_data_out_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 -2.000 358.710 4.000 ;
    END
  END la_data_out_mprj[50]
  PIN la_data_out_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 -2.000 366.070 4.000 ;
    END
  END la_data_out_mprj[51]
  PIN la_data_out_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 -2.000 372.970 4.000 ;
    END
  END la_data_out_mprj[52]
  PIN la_data_out_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 -2.000 380.330 4.000 ;
    END
  END la_data_out_mprj[53]
  PIN la_data_out_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 -2.000 387.230 4.000 ;
    END
  END la_data_out_mprj[54]
  PIN la_data_out_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 -2.000 394.590 4.000 ;
    END
  END la_data_out_mprj[55]
  PIN la_data_out_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 -2.000 401.490 4.000 ;
    END
  END la_data_out_mprj[56]
  PIN la_data_out_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 -2.000 408.850 4.000 ;
    END
  END la_data_out_mprj[57]
  PIN la_data_out_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 -2.000 415.750 4.000 ;
    END
  END la_data_out_mprj[58]
  PIN la_data_out_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 -2.000 423.110 4.000 ;
    END
  END la_data_out_mprj[59]
  PIN la_data_out_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 -2.000 38.090 4.000 ;
    END
  END la_data_out_mprj[5]
  PIN la_data_out_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 -2.000 430.010 4.000 ;
    END
  END la_data_out_mprj[60]
  PIN la_data_out_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 -2.000 437.370 4.000 ;
    END
  END la_data_out_mprj[61]
  PIN la_data_out_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 -2.000 444.270 4.000 ;
    END
  END la_data_out_mprj[62]
  PIN la_data_out_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 -2.000 451.630 4.000 ;
    END
  END la_data_out_mprj[63]
  PIN la_data_out_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 -2.000 458.530 4.000 ;
    END
  END la_data_out_mprj[64]
  PIN la_data_out_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 -2.000 465.890 4.000 ;
    END
  END la_data_out_mprj[65]
  PIN la_data_out_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 -2.000 472.790 4.000 ;
    END
  END la_data_out_mprj[66]
  PIN la_data_out_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 -2.000 480.150 4.000 ;
    END
  END la_data_out_mprj[67]
  PIN la_data_out_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 -2.000 487.050 4.000 ;
    END
  END la_data_out_mprj[68]
  PIN la_data_out_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 -2.000 494.410 4.000 ;
    END
  END la_data_out_mprj[69]
  PIN la_data_out_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 -2.000 44.990 4.000 ;
    END
  END la_data_out_mprj[6]
  PIN la_data_out_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 -2.000 501.310 4.000 ;
    END
  END la_data_out_mprj[70]
  PIN la_data_out_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 -2.000 508.670 4.000 ;
    END
  END la_data_out_mprj[71]
  PIN la_data_out_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 -2.000 515.570 4.000 ;
    END
  END la_data_out_mprj[72]
  PIN la_data_out_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 -2.000 522.930 4.000 ;
    END
  END la_data_out_mprj[73]
  PIN la_data_out_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 -2.000 529.830 4.000 ;
    END
  END la_data_out_mprj[74]
  PIN la_data_out_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 -2.000 537.190 4.000 ;
    END
  END la_data_out_mprj[75]
  PIN la_data_out_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 -2.000 544.090 4.000 ;
    END
  END la_data_out_mprj[76]
  PIN la_data_out_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 -2.000 551.450 4.000 ;
    END
  END la_data_out_mprj[77]
  PIN la_data_out_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 -2.000 558.350 4.000 ;
    END
  END la_data_out_mprj[78]
  PIN la_data_out_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 -2.000 565.710 4.000 ;
    END
  END la_data_out_mprj[79]
  PIN la_data_out_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 -2.000 52.350 4.000 ;
    END
  END la_data_out_mprj[7]
  PIN la_data_out_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 -2.000 572.610 4.000 ;
    END
  END la_data_out_mprj[80]
  PIN la_data_out_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 -2.000 579.970 4.000 ;
    END
  END la_data_out_mprj[81]
  PIN la_data_out_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 -2.000 586.870 4.000 ;
    END
  END la_data_out_mprj[82]
  PIN la_data_out_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 -2.000 594.230 4.000 ;
    END
  END la_data_out_mprj[83]
  PIN la_data_out_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 -2.000 601.130 4.000 ;
    END
  END la_data_out_mprj[84]
  PIN la_data_out_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 -2.000 608.490 4.000 ;
    END
  END la_data_out_mprj[85]
  PIN la_data_out_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 -2.000 615.390 4.000 ;
    END
  END la_data_out_mprj[86]
  PIN la_data_out_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 -2.000 622.750 4.000 ;
    END
  END la_data_out_mprj[87]
  PIN la_data_out_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 -2.000 629.650 4.000 ;
    END
  END la_data_out_mprj[88]
  PIN la_data_out_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 -2.000 637.010 4.000 ;
    END
  END la_data_out_mprj[89]
  PIN la_data_out_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 -2.000 59.250 4.000 ;
    END
  END la_data_out_mprj[8]
  PIN la_data_out_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 -2.000 643.910 4.000 ;
    END
  END la_data_out_mprj[90]
  PIN la_data_out_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 -2.000 651.270 4.000 ;
    END
  END la_data_out_mprj[91]
  PIN la_data_out_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 -2.000 658.170 4.000 ;
    END
  END la_data_out_mprj[92]
  PIN la_data_out_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 -2.000 665.530 4.000 ;
    END
  END la_data_out_mprj[93]
  PIN la_data_out_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 -2.000 672.430 4.000 ;
    END
  END la_data_out_mprj[94]
  PIN la_data_out_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 -2.000 679.790 4.000 ;
    END
  END la_data_out_mprj[95]
  PIN la_data_out_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 -2.000 686.690 4.000 ;
    END
  END la_data_out_mprj[96]
  PIN la_data_out_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 -2.000 694.050 4.000 ;
    END
  END la_data_out_mprj[97]
  PIN la_data_out_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 -2.000 700.950 4.000 ;
    END
  END la_data_out_mprj[98]
  PIN la_data_out_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 -2.000 708.310 4.000 ;
    END
  END la_data_out_mprj[99]
  PIN la_data_out_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 -2.000 66.610 4.000 ;
    END
  END la_data_out_mprj[9]
  PIN la_iena_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 -2.000 4.050 4.000 ;
    END
  END la_iena_mprj[0]
  PIN la_iena_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 -2.000 717.050 4.000 ;
    END
  END la_iena_mprj[100]
  PIN la_iena_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 -2.000 724.410 4.000 ;
    END
  END la_iena_mprj[101]
  PIN la_iena_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 -2.000 731.310 4.000 ;
    END
  END la_iena_mprj[102]
  PIN la_iena_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 -2.000 738.670 4.000 ;
    END
  END la_iena_mprj[103]
  PIN la_iena_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 -2.000 745.570 4.000 ;
    END
  END la_iena_mprj[104]
  PIN la_iena_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 -2.000 752.930 4.000 ;
    END
  END la_iena_mprj[105]
  PIN la_iena_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.550 -2.000 759.830 4.000 ;
    END
  END la_iena_mprj[106]
  PIN la_iena_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 -2.000 767.190 4.000 ;
    END
  END la_iena_mprj[107]
  PIN la_iena_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 -2.000 774.090 4.000 ;
    END
  END la_iena_mprj[108]
  PIN la_iena_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 -2.000 781.450 4.000 ;
    END
  END la_iena_mprj[109]
  PIN la_iena_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 -2.000 75.350 4.000 ;
    END
  END la_iena_mprj[10]
  PIN la_iena_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 -2.000 788.350 4.000 ;
    END
  END la_iena_mprj[110]
  PIN la_iena_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 -2.000 795.710 4.000 ;
    END
  END la_iena_mprj[111]
  PIN la_iena_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 -2.000 802.610 4.000 ;
    END
  END la_iena_mprj[112]
  PIN la_iena_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 -2.000 809.970 4.000 ;
    END
  END la_iena_mprj[113]
  PIN la_iena_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.590 -2.000 816.870 4.000 ;
    END
  END la_iena_mprj[114]
  PIN la_iena_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 -2.000 824.230 4.000 ;
    END
  END la_iena_mprj[115]
  PIN la_iena_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 -2.000 831.130 4.000 ;
    END
  END la_iena_mprj[116]
  PIN la_iena_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 -2.000 838.490 4.000 ;
    END
  END la_iena_mprj[117]
  PIN la_iena_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 -2.000 845.390 4.000 ;
    END
  END la_iena_mprj[118]
  PIN la_iena_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 -2.000 852.750 4.000 ;
    END
  END la_iena_mprj[119]
  PIN la_iena_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 -2.000 82.710 4.000 ;
    END
  END la_iena_mprj[11]
  PIN la_iena_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 -2.000 859.650 4.000 ;
    END
  END la_iena_mprj[120]
  PIN la_iena_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 -2.000 867.010 4.000 ;
    END
  END la_iena_mprj[121]
  PIN la_iena_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 -2.000 873.910 4.000 ;
    END
  END la_iena_mprj[122]
  PIN la_iena_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 -2.000 881.270 4.000 ;
    END
  END la_iena_mprj[123]
  PIN la_iena_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 -2.000 888.170 4.000 ;
    END
  END la_iena_mprj[124]
  PIN la_iena_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 -2.000 895.530 4.000 ;
    END
  END la_iena_mprj[125]
  PIN la_iena_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.150 -2.000 902.430 4.000 ;
    END
  END la_iena_mprj[126]
  PIN la_iena_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 -2.000 909.790 4.000 ;
    END
  END la_iena_mprj[127]
  PIN la_iena_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 -2.000 89.610 4.000 ;
    END
  END la_iena_mprj[12]
  PIN la_iena_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 -2.000 96.970 4.000 ;
    END
  END la_iena_mprj[13]
  PIN la_iena_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 -2.000 103.870 4.000 ;
    END
  END la_iena_mprj[14]
  PIN la_iena_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 -2.000 111.230 4.000 ;
    END
  END la_iena_mprj[15]
  PIN la_iena_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 -2.000 118.130 4.000 ;
    END
  END la_iena_mprj[16]
  PIN la_iena_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 -2.000 125.490 4.000 ;
    END
  END la_iena_mprj[17]
  PIN la_iena_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 -2.000 132.390 4.000 ;
    END
  END la_iena_mprj[18]
  PIN la_iena_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 -2.000 139.750 4.000 ;
    END
  END la_iena_mprj[19]
  PIN la_iena_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 -2.000 11.410 4.000 ;
    END
  END la_iena_mprj[1]
  PIN la_iena_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 -2.000 146.650 4.000 ;
    END
  END la_iena_mprj[20]
  PIN la_iena_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 -2.000 154.010 4.000 ;
    END
  END la_iena_mprj[21]
  PIN la_iena_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 -2.000 160.910 4.000 ;
    END
  END la_iena_mprj[22]
  PIN la_iena_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 -2.000 168.270 4.000 ;
    END
  END la_iena_mprj[23]
  PIN la_iena_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 -2.000 175.170 4.000 ;
    END
  END la_iena_mprj[24]
  PIN la_iena_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 -2.000 182.530 4.000 ;
    END
  END la_iena_mprj[25]
  PIN la_iena_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 -2.000 189.430 4.000 ;
    END
  END la_iena_mprj[26]
  PIN la_iena_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 -2.000 196.790 4.000 ;
    END
  END la_iena_mprj[27]
  PIN la_iena_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 -2.000 203.690 4.000 ;
    END
  END la_iena_mprj[28]
  PIN la_iena_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 -2.000 211.050 4.000 ;
    END
  END la_iena_mprj[29]
  PIN la_iena_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 -2.000 18.310 4.000 ;
    END
  END la_iena_mprj[2]
  PIN la_iena_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 -2.000 217.950 4.000 ;
    END
  END la_iena_mprj[30]
  PIN la_iena_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 -2.000 225.310 4.000 ;
    END
  END la_iena_mprj[31]
  PIN la_iena_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 -2.000 232.210 4.000 ;
    END
  END la_iena_mprj[32]
  PIN la_iena_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 -2.000 239.570 4.000 ;
    END
  END la_iena_mprj[33]
  PIN la_iena_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 -2.000 246.470 4.000 ;
    END
  END la_iena_mprj[34]
  PIN la_iena_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 -2.000 253.830 4.000 ;
    END
  END la_iena_mprj[35]
  PIN la_iena_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 -2.000 260.730 4.000 ;
    END
  END la_iena_mprj[36]
  PIN la_iena_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 -2.000 268.090 4.000 ;
    END
  END la_iena_mprj[37]
  PIN la_iena_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 -2.000 274.990 4.000 ;
    END
  END la_iena_mprj[38]
  PIN la_iena_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 -2.000 282.350 4.000 ;
    END
  END la_iena_mprj[39]
  PIN la_iena_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 -2.000 25.670 4.000 ;
    END
  END la_iena_mprj[3]
  PIN la_iena_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 -2.000 289.250 4.000 ;
    END
  END la_iena_mprj[40]
  PIN la_iena_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 -2.000 296.610 4.000 ;
    END
  END la_iena_mprj[41]
  PIN la_iena_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 -2.000 303.510 4.000 ;
    END
  END la_iena_mprj[42]
  PIN la_iena_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 -2.000 310.870 4.000 ;
    END
  END la_iena_mprj[43]
  PIN la_iena_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 -2.000 317.770 4.000 ;
    END
  END la_iena_mprj[44]
  PIN la_iena_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 -2.000 325.130 4.000 ;
    END
  END la_iena_mprj[45]
  PIN la_iena_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 -2.000 332.030 4.000 ;
    END
  END la_iena_mprj[46]
  PIN la_iena_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 -2.000 339.390 4.000 ;
    END
  END la_iena_mprj[47]
  PIN la_iena_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 -2.000 346.290 4.000 ;
    END
  END la_iena_mprj[48]
  PIN la_iena_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 -2.000 353.650 4.000 ;
    END
  END la_iena_mprj[49]
  PIN la_iena_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 -2.000 32.570 4.000 ;
    END
  END la_iena_mprj[4]
  PIN la_iena_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 -2.000 360.550 4.000 ;
    END
  END la_iena_mprj[50]
  PIN la_iena_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 -2.000 367.910 4.000 ;
    END
  END la_iena_mprj[51]
  PIN la_iena_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 -2.000 374.810 4.000 ;
    END
  END la_iena_mprj[52]
  PIN la_iena_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 -2.000 382.170 4.000 ;
    END
  END la_iena_mprj[53]
  PIN la_iena_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 -2.000 389.070 4.000 ;
    END
  END la_iena_mprj[54]
  PIN la_iena_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 -2.000 396.430 4.000 ;
    END
  END la_iena_mprj[55]
  PIN la_iena_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 -2.000 403.330 4.000 ;
    END
  END la_iena_mprj[56]
  PIN la_iena_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 -2.000 410.690 4.000 ;
    END
  END la_iena_mprj[57]
  PIN la_iena_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 -2.000 417.590 4.000 ;
    END
  END la_iena_mprj[58]
  PIN la_iena_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 -2.000 424.950 4.000 ;
    END
  END la_iena_mprj[59]
  PIN la_iena_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 -2.000 39.930 4.000 ;
    END
  END la_iena_mprj[5]
  PIN la_iena_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 -2.000 431.850 4.000 ;
    END
  END la_iena_mprj[60]
  PIN la_iena_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 -2.000 439.210 4.000 ;
    END
  END la_iena_mprj[61]
  PIN la_iena_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 -2.000 446.110 4.000 ;
    END
  END la_iena_mprj[62]
  PIN la_iena_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 -2.000 453.470 4.000 ;
    END
  END la_iena_mprj[63]
  PIN la_iena_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 -2.000 460.370 4.000 ;
    END
  END la_iena_mprj[64]
  PIN la_iena_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 -2.000 467.730 4.000 ;
    END
  END la_iena_mprj[65]
  PIN la_iena_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 -2.000 474.630 4.000 ;
    END
  END la_iena_mprj[66]
  PIN la_iena_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 -2.000 481.990 4.000 ;
    END
  END la_iena_mprj[67]
  PIN la_iena_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 -2.000 488.890 4.000 ;
    END
  END la_iena_mprj[68]
  PIN la_iena_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 -2.000 496.250 4.000 ;
    END
  END la_iena_mprj[69]
  PIN la_iena_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 -2.000 46.830 4.000 ;
    END
  END la_iena_mprj[6]
  PIN la_iena_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 -2.000 503.150 4.000 ;
    END
  END la_iena_mprj[70]
  PIN la_iena_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 -2.000 510.510 4.000 ;
    END
  END la_iena_mprj[71]
  PIN la_iena_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 -2.000 517.410 4.000 ;
    END
  END la_iena_mprj[72]
  PIN la_iena_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 -2.000 524.770 4.000 ;
    END
  END la_iena_mprj[73]
  PIN la_iena_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 -2.000 531.670 4.000 ;
    END
  END la_iena_mprj[74]
  PIN la_iena_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 -2.000 539.030 4.000 ;
    END
  END la_iena_mprj[75]
  PIN la_iena_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 -2.000 545.930 4.000 ;
    END
  END la_iena_mprj[76]
  PIN la_iena_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 -2.000 553.290 4.000 ;
    END
  END la_iena_mprj[77]
  PIN la_iena_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 -2.000 560.190 4.000 ;
    END
  END la_iena_mprj[78]
  PIN la_iena_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 -2.000 567.550 4.000 ;
    END
  END la_iena_mprj[79]
  PIN la_iena_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 -2.000 54.190 4.000 ;
    END
  END la_iena_mprj[7]
  PIN la_iena_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 -2.000 574.450 4.000 ;
    END
  END la_iena_mprj[80]
  PIN la_iena_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 -2.000 581.810 4.000 ;
    END
  END la_iena_mprj[81]
  PIN la_iena_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 -2.000 588.710 4.000 ;
    END
  END la_iena_mprj[82]
  PIN la_iena_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 -2.000 596.070 4.000 ;
    END
  END la_iena_mprj[83]
  PIN la_iena_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 -2.000 602.970 4.000 ;
    END
  END la_iena_mprj[84]
  PIN la_iena_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 -2.000 610.330 4.000 ;
    END
  END la_iena_mprj[85]
  PIN la_iena_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 -2.000 617.230 4.000 ;
    END
  END la_iena_mprj[86]
  PIN la_iena_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 -2.000 624.590 4.000 ;
    END
  END la_iena_mprj[87]
  PIN la_iena_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 -2.000 631.490 4.000 ;
    END
  END la_iena_mprj[88]
  PIN la_iena_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 -2.000 638.850 4.000 ;
    END
  END la_iena_mprj[89]
  PIN la_iena_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 -2.000 61.090 4.000 ;
    END
  END la_iena_mprj[8]
  PIN la_iena_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 -2.000 645.750 4.000 ;
    END
  END la_iena_mprj[90]
  PIN la_iena_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 -2.000 653.110 4.000 ;
    END
  END la_iena_mprj[91]
  PIN la_iena_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 -2.000 660.010 4.000 ;
    END
  END la_iena_mprj[92]
  PIN la_iena_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 -2.000 667.370 4.000 ;
    END
  END la_iena_mprj[93]
  PIN la_iena_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 -2.000 674.270 4.000 ;
    END
  END la_iena_mprj[94]
  PIN la_iena_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 -2.000 681.630 4.000 ;
    END
  END la_iena_mprj[95]
  PIN la_iena_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 -2.000 688.530 4.000 ;
    END
  END la_iena_mprj[96]
  PIN la_iena_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 -2.000 695.890 4.000 ;
    END
  END la_iena_mprj[97]
  PIN la_iena_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 -2.000 702.790 4.000 ;
    END
  END la_iena_mprj[98]
  PIN la_iena_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.870 -2.000 710.150 4.000 ;
    END
  END la_iena_mprj[99]
  PIN la_iena_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 -2.000 68.450 4.000 ;
    END
  END la_iena_mprj[9]
  PIN la_oenb_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 116.000 241.410 122.000 ;
    END
  END la_oenb_core[0]
  PIN la_oenb_core[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.050 116.000 909.330 122.000 ;
    END
  END la_oenb_core[100]
  PIN la_oenb_core[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 116.000 916.230 122.000 ;
    END
  END la_oenb_core[101]
  PIN la_oenb_core[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 116.000 922.670 122.000 ;
    END
  END la_oenb_core[102]
  PIN la_oenb_core[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 116.000 929.570 122.000 ;
    END
  END la_oenb_core[103]
  PIN la_oenb_core[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730 116.000 936.010 122.000 ;
    END
  END la_oenb_core[104]
  PIN la_oenb_core[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 116.000 942.910 122.000 ;
    END
  END la_oenb_core[105]
  PIN la_oenb_core[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 116.000 949.350 122.000 ;
    END
  END la_oenb_core[106]
  PIN la_oenb_core[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.970 116.000 956.250 122.000 ;
    END
  END la_oenb_core[107]
  PIN la_oenb_core[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.410 116.000 962.690 122.000 ;
    END
  END la_oenb_core[108]
  PIN la_oenb_core[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 116.000 969.590 122.000 ;
    END
  END la_oenb_core[109]
  PIN la_oenb_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 116.000 308.110 122.000 ;
    END
  END la_oenb_core[10]
  PIN la_oenb_core[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 116.000 976.030 122.000 ;
    END
  END la_oenb_core[110]
  PIN la_oenb_core[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 116.000 982.930 122.000 ;
    END
  END la_oenb_core[111]
  PIN la_oenb_core[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.090 116.000 989.370 122.000 ;
    END
  END la_oenb_core[112]
  PIN la_oenb_core[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 116.000 996.270 122.000 ;
    END
  END la_oenb_core[113]
  PIN la_oenb_core[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 116.000 1003.170 122.000 ;
    END
  END la_oenb_core[114]
  PIN la_oenb_core[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.330 116.000 1009.610 122.000 ;
    END
  END la_oenb_core[115]
  PIN la_oenb_core[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.230 116.000 1016.510 122.000 ;
    END
  END la_oenb_core[116]
  PIN la_oenb_core[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.670 116.000 1022.950 122.000 ;
    END
  END la_oenb_core[117]
  PIN la_oenb_core[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.570 116.000 1029.850 122.000 ;
    END
  END la_oenb_core[118]
  PIN la_oenb_core[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 116.000 1036.290 122.000 ;
    END
  END la_oenb_core[119]
  PIN la_oenb_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 116.000 315.010 122.000 ;
    END
  END la_oenb_core[11]
  PIN la_oenb_core[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.910 116.000 1043.190 122.000 ;
    END
  END la_oenb_core[120]
  PIN la_oenb_core[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.350 116.000 1049.630 122.000 ;
    END
  END la_oenb_core[121]
  PIN la_oenb_core[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 116.000 1056.530 122.000 ;
    END
  END la_oenb_core[122]
  PIN la_oenb_core[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 116.000 1062.970 122.000 ;
    END
  END la_oenb_core[123]
  PIN la_oenb_core[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 116.000 1069.870 122.000 ;
    END
  END la_oenb_core[124]
  PIN la_oenb_core[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.030 116.000 1076.310 122.000 ;
    END
  END la_oenb_core[125]
  PIN la_oenb_core[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 116.000 1083.210 122.000 ;
    END
  END la_oenb_core[126]
  PIN la_oenb_core[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 116.000 1089.650 122.000 ;
    END
  END la_oenb_core[127]
  PIN la_oenb_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 116.000 321.450 122.000 ;
    END
  END la_oenb_core[12]
  PIN la_oenb_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 116.000 328.350 122.000 ;
    END
  END la_oenb_core[13]
  PIN la_oenb_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 116.000 335.250 122.000 ;
    END
  END la_oenb_core[14]
  PIN la_oenb_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 116.000 341.690 122.000 ;
    END
  END la_oenb_core[15]
  PIN la_oenb_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 116.000 348.590 122.000 ;
    END
  END la_oenb_core[16]
  PIN la_oenb_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 116.000 355.030 122.000 ;
    END
  END la_oenb_core[17]
  PIN la_oenb_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 116.000 361.930 122.000 ;
    END
  END la_oenb_core[18]
  PIN la_oenb_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 116.000 368.370 122.000 ;
    END
  END la_oenb_core[19]
  PIN la_oenb_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 116.000 248.310 122.000 ;
    END
  END la_oenb_core[1]
  PIN la_oenb_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 116.000 375.270 122.000 ;
    END
  END la_oenb_core[20]
  PIN la_oenb_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 116.000 381.710 122.000 ;
    END
  END la_oenb_core[21]
  PIN la_oenb_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 116.000 388.610 122.000 ;
    END
  END la_oenb_core[22]
  PIN la_oenb_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 116.000 395.050 122.000 ;
    END
  END la_oenb_core[23]
  PIN la_oenb_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 116.000 401.950 122.000 ;
    END
  END la_oenb_core[24]
  PIN la_oenb_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 116.000 408.390 122.000 ;
    END
  END la_oenb_core[25]
  PIN la_oenb_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 116.000 415.290 122.000 ;
    END
  END la_oenb_core[26]
  PIN la_oenb_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 116.000 421.730 122.000 ;
    END
  END la_oenb_core[27]
  PIN la_oenb_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 116.000 428.630 122.000 ;
    END
  END la_oenb_core[28]
  PIN la_oenb_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 116.000 435.070 122.000 ;
    END
  END la_oenb_core[29]
  PIN la_oenb_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 116.000 254.750 122.000 ;
    END
  END la_oenb_core[2]
  PIN la_oenb_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 116.000 441.970 122.000 ;
    END
  END la_oenb_core[30]
  PIN la_oenb_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 116.000 448.410 122.000 ;
    END
  END la_oenb_core[31]
  PIN la_oenb_core[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 116.000 455.310 122.000 ;
    END
  END la_oenb_core[32]
  PIN la_oenb_core[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 116.000 461.750 122.000 ;
    END
  END la_oenb_core[33]
  PIN la_oenb_core[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 116.000 468.650 122.000 ;
    END
  END la_oenb_core[34]
  PIN la_oenb_core[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 116.000 475.090 122.000 ;
    END
  END la_oenb_core[35]
  PIN la_oenb_core[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 116.000 481.990 122.000 ;
    END
  END la_oenb_core[36]
  PIN la_oenb_core[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 116.000 488.430 122.000 ;
    END
  END la_oenb_core[37]
  PIN la_oenb_core[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 116.000 495.330 122.000 ;
    END
  END la_oenb_core[38]
  PIN la_oenb_core[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 116.000 502.230 122.000 ;
    END
  END la_oenb_core[39]
  PIN la_oenb_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 116.000 261.650 122.000 ;
    END
  END la_oenb_core[3]
  PIN la_oenb_core[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 116.000 508.670 122.000 ;
    END
  END la_oenb_core[40]
  PIN la_oenb_core[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 116.000 515.570 122.000 ;
    END
  END la_oenb_core[41]
  PIN la_oenb_core[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 116.000 522.010 122.000 ;
    END
  END la_oenb_core[42]
  PIN la_oenb_core[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 116.000 528.910 122.000 ;
    END
  END la_oenb_core[43]
  PIN la_oenb_core[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 116.000 535.350 122.000 ;
    END
  END la_oenb_core[44]
  PIN la_oenb_core[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 116.000 542.250 122.000 ;
    END
  END la_oenb_core[45]
  PIN la_oenb_core[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 116.000 548.690 122.000 ;
    END
  END la_oenb_core[46]
  PIN la_oenb_core[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 116.000 555.590 122.000 ;
    END
  END la_oenb_core[47]
  PIN la_oenb_core[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 116.000 562.030 122.000 ;
    END
  END la_oenb_core[48]
  PIN la_oenb_core[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 116.000 568.930 122.000 ;
    END
  END la_oenb_core[49]
  PIN la_oenb_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 116.000 268.090 122.000 ;
    END
  END la_oenb_core[4]
  PIN la_oenb_core[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 116.000 575.370 122.000 ;
    END
  END la_oenb_core[50]
  PIN la_oenb_core[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 116.000 582.270 122.000 ;
    END
  END la_oenb_core[51]
  PIN la_oenb_core[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 116.000 588.710 122.000 ;
    END
  END la_oenb_core[52]
  PIN la_oenb_core[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 116.000 595.610 122.000 ;
    END
  END la_oenb_core[53]
  PIN la_oenb_core[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 116.000 602.050 122.000 ;
    END
  END la_oenb_core[54]
  PIN la_oenb_core[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 116.000 608.950 122.000 ;
    END
  END la_oenb_core[55]
  PIN la_oenb_core[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 116.000 615.390 122.000 ;
    END
  END la_oenb_core[56]
  PIN la_oenb_core[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 116.000 622.290 122.000 ;
    END
  END la_oenb_core[57]
  PIN la_oenb_core[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 116.000 628.730 122.000 ;
    END
  END la_oenb_core[58]
  PIN la_oenb_core[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 116.000 635.630 122.000 ;
    END
  END la_oenb_core[59]
  PIN la_oenb_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 116.000 274.990 122.000 ;
    END
  END la_oenb_core[5]
  PIN la_oenb_core[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 116.000 642.070 122.000 ;
    END
  END la_oenb_core[60]
  PIN la_oenb_core[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 116.000 648.970 122.000 ;
    END
  END la_oenb_core[61]
  PIN la_oenb_core[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 116.000 655.410 122.000 ;
    END
  END la_oenb_core[62]
  PIN la_oenb_core[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 116.000 662.310 122.000 ;
    END
  END la_oenb_core[63]
  PIN la_oenb_core[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 116.000 669.210 122.000 ;
    END
  END la_oenb_core[64]
  PIN la_oenb_core[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 116.000 675.650 122.000 ;
    END
  END la_oenb_core[65]
  PIN la_oenb_core[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 116.000 682.550 122.000 ;
    END
  END la_oenb_core[66]
  PIN la_oenb_core[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 116.000 688.990 122.000 ;
    END
  END la_oenb_core[67]
  PIN la_oenb_core[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 116.000 695.890 122.000 ;
    END
  END la_oenb_core[68]
  PIN la_oenb_core[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 116.000 702.330 122.000 ;
    END
  END la_oenb_core[69]
  PIN la_oenb_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 116.000 281.430 122.000 ;
    END
  END la_oenb_core[6]
  PIN la_oenb_core[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 116.000 709.230 122.000 ;
    END
  END la_oenb_core[70]
  PIN la_oenb_core[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 116.000 715.670 122.000 ;
    END
  END la_oenb_core[71]
  PIN la_oenb_core[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 116.000 722.570 122.000 ;
    END
  END la_oenb_core[72]
  PIN la_oenb_core[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 116.000 729.010 122.000 ;
    END
  END la_oenb_core[73]
  PIN la_oenb_core[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 116.000 735.910 122.000 ;
    END
  END la_oenb_core[74]
  PIN la_oenb_core[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 116.000 742.350 122.000 ;
    END
  END la_oenb_core[75]
  PIN la_oenb_core[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 116.000 749.250 122.000 ;
    END
  END la_oenb_core[76]
  PIN la_oenb_core[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 116.000 755.690 122.000 ;
    END
  END la_oenb_core[77]
  PIN la_oenb_core[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 116.000 762.590 122.000 ;
    END
  END la_oenb_core[78]
  PIN la_oenb_core[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 116.000 769.030 122.000 ;
    END
  END la_oenb_core[79]
  PIN la_oenb_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 116.000 288.330 122.000 ;
    END
  END la_oenb_core[7]
  PIN la_oenb_core[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 116.000 775.930 122.000 ;
    END
  END la_oenb_core[80]
  PIN la_oenb_core[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 116.000 782.370 122.000 ;
    END
  END la_oenb_core[81]
  PIN la_oenb_core[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 116.000 789.270 122.000 ;
    END
  END la_oenb_core[82]
  PIN la_oenb_core[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 116.000 795.710 122.000 ;
    END
  END la_oenb_core[83]
  PIN la_oenb_core[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 116.000 802.610 122.000 ;
    END
  END la_oenb_core[84]
  PIN la_oenb_core[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 116.000 809.050 122.000 ;
    END
  END la_oenb_core[85]
  PIN la_oenb_core[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 116.000 815.950 122.000 ;
    END
  END la_oenb_core[86]
  PIN la_oenb_core[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 116.000 822.390 122.000 ;
    END
  END la_oenb_core[87]
  PIN la_oenb_core[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 116.000 829.290 122.000 ;
    END
  END la_oenb_core[88]
  PIN la_oenb_core[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.910 116.000 836.190 122.000 ;
    END
  END la_oenb_core[89]
  PIN la_oenb_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 116.000 294.770 122.000 ;
    END
  END la_oenb_core[8]
  PIN la_oenb_core[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 116.000 842.630 122.000 ;
    END
  END la_oenb_core[90]
  PIN la_oenb_core[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.250 116.000 849.530 122.000 ;
    END
  END la_oenb_core[91]
  PIN la_oenb_core[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 116.000 855.970 122.000 ;
    END
  END la_oenb_core[92]
  PIN la_oenb_core[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 116.000 862.870 122.000 ;
    END
  END la_oenb_core[93]
  PIN la_oenb_core[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.030 116.000 869.310 122.000 ;
    END
  END la_oenb_core[94]
  PIN la_oenb_core[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 116.000 876.210 122.000 ;
    END
  END la_oenb_core[95]
  PIN la_oenb_core[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 116.000 882.650 122.000 ;
    END
  END la_oenb_core[96]
  PIN la_oenb_core[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 116.000 889.550 122.000 ;
    END
  END la_oenb_core[97]
  PIN la_oenb_core[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 116.000 895.990 122.000 ;
    END
  END la_oenb_core[98]
  PIN la_oenb_core[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 116.000 902.890 122.000 ;
    END
  END la_oenb_core[99]
  PIN la_oenb_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 116.000 301.670 122.000 ;
    END
  END la_oenb_core[9]
  PIN la_oenb_mprj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 -2.000 5.890 4.000 ;
    END
  END la_oenb_mprj[0]
  PIN la_oenb_mprj[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 -2.000 718.890 4.000 ;
    END
  END la_oenb_mprj[100]
  PIN la_oenb_mprj[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 -2.000 726.250 4.000 ;
    END
  END la_oenb_mprj[101]
  PIN la_oenb_mprj[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 -2.000 733.150 4.000 ;
    END
  END la_oenb_mprj[102]
  PIN la_oenb_mprj[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 -2.000 740.510 4.000 ;
    END
  END la_oenb_mprj[103]
  PIN la_oenb_mprj[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 -2.000 747.410 4.000 ;
    END
  END la_oenb_mprj[104]
  PIN la_oenb_mprj[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 -2.000 754.770 4.000 ;
    END
  END la_oenb_mprj[105]
  PIN la_oenb_mprj[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 -2.000 761.670 4.000 ;
    END
  END la_oenb_mprj[106]
  PIN la_oenb_mprj[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 -2.000 769.030 4.000 ;
    END
  END la_oenb_mprj[107]
  PIN la_oenb_mprj[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 -2.000 775.930 4.000 ;
    END
  END la_oenb_mprj[108]
  PIN la_oenb_mprj[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 -2.000 783.290 4.000 ;
    END
  END la_oenb_mprj[109]
  PIN la_oenb_mprj[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 -2.000 77.190 4.000 ;
    END
  END la_oenb_mprj[10]
  PIN la_oenb_mprj[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 -2.000 790.190 4.000 ;
    END
  END la_oenb_mprj[110]
  PIN la_oenb_mprj[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 -2.000 797.550 4.000 ;
    END
  END la_oenb_mprj[111]
  PIN la_oenb_mprj[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 -2.000 804.450 4.000 ;
    END
  END la_oenb_mprj[112]
  PIN la_oenb_mprj[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 -2.000 811.810 4.000 ;
    END
  END la_oenb_mprj[113]
  PIN la_oenb_mprj[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 -2.000 818.710 4.000 ;
    END
  END la_oenb_mprj[114]
  PIN la_oenb_mprj[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 -2.000 826.070 4.000 ;
    END
  END la_oenb_mprj[115]
  PIN la_oenb_mprj[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 -2.000 832.970 4.000 ;
    END
  END la_oenb_mprj[116]
  PIN la_oenb_mprj[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 -2.000 840.330 4.000 ;
    END
  END la_oenb_mprj[117]
  PIN la_oenb_mprj[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 -2.000 847.230 4.000 ;
    END
  END la_oenb_mprj[118]
  PIN la_oenb_mprj[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.310 -2.000 854.590 4.000 ;
    END
  END la_oenb_mprj[119]
  PIN la_oenb_mprj[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 -2.000 84.550 4.000 ;
    END
  END la_oenb_mprj[11]
  PIN la_oenb_mprj[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 -2.000 861.490 4.000 ;
    END
  END la_oenb_mprj[120]
  PIN la_oenb_mprj[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.570 -2.000 868.850 4.000 ;
    END
  END la_oenb_mprj[121]
  PIN la_oenb_mprj[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.470 -2.000 875.750 4.000 ;
    END
  END la_oenb_mprj[122]
  PIN la_oenb_mprj[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 -2.000 883.110 4.000 ;
    END
  END la_oenb_mprj[123]
  PIN la_oenb_mprj[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 -2.000 890.010 4.000 ;
    END
  END la_oenb_mprj[124]
  PIN la_oenb_mprj[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 -2.000 897.370 4.000 ;
    END
  END la_oenb_mprj[125]
  PIN la_oenb_mprj[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 -2.000 904.270 4.000 ;
    END
  END la_oenb_mprj[126]
  PIN la_oenb_mprj[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 -2.000 911.630 4.000 ;
    END
  END la_oenb_mprj[127]
  PIN la_oenb_mprj[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 -2.000 91.450 4.000 ;
    END
  END la_oenb_mprj[12]
  PIN la_oenb_mprj[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 -2.000 98.810 4.000 ;
    END
  END la_oenb_mprj[13]
  PIN la_oenb_mprj[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 -2.000 105.710 4.000 ;
    END
  END la_oenb_mprj[14]
  PIN la_oenb_mprj[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 -2.000 113.070 4.000 ;
    END
  END la_oenb_mprj[15]
  PIN la_oenb_mprj[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 -2.000 119.970 4.000 ;
    END
  END la_oenb_mprj[16]
  PIN la_oenb_mprj[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 -2.000 127.330 4.000 ;
    END
  END la_oenb_mprj[17]
  PIN la_oenb_mprj[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 -2.000 134.230 4.000 ;
    END
  END la_oenb_mprj[18]
  PIN la_oenb_mprj[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 -2.000 141.590 4.000 ;
    END
  END la_oenb_mprj[19]
  PIN la_oenb_mprj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 -2.000 13.250 4.000 ;
    END
  END la_oenb_mprj[1]
  PIN la_oenb_mprj[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 -2.000 148.490 4.000 ;
    END
  END la_oenb_mprj[20]
  PIN la_oenb_mprj[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 -2.000 155.850 4.000 ;
    END
  END la_oenb_mprj[21]
  PIN la_oenb_mprj[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 -2.000 162.750 4.000 ;
    END
  END la_oenb_mprj[22]
  PIN la_oenb_mprj[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 -2.000 170.110 4.000 ;
    END
  END la_oenb_mprj[23]
  PIN la_oenb_mprj[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 -2.000 177.010 4.000 ;
    END
  END la_oenb_mprj[24]
  PIN la_oenb_mprj[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 -2.000 184.370 4.000 ;
    END
  END la_oenb_mprj[25]
  PIN la_oenb_mprj[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 -2.000 191.270 4.000 ;
    END
  END la_oenb_mprj[26]
  PIN la_oenb_mprj[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 -2.000 198.630 4.000 ;
    END
  END la_oenb_mprj[27]
  PIN la_oenb_mprj[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 -2.000 205.530 4.000 ;
    END
  END la_oenb_mprj[28]
  PIN la_oenb_mprj[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 -2.000 212.890 4.000 ;
    END
  END la_oenb_mprj[29]
  PIN la_oenb_mprj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 -2.000 20.150 4.000 ;
    END
  END la_oenb_mprj[2]
  PIN la_oenb_mprj[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 -2.000 219.790 4.000 ;
    END
  END la_oenb_mprj[30]
  PIN la_oenb_mprj[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 -2.000 227.150 4.000 ;
    END
  END la_oenb_mprj[31]
  PIN la_oenb_mprj[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 -2.000 234.050 4.000 ;
    END
  END la_oenb_mprj[32]
  PIN la_oenb_mprj[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 -2.000 241.410 4.000 ;
    END
  END la_oenb_mprj[33]
  PIN la_oenb_mprj[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 -2.000 248.310 4.000 ;
    END
  END la_oenb_mprj[34]
  PIN la_oenb_mprj[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 -2.000 255.670 4.000 ;
    END
  END la_oenb_mprj[35]
  PIN la_oenb_mprj[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 -2.000 262.570 4.000 ;
    END
  END la_oenb_mprj[36]
  PIN la_oenb_mprj[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 -2.000 269.930 4.000 ;
    END
  END la_oenb_mprj[37]
  PIN la_oenb_mprj[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 -2.000 276.830 4.000 ;
    END
  END la_oenb_mprj[38]
  PIN la_oenb_mprj[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 -2.000 284.190 4.000 ;
    END
  END la_oenb_mprj[39]
  PIN la_oenb_mprj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 -2.000 27.510 4.000 ;
    END
  END la_oenb_mprj[3]
  PIN la_oenb_mprj[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 -2.000 291.090 4.000 ;
    END
  END la_oenb_mprj[40]
  PIN la_oenb_mprj[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 -2.000 298.450 4.000 ;
    END
  END la_oenb_mprj[41]
  PIN la_oenb_mprj[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 -2.000 305.350 4.000 ;
    END
  END la_oenb_mprj[42]
  PIN la_oenb_mprj[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 -2.000 312.710 4.000 ;
    END
  END la_oenb_mprj[43]
  PIN la_oenb_mprj[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 -2.000 319.610 4.000 ;
    END
  END la_oenb_mprj[44]
  PIN la_oenb_mprj[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 -2.000 326.970 4.000 ;
    END
  END la_oenb_mprj[45]
  PIN la_oenb_mprj[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 -2.000 333.870 4.000 ;
    END
  END la_oenb_mprj[46]
  PIN la_oenb_mprj[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 -2.000 341.230 4.000 ;
    END
  END la_oenb_mprj[47]
  PIN la_oenb_mprj[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 -2.000 348.130 4.000 ;
    END
  END la_oenb_mprj[48]
  PIN la_oenb_mprj[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 -2.000 355.490 4.000 ;
    END
  END la_oenb_mprj[49]
  PIN la_oenb_mprj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 -2.000 34.410 4.000 ;
    END
  END la_oenb_mprj[4]
  PIN la_oenb_mprj[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 -2.000 362.390 4.000 ;
    END
  END la_oenb_mprj[50]
  PIN la_oenb_mprj[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 -2.000 369.750 4.000 ;
    END
  END la_oenb_mprj[51]
  PIN la_oenb_mprj[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 -2.000 376.650 4.000 ;
    END
  END la_oenb_mprj[52]
  PIN la_oenb_mprj[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 -2.000 384.010 4.000 ;
    END
  END la_oenb_mprj[53]
  PIN la_oenb_mprj[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 -2.000 390.910 4.000 ;
    END
  END la_oenb_mprj[54]
  PIN la_oenb_mprj[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 -2.000 398.270 4.000 ;
    END
  END la_oenb_mprj[55]
  PIN la_oenb_mprj[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 -2.000 405.170 4.000 ;
    END
  END la_oenb_mprj[56]
  PIN la_oenb_mprj[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 -2.000 412.530 4.000 ;
    END
  END la_oenb_mprj[57]
  PIN la_oenb_mprj[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 -2.000 419.430 4.000 ;
    END
  END la_oenb_mprj[58]
  PIN la_oenb_mprj[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 -2.000 426.790 4.000 ;
    END
  END la_oenb_mprj[59]
  PIN la_oenb_mprj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 -2.000 41.770 4.000 ;
    END
  END la_oenb_mprj[5]
  PIN la_oenb_mprj[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 -2.000 433.690 4.000 ;
    END
  END la_oenb_mprj[60]
  PIN la_oenb_mprj[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 -2.000 441.050 4.000 ;
    END
  END la_oenb_mprj[61]
  PIN la_oenb_mprj[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 -2.000 447.950 4.000 ;
    END
  END la_oenb_mprj[62]
  PIN la_oenb_mprj[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 -2.000 455.310 4.000 ;
    END
  END la_oenb_mprj[63]
  PIN la_oenb_mprj[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 -2.000 462.210 4.000 ;
    END
  END la_oenb_mprj[64]
  PIN la_oenb_mprj[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 -2.000 469.570 4.000 ;
    END
  END la_oenb_mprj[65]
  PIN la_oenb_mprj[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 -2.000 476.470 4.000 ;
    END
  END la_oenb_mprj[66]
  PIN la_oenb_mprj[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 -2.000 483.830 4.000 ;
    END
  END la_oenb_mprj[67]
  PIN la_oenb_mprj[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 -2.000 490.730 4.000 ;
    END
  END la_oenb_mprj[68]
  PIN la_oenb_mprj[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 -2.000 498.090 4.000 ;
    END
  END la_oenb_mprj[69]
  PIN la_oenb_mprj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 -2.000 48.670 4.000 ;
    END
  END la_oenb_mprj[6]
  PIN la_oenb_mprj[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 -2.000 504.990 4.000 ;
    END
  END la_oenb_mprj[70]
  PIN la_oenb_mprj[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 -2.000 512.350 4.000 ;
    END
  END la_oenb_mprj[71]
  PIN la_oenb_mprj[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 -2.000 519.250 4.000 ;
    END
  END la_oenb_mprj[72]
  PIN la_oenb_mprj[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 -2.000 526.610 4.000 ;
    END
  END la_oenb_mprj[73]
  PIN la_oenb_mprj[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 -2.000 533.510 4.000 ;
    END
  END la_oenb_mprj[74]
  PIN la_oenb_mprj[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 -2.000 540.870 4.000 ;
    END
  END la_oenb_mprj[75]
  PIN la_oenb_mprj[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 -2.000 547.770 4.000 ;
    END
  END la_oenb_mprj[76]
  PIN la_oenb_mprj[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 -2.000 555.130 4.000 ;
    END
  END la_oenb_mprj[77]
  PIN la_oenb_mprj[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 -2.000 562.030 4.000 ;
    END
  END la_oenb_mprj[78]
  PIN la_oenb_mprj[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 -2.000 569.390 4.000 ;
    END
  END la_oenb_mprj[79]
  PIN la_oenb_mprj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 -2.000 56.030 4.000 ;
    END
  END la_oenb_mprj[7]
  PIN la_oenb_mprj[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 -2.000 576.290 4.000 ;
    END
  END la_oenb_mprj[80]
  PIN la_oenb_mprj[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 -2.000 583.650 4.000 ;
    END
  END la_oenb_mprj[81]
  PIN la_oenb_mprj[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 -2.000 590.550 4.000 ;
    END
  END la_oenb_mprj[82]
  PIN la_oenb_mprj[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 -2.000 597.910 4.000 ;
    END
  END la_oenb_mprj[83]
  PIN la_oenb_mprj[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 -2.000 604.810 4.000 ;
    END
  END la_oenb_mprj[84]
  PIN la_oenb_mprj[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 -2.000 612.170 4.000 ;
    END
  END la_oenb_mprj[85]
  PIN la_oenb_mprj[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 -2.000 619.070 4.000 ;
    END
  END la_oenb_mprj[86]
  PIN la_oenb_mprj[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 -2.000 626.430 4.000 ;
    END
  END la_oenb_mprj[87]
  PIN la_oenb_mprj[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 -2.000 633.330 4.000 ;
    END
  END la_oenb_mprj[88]
  PIN la_oenb_mprj[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 -2.000 640.690 4.000 ;
    END
  END la_oenb_mprj[89]
  PIN la_oenb_mprj[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 -2.000 62.930 4.000 ;
    END
  END la_oenb_mprj[8]
  PIN la_oenb_mprj[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 -2.000 647.590 4.000 ;
    END
  END la_oenb_mprj[90]
  PIN la_oenb_mprj[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 -2.000 654.950 4.000 ;
    END
  END la_oenb_mprj[91]
  PIN la_oenb_mprj[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 -2.000 661.850 4.000 ;
    END
  END la_oenb_mprj[92]
  PIN la_oenb_mprj[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 -2.000 669.210 4.000 ;
    END
  END la_oenb_mprj[93]
  PIN la_oenb_mprj[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 -2.000 676.110 4.000 ;
    END
  END la_oenb_mprj[94]
  PIN la_oenb_mprj[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 -2.000 683.470 4.000 ;
    END
  END la_oenb_mprj[95]
  PIN la_oenb_mprj[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 -2.000 690.370 4.000 ;
    END
  END la_oenb_mprj[96]
  PIN la_oenb_mprj[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 -2.000 697.730 4.000 ;
    END
  END la_oenb_mprj[97]
  PIN la_oenb_mprj[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 -2.000 704.630 4.000 ;
    END
  END la_oenb_mprj[98]
  PIN la_oenb_mprj[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 -2.000 711.990 4.000 ;
    END
  END la_oenb_mprj[99]
  PIN la_oenb_mprj[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 -2.000 70.290 4.000 ;
    END
  END la_oenb_mprj[9]
  PIN mprj_ack_i_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.190 -2.000 913.470 4.000 ;
    END
  END mprj_ack_i_core
  PIN mprj_ack_i_user
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 116.000 5.430 122.000 ;
    END
  END mprj_ack_i_user
  PIN mprj_adr_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 -2.000 920.370 4.000 ;
    END
  END mprj_adr_o_core[0]
  PIN mprj_adr_o_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.810 -2.000 981.090 4.000 ;
    END
  END mprj_adr_o_core[10]
  PIN mprj_adr_o_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.870 -2.000 986.150 4.000 ;
    END
  END mprj_adr_o_core[11]
  PIN mprj_adr_o_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 -2.000 991.670 4.000 ;
    END
  END mprj_adr_o_core[12]
  PIN mprj_adr_o_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 -2.000 997.190 4.000 ;
    END
  END mprj_adr_o_core[13]
  PIN mprj_adr_o_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.970 -2.000 1002.250 4.000 ;
    END
  END mprj_adr_o_core[14]
  PIN mprj_adr_o_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.490 -2.000 1007.770 4.000 ;
    END
  END mprj_adr_o_core[15]
  PIN mprj_adr_o_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 -2.000 1013.290 4.000 ;
    END
  END mprj_adr_o_core[16]
  PIN mprj_adr_o_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.070 -2.000 1018.350 4.000 ;
    END
  END mprj_adr_o_core[17]
  PIN mprj_adr_o_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.590 -2.000 1023.870 4.000 ;
    END
  END mprj_adr_o_core[18]
  PIN mprj_adr_o_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.650 -2.000 1028.930 4.000 ;
    END
  END mprj_adr_o_core[19]
  PIN mprj_adr_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 -2.000 927.730 4.000 ;
    END
  END mprj_adr_o_core[1]
  PIN mprj_adr_o_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 -2.000 1034.450 4.000 ;
    END
  END mprj_adr_o_core[20]
  PIN mprj_adr_o_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.690 -2.000 1039.970 4.000 ;
    END
  END mprj_adr_o_core[21]
  PIN mprj_adr_o_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 -2.000 1045.030 4.000 ;
    END
  END mprj_adr_o_core[22]
  PIN mprj_adr_o_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 -2.000 1050.550 4.000 ;
    END
  END mprj_adr_o_core[23]
  PIN mprj_adr_o_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.790 -2.000 1056.070 4.000 ;
    END
  END mprj_adr_o_core[24]
  PIN mprj_adr_o_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.850 -2.000 1061.130 4.000 ;
    END
  END mprj_adr_o_core[25]
  PIN mprj_adr_o_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 -2.000 1066.650 4.000 ;
    END
  END mprj_adr_o_core[26]
  PIN mprj_adr_o_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 -2.000 1071.710 4.000 ;
    END
  END mprj_adr_o_core[27]
  PIN mprj_adr_o_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 -2.000 1077.230 4.000 ;
    END
  END mprj_adr_o_core[28]
  PIN mprj_adr_o_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.470 -2.000 1082.750 4.000 ;
    END
  END mprj_adr_o_core[29]
  PIN mprj_adr_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 -2.000 934.630 4.000 ;
    END
  END mprj_adr_o_core[2]
  PIN mprj_adr_o_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 -2.000 1087.810 4.000 ;
    END
  END mprj_adr_o_core[30]
  PIN mprj_adr_o_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.050 -2.000 1093.330 4.000 ;
    END
  END mprj_adr_o_core[31]
  PIN mprj_adr_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.710 -2.000 941.990 4.000 ;
    END
  END mprj_adr_o_core[3]
  PIN mprj_adr_o_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 -2.000 948.890 4.000 ;
    END
  END mprj_adr_o_core[4]
  PIN mprj_adr_o_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 -2.000 954.410 4.000 ;
    END
  END mprj_adr_o_core[5]
  PIN mprj_adr_o_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 -2.000 959.470 4.000 ;
    END
  END mprj_adr_o_core[6]
  PIN mprj_adr_o_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 -2.000 964.990 4.000 ;
    END
  END mprj_adr_o_core[7]
  PIN mprj_adr_o_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 -2.000 970.510 4.000 ;
    END
  END mprj_adr_o_core[8]
  PIN mprj_adr_o_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 -2.000 975.570 4.000 ;
    END
  END mprj_adr_o_core[9]
  PIN mprj_adr_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 116.000 14.630 122.000 ;
    END
  END mprj_adr_o_user[0]
  PIN mprj_adr_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 116.000 90.070 122.000 ;
    END
  END mprj_adr_o_user[10]
  PIN mprj_adr_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 116.000 96.970 122.000 ;
    END
  END mprj_adr_o_user[11]
  PIN mprj_adr_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 116.000 103.410 122.000 ;
    END
  END mprj_adr_o_user[12]
  PIN mprj_adr_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 116.000 110.310 122.000 ;
    END
  END mprj_adr_o_user[13]
  PIN mprj_adr_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 116.000 116.750 122.000 ;
    END
  END mprj_adr_o_user[14]
  PIN mprj_adr_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 116.000 123.650 122.000 ;
    END
  END mprj_adr_o_user[15]
  PIN mprj_adr_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 116.000 130.090 122.000 ;
    END
  END mprj_adr_o_user[16]
  PIN mprj_adr_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 116.000 136.990 122.000 ;
    END
  END mprj_adr_o_user[17]
  PIN mprj_adr_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 116.000 143.430 122.000 ;
    END
  END mprj_adr_o_user[18]
  PIN mprj_adr_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 116.000 150.330 122.000 ;
    END
  END mprj_adr_o_user[19]
  PIN mprj_adr_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 116.000 23.370 122.000 ;
    END
  END mprj_adr_o_user[1]
  PIN mprj_adr_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 116.000 156.770 122.000 ;
    END
  END mprj_adr_o_user[20]
  PIN mprj_adr_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 116.000 163.670 122.000 ;
    END
  END mprj_adr_o_user[21]
  PIN mprj_adr_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 116.000 170.110 122.000 ;
    END
  END mprj_adr_o_user[22]
  PIN mprj_adr_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 116.000 177.010 122.000 ;
    END
  END mprj_adr_o_user[23]
  PIN mprj_adr_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 116.000 183.450 122.000 ;
    END
  END mprj_adr_o_user[24]
  PIN mprj_adr_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 116.000 190.350 122.000 ;
    END
  END mprj_adr_o_user[25]
  PIN mprj_adr_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 116.000 196.790 122.000 ;
    END
  END mprj_adr_o_user[26]
  PIN mprj_adr_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 116.000 203.690 122.000 ;
    END
  END mprj_adr_o_user[27]
  PIN mprj_adr_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 116.000 210.130 122.000 ;
    END
  END mprj_adr_o_user[28]
  PIN mprj_adr_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 116.000 217.030 122.000 ;
    END
  END mprj_adr_o_user[29]
  PIN mprj_adr_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 116.000 32.110 122.000 ;
    END
  END mprj_adr_o_user[2]
  PIN mprj_adr_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 116.000 223.930 122.000 ;
    END
  END mprj_adr_o_user[30]
  PIN mprj_adr_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 116.000 230.370 122.000 ;
    END
  END mprj_adr_o_user[31]
  PIN mprj_adr_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 116.000 41.310 122.000 ;
    END
  END mprj_adr_o_user[3]
  PIN mprj_adr_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 116.000 50.050 122.000 ;
    END
  END mprj_adr_o_user[4]
  PIN mprj_adr_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 116.000 56.950 122.000 ;
    END
  END mprj_adr_o_user[5]
  PIN mprj_adr_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 116.000 63.390 122.000 ;
    END
  END mprj_adr_o_user[6]
  PIN mprj_adr_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 116.000 70.290 122.000 ;
    END
  END mprj_adr_o_user[7]
  PIN mprj_adr_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 116.000 76.730 122.000 ;
    END
  END mprj_adr_o_user[8]
  PIN mprj_adr_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 116.000 83.630 122.000 ;
    END
  END mprj_adr_o_user[9]
  PIN mprj_cyc_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 -2.000 914.850 4.000 ;
    END
  END mprj_cyc_o_core
  PIN mprj_cyc_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 116.000 7.730 122.000 ;
    END
  END mprj_cyc_o_user
  PIN mprj_dat_i_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 -2.000 922.210 4.000 ;
    END
  END mprj_dat_i_core[0]
  PIN mprj_dat_i_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 -2.000 982.930 4.000 ;
    END
  END mprj_dat_i_core[10]
  PIN mprj_dat_i_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.710 -2.000 987.990 4.000 ;
    END
  END mprj_dat_i_core[11]
  PIN mprj_dat_i_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230 -2.000 993.510 4.000 ;
    END
  END mprj_dat_i_core[12]
  PIN mprj_dat_i_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 -2.000 999.030 4.000 ;
    END
  END mprj_dat_i_core[13]
  PIN mprj_dat_i_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.810 -2.000 1004.090 4.000 ;
    END
  END mprj_dat_i_core[14]
  PIN mprj_dat_i_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.330 -2.000 1009.610 4.000 ;
    END
  END mprj_dat_i_core[15]
  PIN mprj_dat_i_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 -2.000 1014.670 4.000 ;
    END
  END mprj_dat_i_core[16]
  PIN mprj_dat_i_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.910 -2.000 1020.190 4.000 ;
    END
  END mprj_dat_i_core[17]
  PIN mprj_dat_i_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.430 -2.000 1025.710 4.000 ;
    END
  END mprj_dat_i_core[18]
  PIN mprj_dat_i_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 -2.000 1030.770 4.000 ;
    END
  END mprj_dat_i_core[19]
  PIN mprj_dat_i_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 -2.000 929.110 4.000 ;
    END
  END mprj_dat_i_core[1]
  PIN mprj_dat_i_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 -2.000 1036.290 4.000 ;
    END
  END mprj_dat_i_core[20]
  PIN mprj_dat_i_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.530 -2.000 1041.810 4.000 ;
    END
  END mprj_dat_i_core[21]
  PIN mprj_dat_i_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 -2.000 1046.870 4.000 ;
    END
  END mprj_dat_i_core[22]
  PIN mprj_dat_i_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.110 -2.000 1052.390 4.000 ;
    END
  END mprj_dat_i_core[23]
  PIN mprj_dat_i_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.170 -2.000 1057.450 4.000 ;
    END
  END mprj_dat_i_core[24]
  PIN mprj_dat_i_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 -2.000 1062.970 4.000 ;
    END
  END mprj_dat_i_core[25]
  PIN mprj_dat_i_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.210 -2.000 1068.490 4.000 ;
    END
  END mprj_dat_i_core[26]
  PIN mprj_dat_i_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.270 -2.000 1073.550 4.000 ;
    END
  END mprj_dat_i_core[27]
  PIN mprj_dat_i_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 -2.000 1079.070 4.000 ;
    END
  END mprj_dat_i_core[28]
  PIN mprj_dat_i_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 -2.000 1084.590 4.000 ;
    END
  END mprj_dat_i_core[29]
  PIN mprj_dat_i_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.190 -2.000 936.470 4.000 ;
    END
  END mprj_dat_i_core[2]
  PIN mprj_dat_i_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 -2.000 1089.650 4.000 ;
    END
  END mprj_dat_i_core[30]
  PIN mprj_dat_i_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 -2.000 1095.170 4.000 ;
    END
  END mprj_dat_i_core[31]
  PIN mprj_dat_i_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.090 -2.000 943.370 4.000 ;
    END
  END mprj_dat_i_core[3]
  PIN mprj_dat_i_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.450 -2.000 950.730 4.000 ;
    END
  END mprj_dat_i_core[4]
  PIN mprj_dat_i_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.970 -2.000 956.250 4.000 ;
    END
  END mprj_dat_i_core[5]
  PIN mprj_dat_i_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 -2.000 961.310 4.000 ;
    END
  END mprj_dat_i_core[6]
  PIN mprj_dat_i_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 -2.000 966.830 4.000 ;
    END
  END mprj_dat_i_core[7]
  PIN mprj_dat_i_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.610 -2.000 971.890 4.000 ;
    END
  END mprj_dat_i_core[8]
  PIN mprj_dat_i_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 -2.000 977.410 4.000 ;
    END
  END mprj_dat_i_core[9]
  PIN mprj_dat_i_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 116.000 16.470 122.000 ;
    END
  END mprj_dat_i_user[0]
  PIN mprj_dat_i_user[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 116.000 92.370 122.000 ;
    END
  END mprj_dat_i_user[10]
  PIN mprj_dat_i_user[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 116.000 98.810 122.000 ;
    END
  END mprj_dat_i_user[11]
  PIN mprj_dat_i_user[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 116.000 105.710 122.000 ;
    END
  END mprj_dat_i_user[12]
  PIN mprj_dat_i_user[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 116.000 112.610 122.000 ;
    END
  END mprj_dat_i_user[13]
  PIN mprj_dat_i_user[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 116.000 119.050 122.000 ;
    END
  END mprj_dat_i_user[14]
  PIN mprj_dat_i_user[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 116.000 125.950 122.000 ;
    END
  END mprj_dat_i_user[15]
  PIN mprj_dat_i_user[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 116.000 132.390 122.000 ;
    END
  END mprj_dat_i_user[16]
  PIN mprj_dat_i_user[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 116.000 139.290 122.000 ;
    END
  END mprj_dat_i_user[17]
  PIN mprj_dat_i_user[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 116.000 145.730 122.000 ;
    END
  END mprj_dat_i_user[18]
  PIN mprj_dat_i_user[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 116.000 152.630 122.000 ;
    END
  END mprj_dat_i_user[19]
  PIN mprj_dat_i_user[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 116.000 25.670 122.000 ;
    END
  END mprj_dat_i_user[1]
  PIN mprj_dat_i_user[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 116.000 159.070 122.000 ;
    END
  END mprj_dat_i_user[20]
  PIN mprj_dat_i_user[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 116.000 165.970 122.000 ;
    END
  END mprj_dat_i_user[21]
  PIN mprj_dat_i_user[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 116.000 172.410 122.000 ;
    END
  END mprj_dat_i_user[22]
  PIN mprj_dat_i_user[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 116.000 179.310 122.000 ;
    END
  END mprj_dat_i_user[23]
  PIN mprj_dat_i_user[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 116.000 185.750 122.000 ;
    END
  END mprj_dat_i_user[24]
  PIN mprj_dat_i_user[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 116.000 192.650 122.000 ;
    END
  END mprj_dat_i_user[25]
  PIN mprj_dat_i_user[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 116.000 199.090 122.000 ;
    END
  END mprj_dat_i_user[26]
  PIN mprj_dat_i_user[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 116.000 205.990 122.000 ;
    END
  END mprj_dat_i_user[27]
  PIN mprj_dat_i_user[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 116.000 212.430 122.000 ;
    END
  END mprj_dat_i_user[28]
  PIN mprj_dat_i_user[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 116.000 219.330 122.000 ;
    END
  END mprj_dat_i_user[29]
  PIN mprj_dat_i_user[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 116.000 34.410 122.000 ;
    END
  END mprj_dat_i_user[2]
  PIN mprj_dat_i_user[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 116.000 225.770 122.000 ;
    END
  END mprj_dat_i_user[30]
  PIN mprj_dat_i_user[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 116.000 232.670 122.000 ;
    END
  END mprj_dat_i_user[31]
  PIN mprj_dat_i_user[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 116.000 43.150 122.000 ;
    END
  END mprj_dat_i_user[3]
  PIN mprj_dat_i_user[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 116.000 52.350 122.000 ;
    END
  END mprj_dat_i_user[4]
  PIN mprj_dat_i_user[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 116.000 58.790 122.000 ;
    END
  END mprj_dat_i_user[5]
  PIN mprj_dat_i_user[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 116.000 65.690 122.000 ;
    END
  END mprj_dat_i_user[6]
  PIN mprj_dat_i_user[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 116.000 72.130 122.000 ;
    END
  END mprj_dat_i_user[7]
  PIN mprj_dat_i_user[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 116.000 79.030 122.000 ;
    END
  END mprj_dat_i_user[8]
  PIN mprj_dat_i_user[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 116.000 85.470 122.000 ;
    END
  END mprj_dat_i_user[9]
  PIN mprj_dat_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.770 -2.000 924.050 4.000 ;
    END
  END mprj_dat_o_core[0]
  PIN mprj_dat_o_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.490 -2.000 984.770 4.000 ;
    END
  END mprj_dat_o_core[10]
  PIN mprj_dat_o_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 -2.000 989.830 4.000 ;
    END
  END mprj_dat_o_core[11]
  PIN mprj_dat_o_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 -2.000 995.350 4.000 ;
    END
  END mprj_dat_o_core[12]
  PIN mprj_dat_o_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.130 -2.000 1000.410 4.000 ;
    END
  END mprj_dat_o_core[13]
  PIN mprj_dat_o_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.650 -2.000 1005.930 4.000 ;
    END
  END mprj_dat_o_core[14]
  PIN mprj_dat_o_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 -2.000 1011.450 4.000 ;
    END
  END mprj_dat_o_core[15]
  PIN mprj_dat_o_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.230 -2.000 1016.510 4.000 ;
    END
  END mprj_dat_o_core[16]
  PIN mprj_dat_o_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.750 -2.000 1022.030 4.000 ;
    END
  END mprj_dat_o_core[17]
  PIN mprj_dat_o_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 -2.000 1027.550 4.000 ;
    END
  END mprj_dat_o_core[18]
  PIN mprj_dat_o_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.330 -2.000 1032.610 4.000 ;
    END
  END mprj_dat_o_core[19]
  PIN mprj_dat_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 -2.000 930.950 4.000 ;
    END
  END mprj_dat_o_core[1]
  PIN mprj_dat_o_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 -2.000 1038.130 4.000 ;
    END
  END mprj_dat_o_core[20]
  PIN mprj_dat_o_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.910 -2.000 1043.190 4.000 ;
    END
  END mprj_dat_o_core[21]
  PIN mprj_dat_o_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.430 -2.000 1048.710 4.000 ;
    END
  END mprj_dat_o_core[22]
  PIN mprj_dat_o_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.950 -2.000 1054.230 4.000 ;
    END
  END mprj_dat_o_core[23]
  PIN mprj_dat_o_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 -2.000 1059.290 4.000 ;
    END
  END mprj_dat_o_core[24]
  PIN mprj_dat_o_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.530 -2.000 1064.810 4.000 ;
    END
  END mprj_dat_o_core[25]
  PIN mprj_dat_o_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.050 -2.000 1070.330 4.000 ;
    END
  END mprj_dat_o_core[26]
  PIN mprj_dat_o_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.110 -2.000 1075.390 4.000 ;
    END
  END mprj_dat_o_core[27]
  PIN mprj_dat_o_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630 -2.000 1080.910 4.000 ;
    END
  END mprj_dat_o_core[28]
  PIN mprj_dat_o_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.690 -2.000 1085.970 4.000 ;
    END
  END mprj_dat_o_core[29]
  PIN mprj_dat_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 -2.000 938.310 4.000 ;
    END
  END mprj_dat_o_core[2]
  PIN mprj_dat_o_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 -2.000 1091.490 4.000 ;
    END
  END mprj_dat_o_core[30]
  PIN mprj_dat_o_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.730 -2.000 1097.010 4.000 ;
    END
  END mprj_dat_o_core[31]
  PIN mprj_dat_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 -2.000 945.210 4.000 ;
    END
  END mprj_dat_o_core[3]
  PIN mprj_dat_o_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 -2.000 952.570 4.000 ;
    END
  END mprj_dat_o_core[4]
  PIN mprj_dat_o_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 -2.000 957.630 4.000 ;
    END
  END mprj_dat_o_core[5]
  PIN mprj_dat_o_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 -2.000 963.150 4.000 ;
    END
  END mprj_dat_o_core[6]
  PIN mprj_dat_o_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 -2.000 968.670 4.000 ;
    END
  END mprj_dat_o_core[7]
  PIN mprj_dat_o_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.450 -2.000 973.730 4.000 ;
    END
  END mprj_dat_o_core[8]
  PIN mprj_dat_o_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 -2.000 979.250 4.000 ;
    END
  END mprj_dat_o_core[9]
  PIN mprj_dat_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 116.000 18.770 122.000 ;
    END
  END mprj_dat_o_user[0]
  PIN mprj_dat_o_user[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 116.000 94.670 122.000 ;
    END
  END mprj_dat_o_user[10]
  PIN mprj_dat_o_user[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 116.000 101.110 122.000 ;
    END
  END mprj_dat_o_user[11]
  PIN mprj_dat_o_user[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 116.000 108.010 122.000 ;
    END
  END mprj_dat_o_user[12]
  PIN mprj_dat_o_user[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 116.000 114.450 122.000 ;
    END
  END mprj_dat_o_user[13]
  PIN mprj_dat_o_user[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 116.000 121.350 122.000 ;
    END
  END mprj_dat_o_user[14]
  PIN mprj_dat_o_user[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 116.000 127.790 122.000 ;
    END
  END mprj_dat_o_user[15]
  PIN mprj_dat_o_user[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 116.000 134.690 122.000 ;
    END
  END mprj_dat_o_user[16]
  PIN mprj_dat_o_user[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 116.000 141.130 122.000 ;
    END
  END mprj_dat_o_user[17]
  PIN mprj_dat_o_user[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 116.000 148.030 122.000 ;
    END
  END mprj_dat_o_user[18]
  PIN mprj_dat_o_user[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 116.000 154.470 122.000 ;
    END
  END mprj_dat_o_user[19]
  PIN mprj_dat_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 116.000 27.970 122.000 ;
    END
  END mprj_dat_o_user[1]
  PIN mprj_dat_o_user[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 116.000 161.370 122.000 ;
    END
  END mprj_dat_o_user[20]
  PIN mprj_dat_o_user[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 116.000 168.270 122.000 ;
    END
  END mprj_dat_o_user[21]
  PIN mprj_dat_o_user[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 116.000 174.710 122.000 ;
    END
  END mprj_dat_o_user[22]
  PIN mprj_dat_o_user[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 116.000 181.610 122.000 ;
    END
  END mprj_dat_o_user[23]
  PIN mprj_dat_o_user[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 116.000 188.050 122.000 ;
    END
  END mprj_dat_o_user[24]
  PIN mprj_dat_o_user[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 116.000 194.950 122.000 ;
    END
  END mprj_dat_o_user[25]
  PIN mprj_dat_o_user[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 116.000 201.390 122.000 ;
    END
  END mprj_dat_o_user[26]
  PIN mprj_dat_o_user[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 116.000 208.290 122.000 ;
    END
  END mprj_dat_o_user[27]
  PIN mprj_dat_o_user[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 116.000 214.730 122.000 ;
    END
  END mprj_dat_o_user[28]
  PIN mprj_dat_o_user[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 116.000 221.630 122.000 ;
    END
  END mprj_dat_o_user[29]
  PIN mprj_dat_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 116.000 36.710 122.000 ;
    END
  END mprj_dat_o_user[2]
  PIN mprj_dat_o_user[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 116.000 228.070 122.000 ;
    END
  END mprj_dat_o_user[30]
  PIN mprj_dat_o_user[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 116.000 234.970 122.000 ;
    END
  END mprj_dat_o_user[31]
  PIN mprj_dat_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 116.000 45.450 122.000 ;
    END
  END mprj_dat_o_user[3]
  PIN mprj_dat_o_user[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 116.000 54.650 122.000 ;
    END
  END mprj_dat_o_user[4]
  PIN mprj_dat_o_user[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 116.000 61.090 122.000 ;
    END
  END mprj_dat_o_user[5]
  PIN mprj_dat_o_user[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 116.000 67.990 122.000 ;
    END
  END mprj_dat_o_user[6]
  PIN mprj_dat_o_user[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 116.000 74.430 122.000 ;
    END
  END mprj_dat_o_user[7]
  PIN mprj_dat_o_user[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 116.000 81.330 122.000 ;
    END
  END mprj_dat_o_user[8]
  PIN mprj_dat_o_user[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 116.000 87.770 122.000 ;
    END
  END mprj_dat_o_user[9]
  PIN mprj_iena_wb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 -2.000 1098.850 4.000 ;
    END
  END mprj_iena_wb
  PIN mprj_sel_o_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 -2.000 925.890 4.000 ;
    END
  END mprj_sel_o_core[0]
  PIN mprj_sel_o_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 -2.000 932.790 4.000 ;
    END
  END mprj_sel_o_core[1]
  PIN mprj_sel_o_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 -2.000 940.150 4.000 ;
    END
  END mprj_sel_o_core[2]
  PIN mprj_sel_o_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 -2.000 947.050 4.000 ;
    END
  END mprj_sel_o_core[3]
  PIN mprj_sel_o_user[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 116.000 21.070 122.000 ;
    END
  END mprj_sel_o_user[0]
  PIN mprj_sel_o_user[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 116.000 29.810 122.000 ;
    END
  END mprj_sel_o_user[1]
  PIN mprj_sel_o_user[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 116.000 39.010 122.000 ;
    END
  END mprj_sel_o_user[2]
  PIN mprj_sel_o_user[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 116.000 47.750 122.000 ;
    END
  END mprj_sel_o_user[3]
  PIN mprj_stb_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 -2.000 916.690 4.000 ;
    END
  END mprj_stb_o_core
  PIN mprj_stb_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 116.000 10.030 122.000 ;
    END
  END mprj_stb_o_user
  PIN mprj_we_o_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 -2.000 918.530 4.000 ;
    END
  END mprj_we_o_core
  PIN mprj_we_o_user
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 116.000 12.330 122.000 ;
    END
  END mprj_we_o_user
  PIN user1_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 5.480 1102.000 6.080 ;
    END
  END user1_vcc_powergood
  PIN user1_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 17.040 1102.000 17.640 ;
    END
  END user1_vdd_powergood
  PIN user2_vcc_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 29.280 1102.000 29.880 ;
    END
  END user2_vcc_powergood
  PIN user2_vdd_powergood
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 40.840 1102.000 41.440 ;
    END
  END user2_vdd_powergood
  PIN user_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 116.000 1.290 122.000 ;
    END
  END user_clock
  PIN user_clock2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 116.000 1091.950 122.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 53.080 1102.000 53.680 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 65.320 1102.000 65.920 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 76.880 1102.000 77.480 ;
    END
  END user_irq[2]
  PIN user_irq_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.970 116.000 1094.250 122.000 ;
    END
  END user_irq_core[0]
  PIN user_irq_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.270 116.000 1096.550 122.000 ;
    END
  END user_irq_core[1]
  PIN user_irq_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 116.000 1098.850 122.000 ;
    END
  END user_irq_core[2]
  PIN user_irq_ena[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 89.120 1102.000 89.720 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 100.680 1102.000 101.280 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 112.920 1102.000 113.520 ;
    END
  END user_irq_ena[2]
  PIN user_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 116.000 3.130 122.000 ;
    END
  END user_reset
  PIN vccd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.070 5.200 20.970 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 170.570 5.200 171.470 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.070 5.200 321.970 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.570 5.200 472.470 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 622.070 5.200 622.970 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 772.570 5.200 773.470 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.070 5.200 923.970 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.570 5.200 1074.470 114.480 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.170 5.440 25.070 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.670 5.440 175.570 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.170 5.440 326.070 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.670 5.440 476.570 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 626.170 5.440 627.070 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 776.670 5.440 777.570 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.170 5.440 928.070 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1077.670 5.440 1078.570 114.240 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.270 5.440 29.170 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 178.770 5.440 179.670 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 329.270 5.440 330.170 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 479.770 5.440 480.670 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 630.270 5.440 631.170 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 780.770 5.440 781.670 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.270 5.440 932.170 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1081.770 5.440 1082.670 114.240 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 934.070 5.440 934.970 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1084.570 5.440 1085.470 114.240 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 937.070 5.440 937.970 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1087.570 5.440 1088.470 114.240 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1009.320 5.440 1010.220 114.240 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1012.320 5.440 1013.220 114.240 ;
    END
  END vssa2
  PIN vssd
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.320 5.200 96.220 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 245.820 5.200 246.720 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.320 5.200 397.220 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.820 5.200 547.720 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 697.320 5.200 698.220 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 847.820 5.200 848.720 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.320 5.200 999.220 114.480 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 99.420 5.440 100.320 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.920 5.440 250.820 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 400.420 5.440 401.320 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.920 5.440 551.820 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.420 5.440 702.320 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 851.920 5.440 852.820 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1002.420 5.440 1003.320 114.240 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 103.520 5.440 104.420 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.020 5.440 254.920 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.520 5.440 405.420 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 555.020 5.440 555.920 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 705.520 5.440 706.420 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.020 5.440 856.920 114.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1006.520 5.440 1007.420 114.240 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 5.520 0.085 1094.340 119.935 ;
      LAYER met1 ;
        RECT 0.530 0.040 1098.870 119.965 ;
      LAYER met2 ;
        RECT 0.560 115.720 0.730 119.670 ;
        RECT 1.570 115.720 2.570 119.670 ;
        RECT 3.410 115.720 4.870 119.670 ;
        RECT 5.710 115.720 7.170 119.670 ;
        RECT 8.010 115.720 9.470 119.670 ;
        RECT 10.310 115.720 11.770 119.670 ;
        RECT 12.610 115.720 14.070 119.670 ;
        RECT 14.910 115.720 15.910 119.670 ;
        RECT 16.750 115.720 18.210 119.670 ;
        RECT 19.050 115.720 20.510 119.670 ;
        RECT 21.350 115.720 22.810 119.670 ;
        RECT 23.650 115.720 25.110 119.670 ;
        RECT 25.950 115.720 27.410 119.670 ;
        RECT 28.250 115.720 29.250 119.670 ;
        RECT 30.090 115.720 31.550 119.670 ;
        RECT 32.390 115.720 33.850 119.670 ;
        RECT 34.690 115.720 36.150 119.670 ;
        RECT 36.990 115.720 38.450 119.670 ;
        RECT 39.290 115.720 40.750 119.670 ;
        RECT 41.590 115.720 42.590 119.670 ;
        RECT 43.430 115.720 44.890 119.670 ;
        RECT 45.730 115.720 47.190 119.670 ;
        RECT 48.030 115.720 49.490 119.670 ;
        RECT 50.330 115.720 51.790 119.670 ;
        RECT 52.630 115.720 54.090 119.670 ;
        RECT 54.930 115.720 56.390 119.670 ;
        RECT 57.230 115.720 58.230 119.670 ;
        RECT 59.070 115.720 60.530 119.670 ;
        RECT 61.370 115.720 62.830 119.670 ;
        RECT 63.670 115.720 65.130 119.670 ;
        RECT 65.970 115.720 67.430 119.670 ;
        RECT 68.270 115.720 69.730 119.670 ;
        RECT 70.570 115.720 71.570 119.670 ;
        RECT 72.410 115.720 73.870 119.670 ;
        RECT 74.710 115.720 76.170 119.670 ;
        RECT 77.010 115.720 78.470 119.670 ;
        RECT 79.310 115.720 80.770 119.670 ;
        RECT 81.610 115.720 83.070 119.670 ;
        RECT 83.910 115.720 84.910 119.670 ;
        RECT 85.750 115.720 87.210 119.670 ;
        RECT 88.050 115.720 89.510 119.670 ;
        RECT 90.350 115.720 91.810 119.670 ;
        RECT 92.650 115.720 94.110 119.670 ;
        RECT 94.950 115.720 96.410 119.670 ;
        RECT 97.250 115.720 98.250 119.670 ;
        RECT 99.090 115.720 100.550 119.670 ;
        RECT 101.390 115.720 102.850 119.670 ;
        RECT 103.690 115.720 105.150 119.670 ;
        RECT 105.990 115.720 107.450 119.670 ;
        RECT 108.290 115.720 109.750 119.670 ;
        RECT 110.590 115.720 112.050 119.670 ;
        RECT 112.890 115.720 113.890 119.670 ;
        RECT 114.730 115.720 116.190 119.670 ;
        RECT 117.030 115.720 118.490 119.670 ;
        RECT 119.330 115.720 120.790 119.670 ;
        RECT 121.630 115.720 123.090 119.670 ;
        RECT 123.930 115.720 125.390 119.670 ;
        RECT 126.230 115.720 127.230 119.670 ;
        RECT 128.070 115.720 129.530 119.670 ;
        RECT 130.370 115.720 131.830 119.670 ;
        RECT 132.670 115.720 134.130 119.670 ;
        RECT 134.970 115.720 136.430 119.670 ;
        RECT 137.270 115.720 138.730 119.670 ;
        RECT 139.570 115.720 140.570 119.670 ;
        RECT 141.410 115.720 142.870 119.670 ;
        RECT 143.710 115.720 145.170 119.670 ;
        RECT 146.010 115.720 147.470 119.670 ;
        RECT 148.310 115.720 149.770 119.670 ;
        RECT 150.610 115.720 152.070 119.670 ;
        RECT 152.910 115.720 153.910 119.670 ;
        RECT 154.750 115.720 156.210 119.670 ;
        RECT 157.050 115.720 158.510 119.670 ;
        RECT 159.350 115.720 160.810 119.670 ;
        RECT 161.650 115.720 163.110 119.670 ;
        RECT 163.950 115.720 165.410 119.670 ;
        RECT 166.250 115.720 167.710 119.670 ;
        RECT 168.550 115.720 169.550 119.670 ;
        RECT 170.390 115.720 171.850 119.670 ;
        RECT 172.690 115.720 174.150 119.670 ;
        RECT 174.990 115.720 176.450 119.670 ;
        RECT 177.290 115.720 178.750 119.670 ;
        RECT 179.590 115.720 181.050 119.670 ;
        RECT 181.890 115.720 182.890 119.670 ;
        RECT 183.730 115.720 185.190 119.670 ;
        RECT 186.030 115.720 187.490 119.670 ;
        RECT 188.330 115.720 189.790 119.670 ;
        RECT 190.630 115.720 192.090 119.670 ;
        RECT 192.930 115.720 194.390 119.670 ;
        RECT 195.230 115.720 196.230 119.670 ;
        RECT 197.070 115.720 198.530 119.670 ;
        RECT 199.370 115.720 200.830 119.670 ;
        RECT 201.670 115.720 203.130 119.670 ;
        RECT 203.970 115.720 205.430 119.670 ;
        RECT 206.270 115.720 207.730 119.670 ;
        RECT 208.570 115.720 209.570 119.670 ;
        RECT 210.410 115.720 211.870 119.670 ;
        RECT 212.710 115.720 214.170 119.670 ;
        RECT 215.010 115.720 216.470 119.670 ;
        RECT 217.310 115.720 218.770 119.670 ;
        RECT 219.610 115.720 221.070 119.670 ;
        RECT 221.910 115.720 223.370 119.670 ;
        RECT 224.210 115.720 225.210 119.670 ;
        RECT 226.050 115.720 227.510 119.670 ;
        RECT 228.350 115.720 229.810 119.670 ;
        RECT 230.650 115.720 232.110 119.670 ;
        RECT 232.950 115.720 234.410 119.670 ;
        RECT 235.250 115.720 236.710 119.670 ;
        RECT 237.550 115.720 238.550 119.670 ;
        RECT 239.390 115.720 240.850 119.670 ;
        RECT 241.690 115.720 243.150 119.670 ;
        RECT 243.990 115.720 245.450 119.670 ;
        RECT 246.290 115.720 247.750 119.670 ;
        RECT 248.590 115.720 250.050 119.670 ;
        RECT 250.890 115.720 251.890 119.670 ;
        RECT 252.730 115.720 254.190 119.670 ;
        RECT 255.030 115.720 256.490 119.670 ;
        RECT 257.330 115.720 258.790 119.670 ;
        RECT 259.630 115.720 261.090 119.670 ;
        RECT 261.930 115.720 263.390 119.670 ;
        RECT 264.230 115.720 265.230 119.670 ;
        RECT 266.070 115.720 267.530 119.670 ;
        RECT 268.370 115.720 269.830 119.670 ;
        RECT 270.670 115.720 272.130 119.670 ;
        RECT 272.970 115.720 274.430 119.670 ;
        RECT 275.270 115.720 276.730 119.670 ;
        RECT 277.570 115.720 279.030 119.670 ;
        RECT 279.870 115.720 280.870 119.670 ;
        RECT 281.710 115.720 283.170 119.670 ;
        RECT 284.010 115.720 285.470 119.670 ;
        RECT 286.310 115.720 287.770 119.670 ;
        RECT 288.610 115.720 290.070 119.670 ;
        RECT 290.910 115.720 292.370 119.670 ;
        RECT 293.210 115.720 294.210 119.670 ;
        RECT 295.050 115.720 296.510 119.670 ;
        RECT 297.350 115.720 298.810 119.670 ;
        RECT 299.650 115.720 301.110 119.670 ;
        RECT 301.950 115.720 303.410 119.670 ;
        RECT 304.250 115.720 305.710 119.670 ;
        RECT 306.550 115.720 307.550 119.670 ;
        RECT 308.390 115.720 309.850 119.670 ;
        RECT 310.690 115.720 312.150 119.670 ;
        RECT 312.990 115.720 314.450 119.670 ;
        RECT 315.290 115.720 316.750 119.670 ;
        RECT 317.590 115.720 319.050 119.670 ;
        RECT 319.890 115.720 320.890 119.670 ;
        RECT 321.730 115.720 323.190 119.670 ;
        RECT 324.030 115.720 325.490 119.670 ;
        RECT 326.330 115.720 327.790 119.670 ;
        RECT 328.630 115.720 330.090 119.670 ;
        RECT 330.930 115.720 332.390 119.670 ;
        RECT 333.230 115.720 334.690 119.670 ;
        RECT 335.530 115.720 336.530 119.670 ;
        RECT 337.370 115.720 338.830 119.670 ;
        RECT 339.670 115.720 341.130 119.670 ;
        RECT 341.970 115.720 343.430 119.670 ;
        RECT 344.270 115.720 345.730 119.670 ;
        RECT 346.570 115.720 348.030 119.670 ;
        RECT 348.870 115.720 349.870 119.670 ;
        RECT 350.710 115.720 352.170 119.670 ;
        RECT 353.010 115.720 354.470 119.670 ;
        RECT 355.310 115.720 356.770 119.670 ;
        RECT 357.610 115.720 359.070 119.670 ;
        RECT 359.910 115.720 361.370 119.670 ;
        RECT 362.210 115.720 363.210 119.670 ;
        RECT 364.050 115.720 365.510 119.670 ;
        RECT 366.350 115.720 367.810 119.670 ;
        RECT 368.650 115.720 370.110 119.670 ;
        RECT 370.950 115.720 372.410 119.670 ;
        RECT 373.250 115.720 374.710 119.670 ;
        RECT 375.550 115.720 376.550 119.670 ;
        RECT 377.390 115.720 378.850 119.670 ;
        RECT 379.690 115.720 381.150 119.670 ;
        RECT 381.990 115.720 383.450 119.670 ;
        RECT 384.290 115.720 385.750 119.670 ;
        RECT 386.590 115.720 388.050 119.670 ;
        RECT 388.890 115.720 390.350 119.670 ;
        RECT 391.190 115.720 392.190 119.670 ;
        RECT 393.030 115.720 394.490 119.670 ;
        RECT 395.330 115.720 396.790 119.670 ;
        RECT 397.630 115.720 399.090 119.670 ;
        RECT 399.930 115.720 401.390 119.670 ;
        RECT 402.230 115.720 403.690 119.670 ;
        RECT 404.530 115.720 405.530 119.670 ;
        RECT 406.370 115.720 407.830 119.670 ;
        RECT 408.670 115.720 410.130 119.670 ;
        RECT 410.970 115.720 412.430 119.670 ;
        RECT 413.270 115.720 414.730 119.670 ;
        RECT 415.570 115.720 417.030 119.670 ;
        RECT 417.870 115.720 418.870 119.670 ;
        RECT 419.710 115.720 421.170 119.670 ;
        RECT 422.010 115.720 423.470 119.670 ;
        RECT 424.310 115.720 425.770 119.670 ;
        RECT 426.610 115.720 428.070 119.670 ;
        RECT 428.910 115.720 430.370 119.670 ;
        RECT 431.210 115.720 432.210 119.670 ;
        RECT 433.050 115.720 434.510 119.670 ;
        RECT 435.350 115.720 436.810 119.670 ;
        RECT 437.650 115.720 439.110 119.670 ;
        RECT 439.950 115.720 441.410 119.670 ;
        RECT 442.250 115.720 443.710 119.670 ;
        RECT 444.550 115.720 446.010 119.670 ;
        RECT 446.850 115.720 447.850 119.670 ;
        RECT 448.690 115.720 450.150 119.670 ;
        RECT 450.990 115.720 452.450 119.670 ;
        RECT 453.290 115.720 454.750 119.670 ;
        RECT 455.590 115.720 457.050 119.670 ;
        RECT 457.890 115.720 459.350 119.670 ;
        RECT 460.190 115.720 461.190 119.670 ;
        RECT 462.030 115.720 463.490 119.670 ;
        RECT 464.330 115.720 465.790 119.670 ;
        RECT 466.630 115.720 468.090 119.670 ;
        RECT 468.930 115.720 470.390 119.670 ;
        RECT 471.230 115.720 472.690 119.670 ;
        RECT 473.530 115.720 474.530 119.670 ;
        RECT 475.370 115.720 476.830 119.670 ;
        RECT 477.670 115.720 479.130 119.670 ;
        RECT 479.970 115.720 481.430 119.670 ;
        RECT 482.270 115.720 483.730 119.670 ;
        RECT 484.570 115.720 486.030 119.670 ;
        RECT 486.870 115.720 487.870 119.670 ;
        RECT 488.710 115.720 490.170 119.670 ;
        RECT 491.010 115.720 492.470 119.670 ;
        RECT 493.310 115.720 494.770 119.670 ;
        RECT 495.610 115.720 497.070 119.670 ;
        RECT 497.910 115.720 499.370 119.670 ;
        RECT 500.210 115.720 501.670 119.670 ;
        RECT 502.510 115.720 503.510 119.670 ;
        RECT 504.350 115.720 505.810 119.670 ;
        RECT 506.650 115.720 508.110 119.670 ;
        RECT 508.950 115.720 510.410 119.670 ;
        RECT 511.250 115.720 512.710 119.670 ;
        RECT 513.550 115.720 515.010 119.670 ;
        RECT 515.850 115.720 516.850 119.670 ;
        RECT 517.690 115.720 519.150 119.670 ;
        RECT 519.990 115.720 521.450 119.670 ;
        RECT 522.290 115.720 523.750 119.670 ;
        RECT 524.590 115.720 526.050 119.670 ;
        RECT 526.890 115.720 528.350 119.670 ;
        RECT 529.190 115.720 530.190 119.670 ;
        RECT 531.030 115.720 532.490 119.670 ;
        RECT 533.330 115.720 534.790 119.670 ;
        RECT 535.630 115.720 537.090 119.670 ;
        RECT 537.930 115.720 539.390 119.670 ;
        RECT 540.230 115.720 541.690 119.670 ;
        RECT 542.530 115.720 543.530 119.670 ;
        RECT 544.370 115.720 545.830 119.670 ;
        RECT 546.670 115.720 548.130 119.670 ;
        RECT 548.970 115.720 550.430 119.670 ;
        RECT 551.270 115.720 552.730 119.670 ;
        RECT 553.570 115.720 555.030 119.670 ;
        RECT 555.870 115.720 557.330 119.670 ;
        RECT 558.170 115.720 559.170 119.670 ;
        RECT 560.010 115.720 561.470 119.670 ;
        RECT 562.310 115.720 563.770 119.670 ;
        RECT 564.610 115.720 566.070 119.670 ;
        RECT 566.910 115.720 568.370 119.670 ;
        RECT 569.210 115.720 570.670 119.670 ;
        RECT 571.510 115.720 572.510 119.670 ;
        RECT 573.350 115.720 574.810 119.670 ;
        RECT 575.650 115.720 577.110 119.670 ;
        RECT 577.950 115.720 579.410 119.670 ;
        RECT 580.250 115.720 581.710 119.670 ;
        RECT 582.550 115.720 584.010 119.670 ;
        RECT 584.850 115.720 585.850 119.670 ;
        RECT 586.690 115.720 588.150 119.670 ;
        RECT 588.990 115.720 590.450 119.670 ;
        RECT 591.290 115.720 592.750 119.670 ;
        RECT 593.590 115.720 595.050 119.670 ;
        RECT 595.890 115.720 597.350 119.670 ;
        RECT 598.190 115.720 599.190 119.670 ;
        RECT 600.030 115.720 601.490 119.670 ;
        RECT 602.330 115.720 603.790 119.670 ;
        RECT 604.630 115.720 606.090 119.670 ;
        RECT 606.930 115.720 608.390 119.670 ;
        RECT 609.230 115.720 610.690 119.670 ;
        RECT 611.530 115.720 612.990 119.670 ;
        RECT 613.830 115.720 614.830 119.670 ;
        RECT 615.670 115.720 617.130 119.670 ;
        RECT 617.970 115.720 619.430 119.670 ;
        RECT 620.270 115.720 621.730 119.670 ;
        RECT 622.570 115.720 624.030 119.670 ;
        RECT 624.870 115.720 626.330 119.670 ;
        RECT 627.170 115.720 628.170 119.670 ;
        RECT 629.010 115.720 630.470 119.670 ;
        RECT 631.310 115.720 632.770 119.670 ;
        RECT 633.610 115.720 635.070 119.670 ;
        RECT 635.910 115.720 637.370 119.670 ;
        RECT 638.210 115.720 639.670 119.670 ;
        RECT 640.510 115.720 641.510 119.670 ;
        RECT 642.350 115.720 643.810 119.670 ;
        RECT 644.650 115.720 646.110 119.670 ;
        RECT 646.950 115.720 648.410 119.670 ;
        RECT 649.250 115.720 650.710 119.670 ;
        RECT 651.550 115.720 653.010 119.670 ;
        RECT 653.850 115.720 654.850 119.670 ;
        RECT 655.690 115.720 657.150 119.670 ;
        RECT 657.990 115.720 659.450 119.670 ;
        RECT 660.290 115.720 661.750 119.670 ;
        RECT 662.590 115.720 664.050 119.670 ;
        RECT 664.890 115.720 666.350 119.670 ;
        RECT 667.190 115.720 668.650 119.670 ;
        RECT 669.490 115.720 670.490 119.670 ;
        RECT 671.330 115.720 672.790 119.670 ;
        RECT 673.630 115.720 675.090 119.670 ;
        RECT 675.930 115.720 677.390 119.670 ;
        RECT 678.230 115.720 679.690 119.670 ;
        RECT 680.530 115.720 681.990 119.670 ;
        RECT 682.830 115.720 683.830 119.670 ;
        RECT 684.670 115.720 686.130 119.670 ;
        RECT 686.970 115.720 688.430 119.670 ;
        RECT 689.270 115.720 690.730 119.670 ;
        RECT 691.570 115.720 693.030 119.670 ;
        RECT 693.870 115.720 695.330 119.670 ;
        RECT 696.170 115.720 697.170 119.670 ;
        RECT 698.010 115.720 699.470 119.670 ;
        RECT 700.310 115.720 701.770 119.670 ;
        RECT 702.610 115.720 704.070 119.670 ;
        RECT 704.910 115.720 706.370 119.670 ;
        RECT 707.210 115.720 708.670 119.670 ;
        RECT 709.510 115.720 710.510 119.670 ;
        RECT 711.350 115.720 712.810 119.670 ;
        RECT 713.650 115.720 715.110 119.670 ;
        RECT 715.950 115.720 717.410 119.670 ;
        RECT 718.250 115.720 719.710 119.670 ;
        RECT 720.550 115.720 722.010 119.670 ;
        RECT 722.850 115.720 724.310 119.670 ;
        RECT 725.150 115.720 726.150 119.670 ;
        RECT 726.990 115.720 728.450 119.670 ;
        RECT 729.290 115.720 730.750 119.670 ;
        RECT 731.590 115.720 733.050 119.670 ;
        RECT 733.890 115.720 735.350 119.670 ;
        RECT 736.190 115.720 737.650 119.670 ;
        RECT 738.490 115.720 739.490 119.670 ;
        RECT 740.330 115.720 741.790 119.670 ;
        RECT 742.630 115.720 744.090 119.670 ;
        RECT 744.930 115.720 746.390 119.670 ;
        RECT 747.230 115.720 748.690 119.670 ;
        RECT 749.530 115.720 750.990 119.670 ;
        RECT 751.830 115.720 752.830 119.670 ;
        RECT 753.670 115.720 755.130 119.670 ;
        RECT 755.970 115.720 757.430 119.670 ;
        RECT 758.270 115.720 759.730 119.670 ;
        RECT 760.570 115.720 762.030 119.670 ;
        RECT 762.870 115.720 764.330 119.670 ;
        RECT 765.170 115.720 766.170 119.670 ;
        RECT 767.010 115.720 768.470 119.670 ;
        RECT 769.310 115.720 770.770 119.670 ;
        RECT 771.610 115.720 773.070 119.670 ;
        RECT 773.910 115.720 775.370 119.670 ;
        RECT 776.210 115.720 777.670 119.670 ;
        RECT 778.510 115.720 779.970 119.670 ;
        RECT 780.810 115.720 781.810 119.670 ;
        RECT 782.650 115.720 784.110 119.670 ;
        RECT 784.950 115.720 786.410 119.670 ;
        RECT 787.250 115.720 788.710 119.670 ;
        RECT 789.550 115.720 791.010 119.670 ;
        RECT 791.850 115.720 793.310 119.670 ;
        RECT 794.150 115.720 795.150 119.670 ;
        RECT 795.990 115.720 797.450 119.670 ;
        RECT 798.290 115.720 799.750 119.670 ;
        RECT 800.590 115.720 802.050 119.670 ;
        RECT 802.890 115.720 804.350 119.670 ;
        RECT 805.190 115.720 806.650 119.670 ;
        RECT 807.490 115.720 808.490 119.670 ;
        RECT 809.330 115.720 810.790 119.670 ;
        RECT 811.630 115.720 813.090 119.670 ;
        RECT 813.930 115.720 815.390 119.670 ;
        RECT 816.230 115.720 817.690 119.670 ;
        RECT 818.530 115.720 819.990 119.670 ;
        RECT 820.830 115.720 821.830 119.670 ;
        RECT 822.670 115.720 824.130 119.670 ;
        RECT 824.970 115.720 826.430 119.670 ;
        RECT 827.270 115.720 828.730 119.670 ;
        RECT 829.570 115.720 831.030 119.670 ;
        RECT 831.870 115.720 833.330 119.670 ;
        RECT 834.170 115.720 835.630 119.670 ;
        RECT 836.470 115.720 837.470 119.670 ;
        RECT 838.310 115.720 839.770 119.670 ;
        RECT 840.610 115.720 842.070 119.670 ;
        RECT 842.910 115.720 844.370 119.670 ;
        RECT 845.210 115.720 846.670 119.670 ;
        RECT 847.510 115.720 848.970 119.670 ;
        RECT 849.810 115.720 850.810 119.670 ;
        RECT 851.650 115.720 853.110 119.670 ;
        RECT 853.950 115.720 855.410 119.670 ;
        RECT 856.250 115.720 857.710 119.670 ;
        RECT 858.550 115.720 860.010 119.670 ;
        RECT 860.850 115.720 862.310 119.670 ;
        RECT 863.150 115.720 864.150 119.670 ;
        RECT 864.990 115.720 866.450 119.670 ;
        RECT 867.290 115.720 868.750 119.670 ;
        RECT 869.590 115.720 871.050 119.670 ;
        RECT 871.890 115.720 873.350 119.670 ;
        RECT 874.190 115.720 875.650 119.670 ;
        RECT 876.490 115.720 877.490 119.670 ;
        RECT 878.330 115.720 879.790 119.670 ;
        RECT 880.630 115.720 882.090 119.670 ;
        RECT 882.930 115.720 884.390 119.670 ;
        RECT 885.230 115.720 886.690 119.670 ;
        RECT 887.530 115.720 888.990 119.670 ;
        RECT 889.830 115.720 891.290 119.670 ;
        RECT 892.130 115.720 893.130 119.670 ;
        RECT 893.970 115.720 895.430 119.670 ;
        RECT 896.270 115.720 897.730 119.670 ;
        RECT 898.570 115.720 900.030 119.670 ;
        RECT 900.870 115.720 902.330 119.670 ;
        RECT 903.170 115.720 904.630 119.670 ;
        RECT 905.470 115.720 906.470 119.670 ;
        RECT 907.310 115.720 908.770 119.670 ;
        RECT 909.610 115.720 911.070 119.670 ;
        RECT 911.910 115.720 913.370 119.670 ;
        RECT 914.210 115.720 915.670 119.670 ;
        RECT 916.510 115.720 917.970 119.670 ;
        RECT 918.810 115.720 919.810 119.670 ;
        RECT 920.650 115.720 922.110 119.670 ;
        RECT 922.950 115.720 924.410 119.670 ;
        RECT 925.250 115.720 926.710 119.670 ;
        RECT 927.550 115.720 929.010 119.670 ;
        RECT 929.850 115.720 931.310 119.670 ;
        RECT 932.150 115.720 933.150 119.670 ;
        RECT 933.990 115.720 935.450 119.670 ;
        RECT 936.290 115.720 937.750 119.670 ;
        RECT 938.590 115.720 940.050 119.670 ;
        RECT 940.890 115.720 942.350 119.670 ;
        RECT 943.190 115.720 944.650 119.670 ;
        RECT 945.490 115.720 946.950 119.670 ;
        RECT 947.790 115.720 948.790 119.670 ;
        RECT 949.630 115.720 951.090 119.670 ;
        RECT 951.930 115.720 953.390 119.670 ;
        RECT 954.230 115.720 955.690 119.670 ;
        RECT 956.530 115.720 957.990 119.670 ;
        RECT 958.830 115.720 960.290 119.670 ;
        RECT 961.130 115.720 962.130 119.670 ;
        RECT 962.970 115.720 964.430 119.670 ;
        RECT 965.270 115.720 966.730 119.670 ;
        RECT 967.570 115.720 969.030 119.670 ;
        RECT 969.870 115.720 971.330 119.670 ;
        RECT 972.170 115.720 973.630 119.670 ;
        RECT 974.470 115.720 975.470 119.670 ;
        RECT 976.310 115.720 977.770 119.670 ;
        RECT 978.610 115.720 980.070 119.670 ;
        RECT 980.910 115.720 982.370 119.670 ;
        RECT 983.210 115.720 984.670 119.670 ;
        RECT 985.510 115.720 986.970 119.670 ;
        RECT 987.810 115.720 988.810 119.670 ;
        RECT 989.650 115.720 991.110 119.670 ;
        RECT 991.950 115.720 993.410 119.670 ;
        RECT 994.250 115.720 995.710 119.670 ;
        RECT 996.550 115.720 998.010 119.670 ;
        RECT 998.850 115.720 1000.310 119.670 ;
        RECT 1001.150 115.720 1002.610 119.670 ;
        RECT 1003.450 115.720 1004.450 119.670 ;
        RECT 1005.290 115.720 1006.750 119.670 ;
        RECT 1007.590 115.720 1009.050 119.670 ;
        RECT 1009.890 115.720 1011.350 119.670 ;
        RECT 1012.190 115.720 1013.650 119.670 ;
        RECT 1014.490 115.720 1015.950 119.670 ;
        RECT 1016.790 115.720 1017.790 119.670 ;
        RECT 1018.630 115.720 1020.090 119.670 ;
        RECT 1020.930 115.720 1022.390 119.670 ;
        RECT 1023.230 115.720 1024.690 119.670 ;
        RECT 1025.530 115.720 1026.990 119.670 ;
        RECT 1027.830 115.720 1029.290 119.670 ;
        RECT 1030.130 115.720 1031.130 119.670 ;
        RECT 1031.970 115.720 1033.430 119.670 ;
        RECT 1034.270 115.720 1035.730 119.670 ;
        RECT 1036.570 115.720 1038.030 119.670 ;
        RECT 1038.870 115.720 1040.330 119.670 ;
        RECT 1041.170 115.720 1042.630 119.670 ;
        RECT 1043.470 115.720 1044.470 119.670 ;
        RECT 1045.310 115.720 1046.770 119.670 ;
        RECT 1047.610 115.720 1049.070 119.670 ;
        RECT 1049.910 115.720 1051.370 119.670 ;
        RECT 1052.210 115.720 1053.670 119.670 ;
        RECT 1054.510 115.720 1055.970 119.670 ;
        RECT 1056.810 115.720 1058.270 119.670 ;
        RECT 1059.110 115.720 1060.110 119.670 ;
        RECT 1060.950 115.720 1062.410 119.670 ;
        RECT 1063.250 115.720 1064.710 119.670 ;
        RECT 1065.550 115.720 1067.010 119.670 ;
        RECT 1067.850 115.720 1069.310 119.670 ;
        RECT 1070.150 115.720 1071.610 119.670 ;
        RECT 1072.450 115.720 1073.450 119.670 ;
        RECT 1074.290 115.720 1075.750 119.670 ;
        RECT 1076.590 115.720 1078.050 119.670 ;
        RECT 1078.890 115.720 1080.350 119.670 ;
        RECT 1081.190 115.720 1082.650 119.670 ;
        RECT 1083.490 115.720 1084.950 119.670 ;
        RECT 1085.790 115.720 1086.790 119.670 ;
        RECT 1087.630 115.720 1089.090 119.670 ;
        RECT 1089.930 115.720 1091.390 119.670 ;
        RECT 1092.230 115.720 1093.690 119.670 ;
        RECT 1094.530 115.720 1095.990 119.670 ;
        RECT 1096.830 115.720 1098.290 119.670 ;
        RECT 0.560 4.280 1098.840 115.720 ;
        RECT 1.110 0.010 1.650 4.280 ;
        RECT 2.490 0.010 3.490 4.280 ;
        RECT 4.330 0.010 5.330 4.280 ;
        RECT 6.170 0.010 7.170 4.280 ;
        RECT 8.010 0.010 9.010 4.280 ;
        RECT 9.850 0.010 10.850 4.280 ;
        RECT 11.690 0.010 12.690 4.280 ;
        RECT 13.530 0.010 14.530 4.280 ;
        RECT 15.370 0.010 15.910 4.280 ;
        RECT 16.750 0.010 17.750 4.280 ;
        RECT 18.590 0.010 19.590 4.280 ;
        RECT 20.430 0.010 21.430 4.280 ;
        RECT 22.270 0.010 23.270 4.280 ;
        RECT 24.110 0.010 25.110 4.280 ;
        RECT 25.950 0.010 26.950 4.280 ;
        RECT 27.790 0.010 28.790 4.280 ;
        RECT 29.630 0.010 30.170 4.280 ;
        RECT 31.010 0.010 32.010 4.280 ;
        RECT 32.850 0.010 33.850 4.280 ;
        RECT 34.690 0.010 35.690 4.280 ;
        RECT 36.530 0.010 37.530 4.280 ;
        RECT 38.370 0.010 39.370 4.280 ;
        RECT 40.210 0.010 41.210 4.280 ;
        RECT 42.050 0.010 43.050 4.280 ;
        RECT 43.890 0.010 44.430 4.280 ;
        RECT 45.270 0.010 46.270 4.280 ;
        RECT 47.110 0.010 48.110 4.280 ;
        RECT 48.950 0.010 49.950 4.280 ;
        RECT 50.790 0.010 51.790 4.280 ;
        RECT 52.630 0.010 53.630 4.280 ;
        RECT 54.470 0.010 55.470 4.280 ;
        RECT 56.310 0.010 57.310 4.280 ;
        RECT 58.150 0.010 58.690 4.280 ;
        RECT 59.530 0.010 60.530 4.280 ;
        RECT 61.370 0.010 62.370 4.280 ;
        RECT 63.210 0.010 64.210 4.280 ;
        RECT 65.050 0.010 66.050 4.280 ;
        RECT 66.890 0.010 67.890 4.280 ;
        RECT 68.730 0.010 69.730 4.280 ;
        RECT 70.570 0.010 71.570 4.280 ;
        RECT 72.410 0.010 72.950 4.280 ;
        RECT 73.790 0.010 74.790 4.280 ;
        RECT 75.630 0.010 76.630 4.280 ;
        RECT 77.470 0.010 78.470 4.280 ;
        RECT 79.310 0.010 80.310 4.280 ;
        RECT 81.150 0.010 82.150 4.280 ;
        RECT 82.990 0.010 83.990 4.280 ;
        RECT 84.830 0.010 85.830 4.280 ;
        RECT 86.670 0.010 87.210 4.280 ;
        RECT 88.050 0.010 89.050 4.280 ;
        RECT 89.890 0.010 90.890 4.280 ;
        RECT 91.730 0.010 92.730 4.280 ;
        RECT 93.570 0.010 94.570 4.280 ;
        RECT 95.410 0.010 96.410 4.280 ;
        RECT 97.250 0.010 98.250 4.280 ;
        RECT 99.090 0.010 100.090 4.280 ;
        RECT 100.930 0.010 101.470 4.280 ;
        RECT 102.310 0.010 103.310 4.280 ;
        RECT 104.150 0.010 105.150 4.280 ;
        RECT 105.990 0.010 106.990 4.280 ;
        RECT 107.830 0.010 108.830 4.280 ;
        RECT 109.670 0.010 110.670 4.280 ;
        RECT 111.510 0.010 112.510 4.280 ;
        RECT 113.350 0.010 114.350 4.280 ;
        RECT 115.190 0.010 115.730 4.280 ;
        RECT 116.570 0.010 117.570 4.280 ;
        RECT 118.410 0.010 119.410 4.280 ;
        RECT 120.250 0.010 121.250 4.280 ;
        RECT 122.090 0.010 123.090 4.280 ;
        RECT 123.930 0.010 124.930 4.280 ;
        RECT 125.770 0.010 126.770 4.280 ;
        RECT 127.610 0.010 128.610 4.280 ;
        RECT 129.450 0.010 129.990 4.280 ;
        RECT 130.830 0.010 131.830 4.280 ;
        RECT 132.670 0.010 133.670 4.280 ;
        RECT 134.510 0.010 135.510 4.280 ;
        RECT 136.350 0.010 137.350 4.280 ;
        RECT 138.190 0.010 139.190 4.280 ;
        RECT 140.030 0.010 141.030 4.280 ;
        RECT 141.870 0.010 142.870 4.280 ;
        RECT 143.710 0.010 144.250 4.280 ;
        RECT 145.090 0.010 146.090 4.280 ;
        RECT 146.930 0.010 147.930 4.280 ;
        RECT 148.770 0.010 149.770 4.280 ;
        RECT 150.610 0.010 151.610 4.280 ;
        RECT 152.450 0.010 153.450 4.280 ;
        RECT 154.290 0.010 155.290 4.280 ;
        RECT 156.130 0.010 157.130 4.280 ;
        RECT 157.970 0.010 158.510 4.280 ;
        RECT 159.350 0.010 160.350 4.280 ;
        RECT 161.190 0.010 162.190 4.280 ;
        RECT 163.030 0.010 164.030 4.280 ;
        RECT 164.870 0.010 165.870 4.280 ;
        RECT 166.710 0.010 167.710 4.280 ;
        RECT 168.550 0.010 169.550 4.280 ;
        RECT 170.390 0.010 171.390 4.280 ;
        RECT 172.230 0.010 172.770 4.280 ;
        RECT 173.610 0.010 174.610 4.280 ;
        RECT 175.450 0.010 176.450 4.280 ;
        RECT 177.290 0.010 178.290 4.280 ;
        RECT 179.130 0.010 180.130 4.280 ;
        RECT 180.970 0.010 181.970 4.280 ;
        RECT 182.810 0.010 183.810 4.280 ;
        RECT 184.650 0.010 185.650 4.280 ;
        RECT 186.490 0.010 187.030 4.280 ;
        RECT 187.870 0.010 188.870 4.280 ;
        RECT 189.710 0.010 190.710 4.280 ;
        RECT 191.550 0.010 192.550 4.280 ;
        RECT 193.390 0.010 194.390 4.280 ;
        RECT 195.230 0.010 196.230 4.280 ;
        RECT 197.070 0.010 198.070 4.280 ;
        RECT 198.910 0.010 199.910 4.280 ;
        RECT 200.750 0.010 201.290 4.280 ;
        RECT 202.130 0.010 203.130 4.280 ;
        RECT 203.970 0.010 204.970 4.280 ;
        RECT 205.810 0.010 206.810 4.280 ;
        RECT 207.650 0.010 208.650 4.280 ;
        RECT 209.490 0.010 210.490 4.280 ;
        RECT 211.330 0.010 212.330 4.280 ;
        RECT 213.170 0.010 214.170 4.280 ;
        RECT 215.010 0.010 215.550 4.280 ;
        RECT 216.390 0.010 217.390 4.280 ;
        RECT 218.230 0.010 219.230 4.280 ;
        RECT 220.070 0.010 221.070 4.280 ;
        RECT 221.910 0.010 222.910 4.280 ;
        RECT 223.750 0.010 224.750 4.280 ;
        RECT 225.590 0.010 226.590 4.280 ;
        RECT 227.430 0.010 228.430 4.280 ;
        RECT 229.270 0.010 229.810 4.280 ;
        RECT 230.650 0.010 231.650 4.280 ;
        RECT 232.490 0.010 233.490 4.280 ;
        RECT 234.330 0.010 235.330 4.280 ;
        RECT 236.170 0.010 237.170 4.280 ;
        RECT 238.010 0.010 239.010 4.280 ;
        RECT 239.850 0.010 240.850 4.280 ;
        RECT 241.690 0.010 242.690 4.280 ;
        RECT 243.530 0.010 244.070 4.280 ;
        RECT 244.910 0.010 245.910 4.280 ;
        RECT 246.750 0.010 247.750 4.280 ;
        RECT 248.590 0.010 249.590 4.280 ;
        RECT 250.430 0.010 251.430 4.280 ;
        RECT 252.270 0.010 253.270 4.280 ;
        RECT 254.110 0.010 255.110 4.280 ;
        RECT 255.950 0.010 256.950 4.280 ;
        RECT 257.790 0.010 258.330 4.280 ;
        RECT 259.170 0.010 260.170 4.280 ;
        RECT 261.010 0.010 262.010 4.280 ;
        RECT 262.850 0.010 263.850 4.280 ;
        RECT 264.690 0.010 265.690 4.280 ;
        RECT 266.530 0.010 267.530 4.280 ;
        RECT 268.370 0.010 269.370 4.280 ;
        RECT 270.210 0.010 271.210 4.280 ;
        RECT 272.050 0.010 272.590 4.280 ;
        RECT 273.430 0.010 274.430 4.280 ;
        RECT 275.270 0.010 276.270 4.280 ;
        RECT 277.110 0.010 278.110 4.280 ;
        RECT 278.950 0.010 279.950 4.280 ;
        RECT 280.790 0.010 281.790 4.280 ;
        RECT 282.630 0.010 283.630 4.280 ;
        RECT 284.470 0.010 285.470 4.280 ;
        RECT 286.310 0.010 286.850 4.280 ;
        RECT 287.690 0.010 288.690 4.280 ;
        RECT 289.530 0.010 290.530 4.280 ;
        RECT 291.370 0.010 292.370 4.280 ;
        RECT 293.210 0.010 294.210 4.280 ;
        RECT 295.050 0.010 296.050 4.280 ;
        RECT 296.890 0.010 297.890 4.280 ;
        RECT 298.730 0.010 299.730 4.280 ;
        RECT 300.570 0.010 301.110 4.280 ;
        RECT 301.950 0.010 302.950 4.280 ;
        RECT 303.790 0.010 304.790 4.280 ;
        RECT 305.630 0.010 306.630 4.280 ;
        RECT 307.470 0.010 308.470 4.280 ;
        RECT 309.310 0.010 310.310 4.280 ;
        RECT 311.150 0.010 312.150 4.280 ;
        RECT 312.990 0.010 313.990 4.280 ;
        RECT 314.830 0.010 315.370 4.280 ;
        RECT 316.210 0.010 317.210 4.280 ;
        RECT 318.050 0.010 319.050 4.280 ;
        RECT 319.890 0.010 320.890 4.280 ;
        RECT 321.730 0.010 322.730 4.280 ;
        RECT 323.570 0.010 324.570 4.280 ;
        RECT 325.410 0.010 326.410 4.280 ;
        RECT 327.250 0.010 328.250 4.280 ;
        RECT 329.090 0.010 329.630 4.280 ;
        RECT 330.470 0.010 331.470 4.280 ;
        RECT 332.310 0.010 333.310 4.280 ;
        RECT 334.150 0.010 335.150 4.280 ;
        RECT 335.990 0.010 336.990 4.280 ;
        RECT 337.830 0.010 338.830 4.280 ;
        RECT 339.670 0.010 340.670 4.280 ;
        RECT 341.510 0.010 342.510 4.280 ;
        RECT 343.350 0.010 343.890 4.280 ;
        RECT 344.730 0.010 345.730 4.280 ;
        RECT 346.570 0.010 347.570 4.280 ;
        RECT 348.410 0.010 349.410 4.280 ;
        RECT 350.250 0.010 351.250 4.280 ;
        RECT 352.090 0.010 353.090 4.280 ;
        RECT 353.930 0.010 354.930 4.280 ;
        RECT 355.770 0.010 356.770 4.280 ;
        RECT 357.610 0.010 358.150 4.280 ;
        RECT 358.990 0.010 359.990 4.280 ;
        RECT 360.830 0.010 361.830 4.280 ;
        RECT 362.670 0.010 363.670 4.280 ;
        RECT 364.510 0.010 365.510 4.280 ;
        RECT 366.350 0.010 367.350 4.280 ;
        RECT 368.190 0.010 369.190 4.280 ;
        RECT 370.030 0.010 371.030 4.280 ;
        RECT 371.870 0.010 372.410 4.280 ;
        RECT 373.250 0.010 374.250 4.280 ;
        RECT 375.090 0.010 376.090 4.280 ;
        RECT 376.930 0.010 377.930 4.280 ;
        RECT 378.770 0.010 379.770 4.280 ;
        RECT 380.610 0.010 381.610 4.280 ;
        RECT 382.450 0.010 383.450 4.280 ;
        RECT 384.290 0.010 385.290 4.280 ;
        RECT 386.130 0.010 386.670 4.280 ;
        RECT 387.510 0.010 388.510 4.280 ;
        RECT 389.350 0.010 390.350 4.280 ;
        RECT 391.190 0.010 392.190 4.280 ;
        RECT 393.030 0.010 394.030 4.280 ;
        RECT 394.870 0.010 395.870 4.280 ;
        RECT 396.710 0.010 397.710 4.280 ;
        RECT 398.550 0.010 399.550 4.280 ;
        RECT 400.390 0.010 400.930 4.280 ;
        RECT 401.770 0.010 402.770 4.280 ;
        RECT 403.610 0.010 404.610 4.280 ;
        RECT 405.450 0.010 406.450 4.280 ;
        RECT 407.290 0.010 408.290 4.280 ;
        RECT 409.130 0.010 410.130 4.280 ;
        RECT 410.970 0.010 411.970 4.280 ;
        RECT 412.810 0.010 413.810 4.280 ;
        RECT 414.650 0.010 415.190 4.280 ;
        RECT 416.030 0.010 417.030 4.280 ;
        RECT 417.870 0.010 418.870 4.280 ;
        RECT 419.710 0.010 420.710 4.280 ;
        RECT 421.550 0.010 422.550 4.280 ;
        RECT 423.390 0.010 424.390 4.280 ;
        RECT 425.230 0.010 426.230 4.280 ;
        RECT 427.070 0.010 428.070 4.280 ;
        RECT 428.910 0.010 429.450 4.280 ;
        RECT 430.290 0.010 431.290 4.280 ;
        RECT 432.130 0.010 433.130 4.280 ;
        RECT 433.970 0.010 434.970 4.280 ;
        RECT 435.810 0.010 436.810 4.280 ;
        RECT 437.650 0.010 438.650 4.280 ;
        RECT 439.490 0.010 440.490 4.280 ;
        RECT 441.330 0.010 442.330 4.280 ;
        RECT 443.170 0.010 443.710 4.280 ;
        RECT 444.550 0.010 445.550 4.280 ;
        RECT 446.390 0.010 447.390 4.280 ;
        RECT 448.230 0.010 449.230 4.280 ;
        RECT 450.070 0.010 451.070 4.280 ;
        RECT 451.910 0.010 452.910 4.280 ;
        RECT 453.750 0.010 454.750 4.280 ;
        RECT 455.590 0.010 456.590 4.280 ;
        RECT 457.430 0.010 457.970 4.280 ;
        RECT 458.810 0.010 459.810 4.280 ;
        RECT 460.650 0.010 461.650 4.280 ;
        RECT 462.490 0.010 463.490 4.280 ;
        RECT 464.330 0.010 465.330 4.280 ;
        RECT 466.170 0.010 467.170 4.280 ;
        RECT 468.010 0.010 469.010 4.280 ;
        RECT 469.850 0.010 470.850 4.280 ;
        RECT 471.690 0.010 472.230 4.280 ;
        RECT 473.070 0.010 474.070 4.280 ;
        RECT 474.910 0.010 475.910 4.280 ;
        RECT 476.750 0.010 477.750 4.280 ;
        RECT 478.590 0.010 479.590 4.280 ;
        RECT 480.430 0.010 481.430 4.280 ;
        RECT 482.270 0.010 483.270 4.280 ;
        RECT 484.110 0.010 485.110 4.280 ;
        RECT 485.950 0.010 486.490 4.280 ;
        RECT 487.330 0.010 488.330 4.280 ;
        RECT 489.170 0.010 490.170 4.280 ;
        RECT 491.010 0.010 492.010 4.280 ;
        RECT 492.850 0.010 493.850 4.280 ;
        RECT 494.690 0.010 495.690 4.280 ;
        RECT 496.530 0.010 497.530 4.280 ;
        RECT 498.370 0.010 499.370 4.280 ;
        RECT 500.210 0.010 500.750 4.280 ;
        RECT 501.590 0.010 502.590 4.280 ;
        RECT 503.430 0.010 504.430 4.280 ;
        RECT 505.270 0.010 506.270 4.280 ;
        RECT 507.110 0.010 508.110 4.280 ;
        RECT 508.950 0.010 509.950 4.280 ;
        RECT 510.790 0.010 511.790 4.280 ;
        RECT 512.630 0.010 513.630 4.280 ;
        RECT 514.470 0.010 515.010 4.280 ;
        RECT 515.850 0.010 516.850 4.280 ;
        RECT 517.690 0.010 518.690 4.280 ;
        RECT 519.530 0.010 520.530 4.280 ;
        RECT 521.370 0.010 522.370 4.280 ;
        RECT 523.210 0.010 524.210 4.280 ;
        RECT 525.050 0.010 526.050 4.280 ;
        RECT 526.890 0.010 527.890 4.280 ;
        RECT 528.730 0.010 529.270 4.280 ;
        RECT 530.110 0.010 531.110 4.280 ;
        RECT 531.950 0.010 532.950 4.280 ;
        RECT 533.790 0.010 534.790 4.280 ;
        RECT 535.630 0.010 536.630 4.280 ;
        RECT 537.470 0.010 538.470 4.280 ;
        RECT 539.310 0.010 540.310 4.280 ;
        RECT 541.150 0.010 542.150 4.280 ;
        RECT 542.990 0.010 543.530 4.280 ;
        RECT 544.370 0.010 545.370 4.280 ;
        RECT 546.210 0.010 547.210 4.280 ;
        RECT 548.050 0.010 549.050 4.280 ;
        RECT 549.890 0.010 550.890 4.280 ;
        RECT 551.730 0.010 552.730 4.280 ;
        RECT 553.570 0.010 554.570 4.280 ;
        RECT 555.410 0.010 556.410 4.280 ;
        RECT 557.250 0.010 557.790 4.280 ;
        RECT 558.630 0.010 559.630 4.280 ;
        RECT 560.470 0.010 561.470 4.280 ;
        RECT 562.310 0.010 563.310 4.280 ;
        RECT 564.150 0.010 565.150 4.280 ;
        RECT 565.990 0.010 566.990 4.280 ;
        RECT 567.830 0.010 568.830 4.280 ;
        RECT 569.670 0.010 570.670 4.280 ;
        RECT 571.510 0.010 572.050 4.280 ;
        RECT 572.890 0.010 573.890 4.280 ;
        RECT 574.730 0.010 575.730 4.280 ;
        RECT 576.570 0.010 577.570 4.280 ;
        RECT 578.410 0.010 579.410 4.280 ;
        RECT 580.250 0.010 581.250 4.280 ;
        RECT 582.090 0.010 583.090 4.280 ;
        RECT 583.930 0.010 584.930 4.280 ;
        RECT 585.770 0.010 586.310 4.280 ;
        RECT 587.150 0.010 588.150 4.280 ;
        RECT 588.990 0.010 589.990 4.280 ;
        RECT 590.830 0.010 591.830 4.280 ;
        RECT 592.670 0.010 593.670 4.280 ;
        RECT 594.510 0.010 595.510 4.280 ;
        RECT 596.350 0.010 597.350 4.280 ;
        RECT 598.190 0.010 599.190 4.280 ;
        RECT 600.030 0.010 600.570 4.280 ;
        RECT 601.410 0.010 602.410 4.280 ;
        RECT 603.250 0.010 604.250 4.280 ;
        RECT 605.090 0.010 606.090 4.280 ;
        RECT 606.930 0.010 607.930 4.280 ;
        RECT 608.770 0.010 609.770 4.280 ;
        RECT 610.610 0.010 611.610 4.280 ;
        RECT 612.450 0.010 613.450 4.280 ;
        RECT 614.290 0.010 614.830 4.280 ;
        RECT 615.670 0.010 616.670 4.280 ;
        RECT 617.510 0.010 618.510 4.280 ;
        RECT 619.350 0.010 620.350 4.280 ;
        RECT 621.190 0.010 622.190 4.280 ;
        RECT 623.030 0.010 624.030 4.280 ;
        RECT 624.870 0.010 625.870 4.280 ;
        RECT 626.710 0.010 627.710 4.280 ;
        RECT 628.550 0.010 629.090 4.280 ;
        RECT 629.930 0.010 630.930 4.280 ;
        RECT 631.770 0.010 632.770 4.280 ;
        RECT 633.610 0.010 634.610 4.280 ;
        RECT 635.450 0.010 636.450 4.280 ;
        RECT 637.290 0.010 638.290 4.280 ;
        RECT 639.130 0.010 640.130 4.280 ;
        RECT 640.970 0.010 641.970 4.280 ;
        RECT 642.810 0.010 643.350 4.280 ;
        RECT 644.190 0.010 645.190 4.280 ;
        RECT 646.030 0.010 647.030 4.280 ;
        RECT 647.870 0.010 648.870 4.280 ;
        RECT 649.710 0.010 650.710 4.280 ;
        RECT 651.550 0.010 652.550 4.280 ;
        RECT 653.390 0.010 654.390 4.280 ;
        RECT 655.230 0.010 656.230 4.280 ;
        RECT 657.070 0.010 657.610 4.280 ;
        RECT 658.450 0.010 659.450 4.280 ;
        RECT 660.290 0.010 661.290 4.280 ;
        RECT 662.130 0.010 663.130 4.280 ;
        RECT 663.970 0.010 664.970 4.280 ;
        RECT 665.810 0.010 666.810 4.280 ;
        RECT 667.650 0.010 668.650 4.280 ;
        RECT 669.490 0.010 670.490 4.280 ;
        RECT 671.330 0.010 671.870 4.280 ;
        RECT 672.710 0.010 673.710 4.280 ;
        RECT 674.550 0.010 675.550 4.280 ;
        RECT 676.390 0.010 677.390 4.280 ;
        RECT 678.230 0.010 679.230 4.280 ;
        RECT 680.070 0.010 681.070 4.280 ;
        RECT 681.910 0.010 682.910 4.280 ;
        RECT 683.750 0.010 684.750 4.280 ;
        RECT 685.590 0.010 686.130 4.280 ;
        RECT 686.970 0.010 687.970 4.280 ;
        RECT 688.810 0.010 689.810 4.280 ;
        RECT 690.650 0.010 691.650 4.280 ;
        RECT 692.490 0.010 693.490 4.280 ;
        RECT 694.330 0.010 695.330 4.280 ;
        RECT 696.170 0.010 697.170 4.280 ;
        RECT 698.010 0.010 699.010 4.280 ;
        RECT 699.850 0.010 700.390 4.280 ;
        RECT 701.230 0.010 702.230 4.280 ;
        RECT 703.070 0.010 704.070 4.280 ;
        RECT 704.910 0.010 705.910 4.280 ;
        RECT 706.750 0.010 707.750 4.280 ;
        RECT 708.590 0.010 709.590 4.280 ;
        RECT 710.430 0.010 711.430 4.280 ;
        RECT 712.270 0.010 713.270 4.280 ;
        RECT 714.110 0.010 714.650 4.280 ;
        RECT 715.490 0.010 716.490 4.280 ;
        RECT 717.330 0.010 718.330 4.280 ;
        RECT 719.170 0.010 720.170 4.280 ;
        RECT 721.010 0.010 722.010 4.280 ;
        RECT 722.850 0.010 723.850 4.280 ;
        RECT 724.690 0.010 725.690 4.280 ;
        RECT 726.530 0.010 727.530 4.280 ;
        RECT 728.370 0.010 728.910 4.280 ;
        RECT 729.750 0.010 730.750 4.280 ;
        RECT 731.590 0.010 732.590 4.280 ;
        RECT 733.430 0.010 734.430 4.280 ;
        RECT 735.270 0.010 736.270 4.280 ;
        RECT 737.110 0.010 738.110 4.280 ;
        RECT 738.950 0.010 739.950 4.280 ;
        RECT 740.790 0.010 741.790 4.280 ;
        RECT 742.630 0.010 743.170 4.280 ;
        RECT 744.010 0.010 745.010 4.280 ;
        RECT 745.850 0.010 746.850 4.280 ;
        RECT 747.690 0.010 748.690 4.280 ;
        RECT 749.530 0.010 750.530 4.280 ;
        RECT 751.370 0.010 752.370 4.280 ;
        RECT 753.210 0.010 754.210 4.280 ;
        RECT 755.050 0.010 756.050 4.280 ;
        RECT 756.890 0.010 757.430 4.280 ;
        RECT 758.270 0.010 759.270 4.280 ;
        RECT 760.110 0.010 761.110 4.280 ;
        RECT 761.950 0.010 762.950 4.280 ;
        RECT 763.790 0.010 764.790 4.280 ;
        RECT 765.630 0.010 766.630 4.280 ;
        RECT 767.470 0.010 768.470 4.280 ;
        RECT 769.310 0.010 770.310 4.280 ;
        RECT 771.150 0.010 771.690 4.280 ;
        RECT 772.530 0.010 773.530 4.280 ;
        RECT 774.370 0.010 775.370 4.280 ;
        RECT 776.210 0.010 777.210 4.280 ;
        RECT 778.050 0.010 779.050 4.280 ;
        RECT 779.890 0.010 780.890 4.280 ;
        RECT 781.730 0.010 782.730 4.280 ;
        RECT 783.570 0.010 784.570 4.280 ;
        RECT 785.410 0.010 785.950 4.280 ;
        RECT 786.790 0.010 787.790 4.280 ;
        RECT 788.630 0.010 789.630 4.280 ;
        RECT 790.470 0.010 791.470 4.280 ;
        RECT 792.310 0.010 793.310 4.280 ;
        RECT 794.150 0.010 795.150 4.280 ;
        RECT 795.990 0.010 796.990 4.280 ;
        RECT 797.830 0.010 798.830 4.280 ;
        RECT 799.670 0.010 800.210 4.280 ;
        RECT 801.050 0.010 802.050 4.280 ;
        RECT 802.890 0.010 803.890 4.280 ;
        RECT 804.730 0.010 805.730 4.280 ;
        RECT 806.570 0.010 807.570 4.280 ;
        RECT 808.410 0.010 809.410 4.280 ;
        RECT 810.250 0.010 811.250 4.280 ;
        RECT 812.090 0.010 813.090 4.280 ;
        RECT 813.930 0.010 814.470 4.280 ;
        RECT 815.310 0.010 816.310 4.280 ;
        RECT 817.150 0.010 818.150 4.280 ;
        RECT 818.990 0.010 819.990 4.280 ;
        RECT 820.830 0.010 821.830 4.280 ;
        RECT 822.670 0.010 823.670 4.280 ;
        RECT 824.510 0.010 825.510 4.280 ;
        RECT 826.350 0.010 827.350 4.280 ;
        RECT 828.190 0.010 828.730 4.280 ;
        RECT 829.570 0.010 830.570 4.280 ;
        RECT 831.410 0.010 832.410 4.280 ;
        RECT 833.250 0.010 834.250 4.280 ;
        RECT 835.090 0.010 836.090 4.280 ;
        RECT 836.930 0.010 837.930 4.280 ;
        RECT 838.770 0.010 839.770 4.280 ;
        RECT 840.610 0.010 841.610 4.280 ;
        RECT 842.450 0.010 842.990 4.280 ;
        RECT 843.830 0.010 844.830 4.280 ;
        RECT 845.670 0.010 846.670 4.280 ;
        RECT 847.510 0.010 848.510 4.280 ;
        RECT 849.350 0.010 850.350 4.280 ;
        RECT 851.190 0.010 852.190 4.280 ;
        RECT 853.030 0.010 854.030 4.280 ;
        RECT 854.870 0.010 855.870 4.280 ;
        RECT 856.710 0.010 857.250 4.280 ;
        RECT 858.090 0.010 859.090 4.280 ;
        RECT 859.930 0.010 860.930 4.280 ;
        RECT 861.770 0.010 862.770 4.280 ;
        RECT 863.610 0.010 864.610 4.280 ;
        RECT 865.450 0.010 866.450 4.280 ;
        RECT 867.290 0.010 868.290 4.280 ;
        RECT 869.130 0.010 870.130 4.280 ;
        RECT 870.970 0.010 871.510 4.280 ;
        RECT 872.350 0.010 873.350 4.280 ;
        RECT 874.190 0.010 875.190 4.280 ;
        RECT 876.030 0.010 877.030 4.280 ;
        RECT 877.870 0.010 878.870 4.280 ;
        RECT 879.710 0.010 880.710 4.280 ;
        RECT 881.550 0.010 882.550 4.280 ;
        RECT 883.390 0.010 884.390 4.280 ;
        RECT 885.230 0.010 885.770 4.280 ;
        RECT 886.610 0.010 887.610 4.280 ;
        RECT 888.450 0.010 889.450 4.280 ;
        RECT 890.290 0.010 891.290 4.280 ;
        RECT 892.130 0.010 893.130 4.280 ;
        RECT 893.970 0.010 894.970 4.280 ;
        RECT 895.810 0.010 896.810 4.280 ;
        RECT 897.650 0.010 898.650 4.280 ;
        RECT 899.490 0.010 900.030 4.280 ;
        RECT 900.870 0.010 901.870 4.280 ;
        RECT 902.710 0.010 903.710 4.280 ;
        RECT 904.550 0.010 905.550 4.280 ;
        RECT 906.390 0.010 907.390 4.280 ;
        RECT 908.230 0.010 909.230 4.280 ;
        RECT 910.070 0.010 911.070 4.280 ;
        RECT 911.910 0.010 912.910 4.280 ;
        RECT 913.750 0.010 914.290 4.280 ;
        RECT 915.130 0.010 916.130 4.280 ;
        RECT 916.970 0.010 917.970 4.280 ;
        RECT 918.810 0.010 919.810 4.280 ;
        RECT 920.650 0.010 921.650 4.280 ;
        RECT 922.490 0.010 923.490 4.280 ;
        RECT 924.330 0.010 925.330 4.280 ;
        RECT 926.170 0.010 927.170 4.280 ;
        RECT 928.010 0.010 928.550 4.280 ;
        RECT 929.390 0.010 930.390 4.280 ;
        RECT 931.230 0.010 932.230 4.280 ;
        RECT 933.070 0.010 934.070 4.280 ;
        RECT 934.910 0.010 935.910 4.280 ;
        RECT 936.750 0.010 937.750 4.280 ;
        RECT 938.590 0.010 939.590 4.280 ;
        RECT 940.430 0.010 941.430 4.280 ;
        RECT 942.270 0.010 942.810 4.280 ;
        RECT 943.650 0.010 944.650 4.280 ;
        RECT 945.490 0.010 946.490 4.280 ;
        RECT 947.330 0.010 948.330 4.280 ;
        RECT 949.170 0.010 950.170 4.280 ;
        RECT 951.010 0.010 952.010 4.280 ;
        RECT 952.850 0.010 953.850 4.280 ;
        RECT 954.690 0.010 955.690 4.280 ;
        RECT 956.530 0.010 957.070 4.280 ;
        RECT 957.910 0.010 958.910 4.280 ;
        RECT 959.750 0.010 960.750 4.280 ;
        RECT 961.590 0.010 962.590 4.280 ;
        RECT 963.430 0.010 964.430 4.280 ;
        RECT 965.270 0.010 966.270 4.280 ;
        RECT 967.110 0.010 968.110 4.280 ;
        RECT 968.950 0.010 969.950 4.280 ;
        RECT 970.790 0.010 971.330 4.280 ;
        RECT 972.170 0.010 973.170 4.280 ;
        RECT 974.010 0.010 975.010 4.280 ;
        RECT 975.850 0.010 976.850 4.280 ;
        RECT 977.690 0.010 978.690 4.280 ;
        RECT 979.530 0.010 980.530 4.280 ;
        RECT 981.370 0.010 982.370 4.280 ;
        RECT 983.210 0.010 984.210 4.280 ;
        RECT 985.050 0.010 985.590 4.280 ;
        RECT 986.430 0.010 987.430 4.280 ;
        RECT 988.270 0.010 989.270 4.280 ;
        RECT 990.110 0.010 991.110 4.280 ;
        RECT 991.950 0.010 992.950 4.280 ;
        RECT 993.790 0.010 994.790 4.280 ;
        RECT 995.630 0.010 996.630 4.280 ;
        RECT 997.470 0.010 998.470 4.280 ;
        RECT 999.310 0.010 999.850 4.280 ;
        RECT 1000.690 0.010 1001.690 4.280 ;
        RECT 1002.530 0.010 1003.530 4.280 ;
        RECT 1004.370 0.010 1005.370 4.280 ;
        RECT 1006.210 0.010 1007.210 4.280 ;
        RECT 1008.050 0.010 1009.050 4.280 ;
        RECT 1009.890 0.010 1010.890 4.280 ;
        RECT 1011.730 0.010 1012.730 4.280 ;
        RECT 1013.570 0.010 1014.110 4.280 ;
        RECT 1014.950 0.010 1015.950 4.280 ;
        RECT 1016.790 0.010 1017.790 4.280 ;
        RECT 1018.630 0.010 1019.630 4.280 ;
        RECT 1020.470 0.010 1021.470 4.280 ;
        RECT 1022.310 0.010 1023.310 4.280 ;
        RECT 1024.150 0.010 1025.150 4.280 ;
        RECT 1025.990 0.010 1026.990 4.280 ;
        RECT 1027.830 0.010 1028.370 4.280 ;
        RECT 1029.210 0.010 1030.210 4.280 ;
        RECT 1031.050 0.010 1032.050 4.280 ;
        RECT 1032.890 0.010 1033.890 4.280 ;
        RECT 1034.730 0.010 1035.730 4.280 ;
        RECT 1036.570 0.010 1037.570 4.280 ;
        RECT 1038.410 0.010 1039.410 4.280 ;
        RECT 1040.250 0.010 1041.250 4.280 ;
        RECT 1042.090 0.010 1042.630 4.280 ;
        RECT 1043.470 0.010 1044.470 4.280 ;
        RECT 1045.310 0.010 1046.310 4.280 ;
        RECT 1047.150 0.010 1048.150 4.280 ;
        RECT 1048.990 0.010 1049.990 4.280 ;
        RECT 1050.830 0.010 1051.830 4.280 ;
        RECT 1052.670 0.010 1053.670 4.280 ;
        RECT 1054.510 0.010 1055.510 4.280 ;
        RECT 1056.350 0.010 1056.890 4.280 ;
        RECT 1057.730 0.010 1058.730 4.280 ;
        RECT 1059.570 0.010 1060.570 4.280 ;
        RECT 1061.410 0.010 1062.410 4.280 ;
        RECT 1063.250 0.010 1064.250 4.280 ;
        RECT 1065.090 0.010 1066.090 4.280 ;
        RECT 1066.930 0.010 1067.930 4.280 ;
        RECT 1068.770 0.010 1069.770 4.280 ;
        RECT 1070.610 0.010 1071.150 4.280 ;
        RECT 1071.990 0.010 1072.990 4.280 ;
        RECT 1073.830 0.010 1074.830 4.280 ;
        RECT 1075.670 0.010 1076.670 4.280 ;
        RECT 1077.510 0.010 1078.510 4.280 ;
        RECT 1079.350 0.010 1080.350 4.280 ;
        RECT 1081.190 0.010 1082.190 4.280 ;
        RECT 1083.030 0.010 1084.030 4.280 ;
        RECT 1084.870 0.010 1085.410 4.280 ;
        RECT 1086.250 0.010 1087.250 4.280 ;
        RECT 1088.090 0.010 1089.090 4.280 ;
        RECT 1089.930 0.010 1090.930 4.280 ;
        RECT 1091.770 0.010 1092.770 4.280 ;
        RECT 1093.610 0.010 1094.610 4.280 ;
        RECT 1095.450 0.010 1096.450 4.280 ;
        RECT 1097.290 0.010 1098.290 4.280 ;
      LAYER met3 ;
        RECT 4.000 113.920 1096.000 119.505 ;
        RECT 4.000 112.520 1095.600 113.920 ;
        RECT 4.000 101.680 1096.000 112.520 ;
        RECT 4.000 100.320 1095.600 101.680 ;
        RECT 4.400 100.280 1095.600 100.320 ;
        RECT 4.400 98.920 1096.000 100.280 ;
        RECT 4.000 90.120 1096.000 98.920 ;
        RECT 4.000 88.720 1095.600 90.120 ;
        RECT 4.000 77.880 1096.000 88.720 ;
        RECT 4.000 76.480 1095.600 77.880 ;
        RECT 4.000 66.320 1096.000 76.480 ;
        RECT 4.000 64.920 1095.600 66.320 ;
        RECT 4.000 60.200 1096.000 64.920 ;
        RECT 4.400 58.800 1096.000 60.200 ;
        RECT 4.000 54.080 1096.000 58.800 ;
        RECT 4.000 52.680 1095.600 54.080 ;
        RECT 4.000 41.840 1096.000 52.680 ;
        RECT 4.000 40.440 1095.600 41.840 ;
        RECT 4.000 30.280 1096.000 40.440 ;
        RECT 4.000 28.880 1095.600 30.280 ;
        RECT 4.000 20.760 1096.000 28.880 ;
        RECT 4.400 19.360 1096.000 20.760 ;
        RECT 4.000 18.040 1096.000 19.360 ;
        RECT 4.000 16.640 1095.600 18.040 ;
        RECT 4.000 6.480 1096.000 16.640 ;
        RECT 4.000 5.080 1095.600 6.480 ;
        RECT 4.000 0.175 1096.000 5.080 ;
      LAYER met4 ;
        RECT 230.295 114.880 1080.705 119.505 ;
        RECT 230.295 4.800 245.420 114.880 ;
        RECT 247.120 114.640 320.670 114.880 ;
        RECT 247.120 5.040 249.520 114.640 ;
        RECT 251.220 5.040 253.620 114.640 ;
        RECT 255.320 5.040 320.670 114.640 ;
        RECT 247.120 4.800 320.670 5.040 ;
        RECT 322.370 114.640 395.920 114.880 ;
        RECT 322.370 5.040 324.770 114.640 ;
        RECT 326.470 5.040 328.870 114.640 ;
        RECT 330.570 5.040 395.920 114.640 ;
        RECT 322.370 4.800 395.920 5.040 ;
        RECT 397.620 114.640 471.170 114.880 ;
        RECT 397.620 5.040 400.020 114.640 ;
        RECT 401.720 5.040 404.120 114.640 ;
        RECT 405.820 5.040 471.170 114.640 ;
        RECT 397.620 4.800 471.170 5.040 ;
        RECT 472.870 114.640 546.420 114.880 ;
        RECT 472.870 5.040 475.270 114.640 ;
        RECT 476.970 5.040 479.370 114.640 ;
        RECT 481.070 5.040 546.420 114.640 ;
        RECT 472.870 4.800 546.420 5.040 ;
        RECT 548.120 114.640 621.670 114.880 ;
        RECT 548.120 5.040 550.520 114.640 ;
        RECT 552.220 5.040 554.620 114.640 ;
        RECT 556.320 5.040 621.670 114.640 ;
        RECT 548.120 4.800 621.670 5.040 ;
        RECT 623.370 114.640 696.920 114.880 ;
        RECT 623.370 5.040 625.770 114.640 ;
        RECT 627.470 5.040 629.870 114.640 ;
        RECT 631.570 5.040 696.920 114.640 ;
        RECT 623.370 4.800 696.920 5.040 ;
        RECT 698.620 114.640 772.170 114.880 ;
        RECT 698.620 5.040 701.020 114.640 ;
        RECT 702.720 5.040 705.120 114.640 ;
        RECT 706.820 5.040 772.170 114.640 ;
        RECT 698.620 4.800 772.170 5.040 ;
        RECT 773.870 114.640 847.420 114.880 ;
        RECT 773.870 5.040 776.270 114.640 ;
        RECT 777.970 5.040 780.370 114.640 ;
        RECT 782.070 5.040 847.420 114.640 ;
        RECT 773.870 4.800 847.420 5.040 ;
        RECT 849.120 114.640 922.670 114.880 ;
        RECT 849.120 5.040 851.520 114.640 ;
        RECT 853.220 5.040 855.620 114.640 ;
        RECT 857.320 5.040 922.670 114.640 ;
        RECT 849.120 4.800 922.670 5.040 ;
        RECT 924.370 114.640 997.920 114.880 ;
        RECT 924.370 5.040 926.770 114.640 ;
        RECT 928.470 5.040 930.870 114.640 ;
        RECT 932.570 5.040 933.670 114.640 ;
        RECT 935.370 5.040 936.670 114.640 ;
        RECT 938.370 5.040 997.920 114.640 ;
        RECT 924.370 4.800 997.920 5.040 ;
        RECT 999.620 114.640 1073.170 114.880 ;
        RECT 999.620 5.040 1002.020 114.640 ;
        RECT 1003.720 5.040 1006.120 114.640 ;
        RECT 1007.820 5.040 1008.920 114.640 ;
        RECT 1010.620 5.040 1011.920 114.640 ;
        RECT 1013.620 5.040 1073.170 114.640 ;
        RECT 999.620 4.800 1073.170 5.040 ;
        RECT 1074.870 114.640 1080.705 114.880 ;
        RECT 1074.870 5.040 1077.270 114.640 ;
        RECT 1078.970 5.040 1080.705 114.640 ;
        RECT 1074.870 4.800 1080.705 5.040 ;
        RECT 230.295 0.175 1080.705 4.800 ;
  END
END mgmt_protect
END LIBRARY

