magic
tech sky130A
magscale 1 2
timestamp 1637275745
<< metal1 >>
rect 425974 1006000 425980 1006052
rect 426032 1006040 426038 1006052
rect 458910 1006040 458916 1006052
rect 426032 1006012 458916 1006040
rect 426032 1006000 426038 1006012
rect 458910 1006000 458916 1006012
rect 458968 1006000 458974 1006052
rect 424318 1005864 424324 1005916
rect 424376 1005904 424382 1005916
rect 440418 1005904 440424 1005916
rect 424376 1005876 440424 1005904
rect 424376 1005864 424382 1005876
rect 440418 1005864 440424 1005876
rect 440476 1005864 440482 1005916
rect 423858 1005796 423864 1005848
rect 423916 1005836 423922 1005848
rect 440234 1005836 440240 1005848
rect 423916 1005808 440240 1005836
rect 423916 1005796 423922 1005808
rect 440234 1005796 440240 1005808
rect 440292 1005796 440298 1005848
rect 504542 1005660 504548 1005712
rect 504600 1005700 504606 1005712
rect 519722 1005700 519728 1005712
rect 504600 1005672 519728 1005700
rect 504600 1005660 504606 1005672
rect 519722 1005660 519728 1005672
rect 519780 1005660 519786 1005712
rect 356054 1005592 356060 1005644
rect 356112 1005632 356118 1005644
rect 373166 1005632 373172 1005644
rect 356112 1005604 373172 1005632
rect 356112 1005592 356118 1005604
rect 373166 1005592 373172 1005604
rect 373224 1005592 373230 1005644
rect 505002 1005592 505008 1005644
rect 505060 1005632 505066 1005644
rect 517422 1005632 517428 1005644
rect 505060 1005604 517428 1005632
rect 505060 1005592 505066 1005604
rect 517422 1005592 517428 1005604
rect 517480 1005592 517486 1005644
rect 356882 1005524 356888 1005576
rect 356940 1005564 356946 1005576
rect 378042 1005564 378048 1005576
rect 356940 1005536 378048 1005564
rect 356940 1005524 356946 1005536
rect 378042 1005524 378048 1005536
rect 378100 1005524 378106 1005576
rect 505370 1005524 505376 1005576
rect 505428 1005564 505434 1005576
rect 518802 1005564 518808 1005576
rect 505428 1005536 518808 1005564
rect 505428 1005524 505434 1005536
rect 518802 1005524 518808 1005536
rect 518860 1005524 518866 1005576
rect 502978 1005456 502984 1005508
rect 503036 1005496 503042 1005508
rect 523034 1005496 523040 1005508
rect 503036 1005468 523040 1005496
rect 503036 1005456 503042 1005468
rect 523034 1005456 523040 1005468
rect 523092 1005456 523098 1005508
rect 144822 1005388 144828 1005440
rect 144880 1005428 144886 1005440
rect 160278 1005428 160284 1005440
rect 144880 1005400 160284 1005428
rect 144880 1005388 144886 1005400
rect 160278 1005388 160284 1005400
rect 160336 1005388 160342 1005440
rect 356514 1005388 356520 1005440
rect 356572 1005428 356578 1005440
rect 376662 1005428 376668 1005440
rect 356572 1005400 376668 1005428
rect 356572 1005388 356578 1005400
rect 376662 1005388 376668 1005400
rect 376720 1005388 376726 1005440
rect 425146 1005388 425152 1005440
rect 425204 1005428 425210 1005440
rect 467926 1005428 467932 1005440
rect 425204 1005400 467932 1005428
rect 425204 1005388 425210 1005400
rect 467926 1005388 467932 1005400
rect 467984 1005388 467990 1005440
rect 209222 1005320 209228 1005372
rect 209280 1005360 209286 1005372
rect 227714 1005360 227720 1005372
rect 209280 1005332 227720 1005360
rect 209280 1005320 209286 1005332
rect 227714 1005320 227720 1005332
rect 227772 1005320 227778 1005372
rect 253290 1005320 253296 1005372
rect 253348 1005360 253354 1005372
rect 280062 1005360 280068 1005372
rect 253348 1005332 280068 1005360
rect 253348 1005320 253354 1005332
rect 280062 1005320 280068 1005332
rect 280120 1005320 280126 1005372
rect 361022 1005320 361028 1005372
rect 361080 1005360 361086 1005372
rect 377950 1005360 377956 1005372
rect 361080 1005332 377956 1005360
rect 361080 1005320 361086 1005332
rect 377950 1005320 377956 1005332
rect 378008 1005320 378014 1005372
rect 428366 1005320 428372 1005372
rect 428424 1005360 428430 1005372
rect 453942 1005360 453948 1005372
rect 428424 1005332 453948 1005360
rect 428424 1005320 428430 1005332
rect 453942 1005320 453948 1005332
rect 454000 1005320 454006 1005372
rect 505830 1005320 505836 1005372
rect 505888 1005360 505894 1005372
rect 517054 1005360 517060 1005372
rect 505888 1005332 517060 1005360
rect 505888 1005320 505894 1005332
rect 517054 1005320 517060 1005332
rect 517112 1005320 517118 1005372
rect 92658 1005252 92664 1005304
rect 92716 1005292 92722 1005304
rect 109310 1005292 109316 1005304
rect 92716 1005264 109316 1005292
rect 92716 1005252 92722 1005264
rect 109310 1005252 109316 1005264
rect 109368 1005252 109374 1005304
rect 259822 1005252 259828 1005304
rect 259880 1005292 259886 1005304
rect 280246 1005292 280252 1005304
rect 259880 1005264 280252 1005292
rect 259880 1005252 259886 1005264
rect 280246 1005252 280252 1005264
rect 280304 1005252 280310 1005304
rect 106458 1005184 106464 1005236
rect 106516 1005224 106522 1005236
rect 125778 1005224 125784 1005236
rect 106516 1005196 125784 1005224
rect 106516 1005184 106522 1005196
rect 125778 1005184 125784 1005196
rect 125836 1005184 125842 1005236
rect 260190 1005184 260196 1005236
rect 260248 1005224 260254 1005236
rect 265066 1005224 265072 1005236
rect 260248 1005196 265072 1005224
rect 260248 1005184 260254 1005196
rect 265066 1005184 265072 1005196
rect 265124 1005184 265130 1005236
rect 360194 1005184 360200 1005236
rect 360252 1005224 360258 1005236
rect 380802 1005224 380808 1005236
rect 360252 1005196 380808 1005224
rect 360252 1005184 360258 1005196
rect 380802 1005184 380808 1005196
rect 380860 1005184 380866 1005236
rect 105630 1005116 105636 1005168
rect 105688 1005156 105694 1005168
rect 125594 1005156 125600 1005168
rect 105688 1005128 125600 1005156
rect 105688 1005116 105694 1005128
rect 125594 1005116 125600 1005128
rect 125652 1005116 125658 1005168
rect 195330 1005116 195336 1005168
rect 195388 1005156 195394 1005168
rect 209590 1005156 209596 1005168
rect 195388 1005128 209596 1005156
rect 195388 1005116 195394 1005128
rect 209590 1005116 209596 1005128
rect 209648 1005116 209654 1005168
rect 210878 1005116 210884 1005168
rect 210936 1005156 210942 1005168
rect 227898 1005156 227904 1005168
rect 210936 1005128 227904 1005156
rect 210936 1005116 210942 1005128
rect 227898 1005116 227904 1005128
rect 227956 1005116 227962 1005168
rect 263042 1005116 263048 1005168
rect 263100 1005156 263106 1005168
rect 264330 1005156 264336 1005168
rect 263100 1005128 264336 1005156
rect 263100 1005116 263106 1005128
rect 264330 1005116 264336 1005128
rect 264388 1005116 264394 1005168
rect 427538 1005116 427544 1005168
rect 427596 1005156 427602 1005168
rect 460842 1005156 460848 1005168
rect 427596 1005128 460848 1005156
rect 427596 1005116 427602 1005128
rect 460842 1005116 460848 1005128
rect 460900 1005116 460906 1005168
rect 201494 1005048 201500 1005100
rect 201552 1005088 201558 1005100
rect 202322 1005088 202328 1005100
rect 201552 1005060 202328 1005088
rect 201552 1005048 201558 1005060
rect 202322 1005048 202328 1005060
rect 202380 1005088 202386 1005100
rect 227622 1005088 227628 1005100
rect 202380 1005060 227628 1005088
rect 202380 1005048 202386 1005060
rect 227622 1005048 227628 1005060
rect 227680 1005048 227686 1005100
rect 261018 1005048 261024 1005100
rect 261076 1005088 261082 1005100
rect 265250 1005088 265256 1005100
rect 261076 1005060 265256 1005088
rect 261076 1005048 261082 1005060
rect 265250 1005048 265256 1005060
rect 265308 1005048 265314 1005100
rect 428826 1005048 428832 1005100
rect 428884 1005088 428890 1005100
rect 465258 1005088 465264 1005100
rect 428884 1005060 465264 1005088
rect 428884 1005048 428890 1005060
rect 465258 1005048 465264 1005060
rect 465316 1005048 465322 1005100
rect 502518 1005048 502524 1005100
rect 502576 1005088 502582 1005100
rect 523218 1005088 523224 1005100
rect 502576 1005060 523224 1005088
rect 502576 1005048 502582 1005060
rect 523218 1005048 523224 1005060
rect 523276 1005048 523282 1005100
rect 150894 1004980 150900 1005032
rect 150952 1005020 150958 1005032
rect 175182 1005020 175188 1005032
rect 150952 1004992 175188 1005020
rect 150952 1004980 150958 1004992
rect 175182 1004980 175188 1004992
rect 175240 1004980 175246 1005032
rect 252830 1004980 252836 1005032
rect 252888 1005020 252894 1005032
rect 253290 1005020 253296 1005032
rect 252888 1004992 253296 1005020
rect 252888 1004980 252894 1004992
rect 253290 1004980 253296 1004992
rect 253348 1004980 253354 1005032
rect 260650 1004980 260656 1005032
rect 260708 1005020 260714 1005032
rect 260708 1004992 264974 1005020
rect 260708 1004980 260714 1004992
rect 157794 1004912 157800 1004964
rect 157852 1004952 157858 1004964
rect 174078 1004952 174084 1004964
rect 157852 1004924 174084 1004952
rect 157852 1004912 157858 1004924
rect 174078 1004912 174084 1004924
rect 174136 1004912 174142 1004964
rect 208394 1004912 208400 1004964
rect 208452 1004952 208458 1004964
rect 227806 1004952 227812 1004964
rect 208452 1004924 227812 1004952
rect 208452 1004912 208458 1004924
rect 227806 1004912 227812 1004924
rect 227864 1004912 227870 1004964
rect 262674 1004912 262680 1004964
rect 262732 1004952 262738 1004964
rect 264330 1004952 264336 1004964
rect 262732 1004924 264336 1004952
rect 262732 1004912 262738 1004924
rect 264330 1004912 264336 1004924
rect 264388 1004912 264394 1004964
rect 264946 1004952 264974 1004992
rect 358170 1004980 358176 1005032
rect 358228 1005020 358234 1005032
rect 383286 1005020 383292 1005032
rect 358228 1004992 383292 1005020
rect 358228 1004980 358234 1004992
rect 383286 1004980 383292 1004992
rect 383344 1004980 383350 1005032
rect 426802 1004980 426808 1005032
rect 426860 1005020 426866 1005032
rect 455598 1005020 455604 1005032
rect 426860 1004992 455604 1005020
rect 426860 1004980 426866 1004992
rect 455598 1004980 455604 1004992
rect 455656 1004980 455662 1005032
rect 504174 1004980 504180 1005032
rect 504232 1005020 504238 1005032
rect 519078 1005020 519084 1005032
rect 504232 1004992 519084 1005020
rect 504232 1004980 504238 1004992
rect 519078 1004980 519084 1004992
rect 519136 1004980 519142 1005032
rect 280154 1004952 280160 1004964
rect 264946 1004924 280160 1004952
rect 280154 1004912 280160 1004924
rect 280212 1004912 280218 1004964
rect 425514 1004912 425520 1004964
rect 425572 1004952 425578 1004964
rect 455414 1004952 455420 1004964
rect 425572 1004924 455420 1004952
rect 425572 1004912 425578 1004924
rect 455414 1004912 455420 1004924
rect 455472 1004912 455478 1004964
rect 552750 1004912 552756 1004964
rect 552808 1004952 552814 1004964
rect 568574 1004952 568580 1004964
rect 552808 1004924 568580 1004952
rect 552808 1004912 552814 1004924
rect 568574 1004912 568580 1004924
rect 568632 1004912 568638 1004964
rect 108022 1004844 108028 1004896
rect 108080 1004884 108086 1004896
rect 109678 1004884 109684 1004896
rect 108080 1004856 109684 1004884
rect 108080 1004844 108086 1004856
rect 109678 1004844 109684 1004856
rect 109736 1004844 109742 1004896
rect 261846 1004844 261852 1004896
rect 261904 1004884 261910 1004896
rect 266262 1004884 266268 1004896
rect 261904 1004856 266268 1004884
rect 261904 1004844 261910 1004856
rect 266262 1004844 266268 1004856
rect 266320 1004844 266326 1004896
rect 427170 1004844 427176 1004896
rect 427228 1004884 427234 1004896
rect 455506 1004884 455512 1004896
rect 427228 1004856 455512 1004884
rect 427228 1004844 427234 1004856
rect 455506 1004844 455512 1004856
rect 455564 1004844 455570 1004896
rect 114646 1004776 114652 1004828
rect 114704 1004816 114710 1004828
rect 125686 1004816 125692 1004828
rect 114704 1004788 125692 1004816
rect 114704 1004776 114710 1004788
rect 125686 1004776 125692 1004788
rect 125744 1004776 125750 1004828
rect 156966 1004776 156972 1004828
rect 157024 1004816 157030 1004828
rect 173986 1004816 173992 1004828
rect 157024 1004788 173992 1004816
rect 157024 1004776 157030 1004788
rect 173986 1004776 173992 1004788
rect 174044 1004776 174050 1004828
rect 423490 1004776 423496 1004828
rect 423548 1004816 423554 1004828
rect 467742 1004816 467748 1004828
rect 423548 1004788 467748 1004816
rect 423548 1004776 423554 1004788
rect 467742 1004776 467748 1004788
rect 467800 1004776 467806 1004828
rect 553118 1004776 553124 1004828
rect 553176 1004816 553182 1004828
rect 557442 1004816 557448 1004828
rect 553176 1004788 557448 1004816
rect 553176 1004776 553182 1004788
rect 557442 1004776 557448 1004788
rect 557500 1004776 557506 1004828
rect 99466 1004708 99472 1004760
rect 99524 1004748 99530 1004760
rect 99524 1004720 121454 1004748
rect 99524 1004708 99530 1004720
rect 92934 1004640 92940 1004692
rect 92992 1004680 92998 1004692
rect 108850 1004680 108856 1004692
rect 92992 1004652 108856 1004680
rect 92992 1004640 92998 1004652
rect 108850 1004640 108856 1004652
rect 108908 1004640 108914 1004692
rect 121426 1004680 121454 1004720
rect 154482 1004708 154488 1004760
rect 154540 1004748 154546 1004760
rect 154540 1004720 155080 1004748
rect 154540 1004708 154546 1004720
rect 125502 1004680 125508 1004692
rect 121426 1004652 125508 1004680
rect 125502 1004640 125508 1004652
rect 125560 1004640 125566 1004692
rect 146018 1004640 146024 1004692
rect 146076 1004680 146082 1004692
rect 154942 1004680 154948 1004692
rect 146076 1004652 154948 1004680
rect 146076 1004640 146082 1004652
rect 154942 1004640 154948 1004652
rect 155000 1004640 155006 1004692
rect 155052 1004680 155080 1004720
rect 159450 1004708 159456 1004760
rect 159508 1004748 159514 1004760
rect 173894 1004748 173900 1004760
rect 159508 1004720 173900 1004748
rect 159508 1004708 159514 1004720
rect 173894 1004708 173900 1004720
rect 173952 1004708 173958 1004760
rect 195974 1004708 195980 1004760
rect 196032 1004748 196038 1004760
rect 206370 1004748 206376 1004760
rect 196032 1004720 206376 1004748
rect 196032 1004708 196038 1004720
rect 206370 1004708 206376 1004720
rect 206428 1004708 206434 1004760
rect 262214 1004708 262220 1004760
rect 262272 1004748 262278 1004760
rect 280338 1004748 280344 1004760
rect 262272 1004720 280344 1004748
rect 262272 1004708 262278 1004720
rect 280338 1004708 280344 1004720
rect 280396 1004708 280402 1004760
rect 358538 1004708 358544 1004760
rect 358596 1004748 358602 1004760
rect 358596 1004720 372614 1004748
rect 358596 1004708 358602 1004720
rect 160646 1004680 160652 1004692
rect 155052 1004652 160652 1004680
rect 160646 1004640 160652 1004652
rect 160704 1004640 160710 1004692
rect 195698 1004640 195704 1004692
rect 195756 1004680 195762 1004692
rect 205174 1004680 205180 1004692
rect 195756 1004652 205180 1004680
rect 195756 1004640 195762 1004652
rect 205174 1004640 205180 1004652
rect 205232 1004640 205238 1004692
rect 261478 1004640 261484 1004692
rect 261536 1004680 261542 1004692
rect 265158 1004680 265164 1004692
rect 261536 1004652 265164 1004680
rect 261536 1004640 261542 1004652
rect 265158 1004640 265164 1004652
rect 265216 1004640 265222 1004692
rect 315114 1004640 315120 1004692
rect 315172 1004680 315178 1004692
rect 331214 1004680 331220 1004692
rect 315172 1004652 331220 1004680
rect 315172 1004640 315178 1004652
rect 331214 1004640 331220 1004652
rect 331272 1004640 331278 1004692
rect 359734 1004640 359740 1004692
rect 359792 1004680 359798 1004692
rect 369854 1004680 369860 1004692
rect 359792 1004652 369860 1004680
rect 359792 1004640 359798 1004652
rect 369854 1004640 369860 1004652
rect 369912 1004640 369918 1004692
rect 372586 1004680 372614 1004720
rect 424686 1004708 424692 1004760
rect 424744 1004748 424750 1004760
rect 467834 1004748 467840 1004760
rect 424744 1004720 467840 1004748
rect 424744 1004708 424750 1004720
rect 467834 1004708 467840 1004720
rect 467892 1004708 467898 1004760
rect 501690 1004708 501696 1004760
rect 501748 1004748 501754 1004760
rect 509142 1004748 509148 1004760
rect 501748 1004720 509148 1004748
rect 501748 1004708 501754 1004720
rect 509142 1004708 509148 1004720
rect 509200 1004708 509206 1004760
rect 551922 1004708 551928 1004760
rect 551980 1004748 551986 1004760
rect 558730 1004748 558736 1004760
rect 551980 1004720 558736 1004748
rect 551980 1004708 551986 1004720
rect 558730 1004708 558736 1004720
rect 558788 1004708 558794 1004760
rect 381722 1004680 381728 1004692
rect 372586 1004652 381728 1004680
rect 381722 1004640 381728 1004652
rect 381780 1004640 381786 1004692
rect 419442 1004640 419448 1004692
rect 419500 1004680 419506 1004692
rect 422294 1004680 422300 1004692
rect 419500 1004652 422300 1004680
rect 419500 1004640 419506 1004652
rect 422294 1004640 422300 1004652
rect 422352 1004640 422358 1004692
rect 458910 1004640 458916 1004692
rect 458968 1004680 458974 1004692
rect 472342 1004680 472348 1004692
rect 458968 1004652 472348 1004680
rect 458968 1004640 458974 1004652
rect 472342 1004640 472348 1004652
rect 472400 1004640 472406 1004692
rect 496722 1004640 496728 1004692
rect 496780 1004680 496786 1004692
rect 499298 1004680 499304 1004692
rect 496780 1004652 499304 1004680
rect 496780 1004640 496786 1004652
rect 499298 1004640 499304 1004652
rect 499356 1004640 499362 1004692
rect 502150 1004640 502156 1004692
rect 502208 1004680 502214 1004692
rect 509234 1004680 509240 1004692
rect 502208 1004652 509240 1004680
rect 502208 1004640 502214 1004652
rect 509234 1004640 509240 1004652
rect 509292 1004640 509298 1004692
rect 554314 1004640 554320 1004692
rect 554372 1004680 554378 1004692
rect 554372 1004652 557488 1004680
rect 554372 1004640 554378 1004652
rect 195146 1004572 195152 1004624
rect 195204 1004612 195210 1004624
rect 205910 1004612 205916 1004624
rect 195204 1004584 205916 1004612
rect 195204 1004572 195210 1004584
rect 205910 1004572 205916 1004584
rect 205968 1004572 205974 1004624
rect 517422 1004572 517428 1004624
rect 517480 1004612 517486 1004624
rect 523954 1004612 523960 1004624
rect 517480 1004584 523960 1004612
rect 517480 1004572 517486 1004584
rect 523954 1004572 523960 1004584
rect 524012 1004572 524018 1004624
rect 557460 1004612 557488 1004652
rect 561306 1004640 561312 1004692
rect 561364 1004680 561370 1004692
rect 567470 1004680 567476 1004692
rect 561364 1004652 567476 1004680
rect 561364 1004640 561370 1004652
rect 567470 1004640 567476 1004652
rect 567528 1004640 567534 1004692
rect 571334 1004612 571340 1004624
rect 557460 1004584 571340 1004612
rect 571334 1004572 571340 1004584
rect 571392 1004572 571398 1004624
rect 557442 1004096 557448 1004148
rect 557500 1004136 557506 1004148
rect 570138 1004136 570144 1004148
rect 557500 1004108 570144 1004136
rect 557500 1004096 557506 1004108
rect 570138 1004096 570144 1004108
rect 570196 1004096 570202 1004148
rect 553946 1003892 553952 1003944
rect 554004 1003932 554010 1003944
rect 571426 1003932 571432 1003944
rect 554004 1003904 571432 1003932
rect 554004 1003892 554010 1003904
rect 571426 1003892 571432 1003904
rect 571484 1003892 571490 1003944
rect 455414 1003348 455420 1003400
rect 455472 1003388 455478 1003400
rect 464246 1003388 464252 1003400
rect 455472 1003360 464252 1003388
rect 455472 1003348 455478 1003360
rect 464246 1003348 464252 1003360
rect 464304 1003348 464310 1003400
rect 455506 1003280 455512 1003332
rect 455564 1003320 455570 1003332
rect 469122 1003320 469128 1003332
rect 455564 1003292 469128 1003320
rect 455564 1003280 455570 1003292
rect 469122 1003280 469128 1003292
rect 469180 1003280 469186 1003332
rect 555510 1003280 555516 1003332
rect 555568 1003320 555574 1003332
rect 574002 1003320 574008 1003332
rect 555568 1003292 574008 1003320
rect 555568 1003280 555574 1003292
rect 574002 1003280 574008 1003292
rect 574060 1003280 574066 1003332
rect 455598 1003212 455604 1003264
rect 455656 1003252 455662 1003264
rect 466454 1003252 466460 1003264
rect 455656 1003224 466460 1003252
rect 455656 1003212 455662 1003224
rect 466454 1003212 466460 1003224
rect 466512 1003212 466518 1003264
rect 554774 1003212 554780 1003264
rect 554832 1003252 554838 1003264
rect 569954 1003252 569960 1003264
rect 554832 1003224 569960 1003252
rect 554832 1003212 554838 1003224
rect 569954 1003212 569960 1003224
rect 570012 1003212 570018 1003264
rect 440418 1001988 440424 1002040
rect 440476 1002028 440482 1002040
rect 440476 1002000 444512 1002028
rect 440476 1001988 440482 1002000
rect 440234 1001920 440240 1001972
rect 440292 1001960 440298 1001972
rect 444484 1001960 444512 1002000
rect 440292 1001932 444420 1001960
rect 444484 1001932 447272 1001960
rect 440292 1001920 440298 1001932
rect 444392 1001892 444420 1001932
rect 447134 1001892 447140 1001904
rect 444392 1001864 447140 1001892
rect 447134 1001852 447140 1001864
rect 447192 1001852 447198 1001904
rect 447244 1001892 447272 1001932
rect 447318 1001892 447324 1001904
rect 447244 1001864 447324 1001892
rect 447318 1001852 447324 1001864
rect 447376 1001852 447382 1001904
rect 466454 1001852 466460 1001904
rect 466512 1001892 466518 1001904
rect 469766 1001892 469772 1001904
rect 466512 1001864 469772 1001892
rect 466512 1001852 466518 1001864
rect 469766 1001852 469772 1001864
rect 469824 1001852 469830 1001904
rect 517054 1001852 517060 1001904
rect 517112 1001892 517118 1001904
rect 519538 1001892 519544 1001904
rect 517112 1001864 519544 1001892
rect 517112 1001852 517118 1001864
rect 519538 1001852 519544 1001864
rect 519596 1001852 519602 1001904
rect 519722 1001852 519728 1001904
rect 519780 1001892 519786 1001904
rect 523862 1001892 523868 1001904
rect 519780 1001864 523868 1001892
rect 519780 1001852 519786 1001864
rect 523862 1001852 523868 1001864
rect 523920 1001852 523926 1001904
rect 558730 1001852 558736 1001904
rect 558788 1001892 558794 1001904
rect 569862 1001892 569868 1001904
rect 558788 1001864 569868 1001892
rect 558788 1001852 558794 1001864
rect 569862 1001852 569868 1001864
rect 569920 1001852 569926 1001904
rect 568574 1001784 568580 1001836
rect 568632 1001824 568638 1001836
rect 572622 1001824 572628 1001836
rect 568632 1001796 572628 1001824
rect 568632 1001784 568638 1001796
rect 572622 1001784 572628 1001796
rect 572680 1001784 572686 1001836
rect 464246 1001716 464252 1001768
rect 464304 1001756 464310 1001768
rect 471698 1001756 471704 1001768
rect 464304 1001728 471704 1001756
rect 464304 1001716 464310 1001728
rect 471698 1001716 471704 1001728
rect 471756 1001716 471762 1001768
rect 376662 1001104 376668 1001156
rect 376720 1001144 376726 1001156
rect 378318 1001144 378324 1001156
rect 376720 1001116 378324 1001144
rect 376720 1001104 376726 1001116
rect 378318 1001104 378324 1001116
rect 378376 1001104 378382 1001156
rect 373166 1001036 373172 1001088
rect 373224 1001076 373230 1001088
rect 381262 1001076 381268 1001088
rect 373224 1001048 381268 1001076
rect 373224 1001036 373230 1001048
rect 381262 1001036 381268 1001048
rect 381320 1001036 381326 1001088
rect 360562 1000696 360568 1000748
rect 360620 1000736 360626 1000748
rect 383562 1000736 383568 1000748
rect 360620 1000708 383568 1000736
rect 360620 1000696 360626 1000708
rect 383562 1000696 383568 1000708
rect 383620 1000696 383626 1000748
rect 361390 1000628 361396 1000680
rect 361448 1000668 361454 1000680
rect 383378 1000668 383384 1000680
rect 361448 1000640 383384 1000668
rect 361448 1000628 361454 1000640
rect 383378 1000628 383384 1000640
rect 383436 1000628 383442 1000680
rect 369854 1000560 369860 1000612
rect 369912 1000600 369918 1000612
rect 383470 1000600 383476 1000612
rect 369912 1000572 383476 1000600
rect 369912 1000560 369918 1000572
rect 383470 1000560 383476 1000572
rect 383528 1000560 383534 1000612
rect 427998 1000560 428004 1000612
rect 428056 1000600 428062 1000612
rect 472618 1000600 472624 1000612
rect 428056 1000572 472624 1000600
rect 428056 1000560 428062 1000572
rect 472618 1000560 472624 1000572
rect 472676 1000560 472682 1000612
rect 358906 1000492 358912 1000544
rect 358964 1000532 358970 1000544
rect 383562 1000532 383568 1000544
rect 358964 1000504 383568 1000532
rect 358964 1000492 358970 1000504
rect 383562 1000492 383568 1000504
rect 383620 1000492 383626 1000544
rect 426342 1000492 426348 1000544
rect 426400 1000532 426406 1000544
rect 472526 1000532 472532 1000544
rect 426400 1000504 472532 1000532
rect 426400 1000492 426406 1000504
rect 472526 1000492 472532 1000504
rect 472584 1000492 472590 1000544
rect 380894 1000288 380900 1000340
rect 380952 1000328 380958 1000340
rect 383562 1000328 383568 1000340
rect 380952 1000300 383568 1000328
rect 380952 1000288 380958 1000300
rect 383562 1000288 383568 1000300
rect 383620 1000288 383626 1000340
rect 566550 1000056 566556 1000068
rect 546466 1000028 566556 1000056
rect 503346 999948 503352 1000000
rect 503404 999988 503410 1000000
rect 516042 999988 516048 1000000
rect 503404 999960 516048 999988
rect 503404 999948 503410 999960
rect 516042 999948 516048 999960
rect 516100 999948 516106 1000000
rect 92566 999880 92572 999932
rect 92624 999920 92630 999932
rect 116026 999920 116032 999932
rect 92624 999892 116032 999920
rect 92624 999880 92630 999892
rect 116026 999880 116032 999892
rect 116084 999880 116090 999932
rect 246758 999880 246764 999932
rect 246816 999920 246822 999932
rect 258626 999920 258632 999932
rect 246816 999892 258632 999920
rect 246816 999880 246822 999892
rect 258626 999880 258632 999892
rect 258684 999880 258690 999932
rect 92474 999812 92480 999864
rect 92532 999852 92538 999864
rect 104342 999852 104348 999864
rect 92532 999824 104348 999852
rect 92532 999812 92538 999824
rect 104342 999812 104348 999824
rect 104400 999812 104406 999864
rect 246574 999812 246580 999864
rect 246632 999852 246638 999864
rect 257338 999852 257344 999864
rect 246632 999824 257344 999852
rect 246632 999812 246638 999824
rect 257338 999812 257344 999824
rect 257396 999812 257402 999864
rect 312170 999812 312176 999864
rect 312228 999852 312234 999864
rect 318886 999852 318892 999864
rect 312228 999824 318892 999852
rect 312228 999812 312234 999824
rect 318886 999812 318892 999824
rect 318944 999812 318950 999864
rect 434622 999852 434628 999864
rect 400186 999824 434628 999852
rect 92290 999744 92296 999796
rect 92348 999784 92354 999796
rect 102778 999784 102784 999796
rect 92348 999756 102784 999784
rect 92348 999744 92354 999756
rect 102778 999744 102784 999756
rect 102836 999744 102842 999796
rect 246666 999744 246672 999796
rect 246724 999784 246730 999796
rect 256970 999784 256976 999796
rect 246724 999756 256976 999784
rect 246724 999744 246730 999756
rect 256970 999744 256976 999756
rect 257028 999744 257034 999796
rect 311434 999744 311440 999796
rect 311492 999784 311498 999796
rect 315942 999784 315948 999796
rect 311492 999756 315948 999784
rect 311492 999744 311498 999756
rect 315942 999744 315948 999756
rect 316000 999744 316006 999796
rect 246942 999676 246948 999728
rect 247000 999716 247006 999728
rect 257798 999716 257804 999728
rect 247000 999688 257804 999716
rect 247000 999676 247006 999688
rect 257798 999676 257804 999688
rect 257856 999676 257862 999728
rect 313826 999676 313832 999728
rect 313884 999716 313890 999728
rect 318702 999716 318708 999728
rect 313884 999688 318708 999716
rect 313884 999676 313890 999688
rect 318702 999676 318708 999688
rect 318760 999676 318766 999728
rect 92382 999608 92388 999660
rect 92440 999648 92446 999660
rect 102318 999648 102324 999660
rect 92440 999620 102324 999648
rect 92440 999608 92446 999620
rect 102318 999608 102324 999620
rect 102376 999608 102382 999660
rect 195238 999608 195244 999660
rect 195296 999648 195302 999660
rect 205542 999648 205548 999660
rect 195296 999620 205548 999648
rect 195296 999608 195302 999620
rect 205542 999608 205548 999620
rect 205600 999608 205606 999660
rect 310146 999608 310152 999660
rect 310204 999648 310210 999660
rect 314930 999648 314936 999660
rect 310204 999620 314936 999648
rect 310204 999608 310210 999620
rect 314930 999608 314936 999620
rect 314988 999608 314994 999660
rect 155770 999540 155776 999592
rect 155828 999580 155834 999592
rect 160278 999580 160284 999592
rect 155828 999552 160284 999580
rect 155828 999540 155834 999552
rect 160278 999540 160284 999552
rect 160336 999540 160342 999592
rect 195606 999540 195612 999592
rect 195664 999580 195670 999592
rect 203518 999580 203524 999592
rect 195664 999552 203524 999580
rect 195664 999540 195670 999552
rect 203518 999540 203524 999552
rect 203576 999540 203582 999592
rect 312998 999540 313004 999592
rect 313056 999580 313062 999592
rect 317598 999580 317604 999592
rect 313056 999552 317604 999580
rect 313056 999540 313062 999552
rect 317598 999540 317604 999552
rect 317656 999540 317662 999592
rect 92750 999472 92756 999524
rect 92808 999512 92814 999524
rect 101950 999512 101956 999524
rect 92808 999484 101956 999512
rect 92808 999472 92814 999484
rect 101950 999472 101956 999484
rect 102008 999472 102014 999524
rect 159082 999472 159088 999524
rect 159140 999512 159146 999524
rect 162854 999512 162860 999524
rect 159140 999484 162860 999512
rect 159140 999472 159146 999484
rect 162854 999472 162860 999484
rect 162912 999472 162918 999524
rect 195422 999472 195428 999524
rect 195480 999512 195486 999524
rect 203886 999512 203892 999524
rect 195480 999484 203892 999512
rect 195480 999472 195486 999484
rect 203886 999472 203892 999484
rect 203944 999472 203950 999524
rect 314654 999472 314660 999524
rect 314712 999512 314718 999524
rect 319070 999512 319076 999524
rect 314712 999484 319076 999512
rect 314712 999472 314718 999484
rect 319070 999472 319076 999484
rect 319128 999472 319134 999524
rect 99282 999404 99288 999456
rect 99340 999444 99346 999456
rect 103146 999444 103152 999456
rect 99340 999416 103152 999444
rect 99340 999404 99346 999416
rect 103146 999404 103152 999416
rect 103204 999404 103210 999456
rect 195514 999404 195520 999456
rect 195572 999444 195578 999456
rect 202322 999444 202328 999456
rect 195572 999416 202328 999444
rect 195572 999404 195578 999416
rect 202322 999404 202328 999416
rect 202380 999404 202386 999456
rect 309778 999404 309784 999456
rect 309836 999444 309842 999456
rect 314838 999444 314844 999456
rect 309836 999416 314844 999444
rect 309836 999404 309842 999416
rect 314838 999404 314844 999416
rect 314896 999404 314902 999456
rect 198366 999336 198372 999388
rect 198424 999376 198430 999388
rect 204714 999376 204720 999388
rect 198424 999348 204720 999376
rect 198424 999336 198430 999348
rect 204714 999336 204720 999348
rect 204772 999336 204778 999388
rect 312630 999336 312636 999388
rect 312688 999376 312694 999388
rect 317414 999376 317420 999388
rect 312688 999348 317420 999376
rect 312688 999336 312694 999348
rect 317414 999336 317420 999348
rect 317472 999336 317478 999388
rect 198458 999268 198464 999320
rect 198516 999308 198522 999320
rect 204346 999308 204352 999320
rect 198516 999280 204352 999308
rect 198516 999268 198522 999280
rect 204346 999268 204352 999280
rect 204404 999268 204410 999320
rect 310974 999268 310980 999320
rect 311032 999308 311038 999320
rect 315022 999308 315028 999320
rect 311032 999280 315028 999308
rect 311032 999268 311038 999280
rect 315022 999268 315028 999280
rect 315080 999268 315086 999320
rect 198642 999200 198648 999252
rect 198700 999240 198706 999252
rect 202690 999240 202696 999252
rect 198700 999212 202696 999240
rect 198700 999200 198706 999212
rect 202690 999200 202696 999212
rect 202748 999200 202754 999252
rect 253842 999200 253848 999252
rect 253900 999240 253906 999252
rect 256510 999240 256516 999252
rect 253900 999212 256516 999240
rect 253900 999200 253906 999212
rect 256510 999200 256516 999212
rect 256568 999200 256574 999252
rect 311802 999200 311808 999252
rect 311860 999240 311866 999252
rect 315114 999240 315120 999252
rect 311860 999212 315120 999240
rect 311860 999200 311866 999212
rect 315114 999200 315120 999212
rect 315172 999200 315178 999252
rect 357342 999200 357348 999252
rect 357400 999240 357406 999252
rect 364886 999240 364892 999252
rect 357400 999212 364892 999240
rect 357400 999200 357406 999212
rect 364886 999200 364892 999212
rect 364944 999200 364950 999252
rect 198550 999132 198556 999184
rect 198608 999172 198614 999184
rect 203058 999172 203064 999184
rect 198608 999144 203064 999172
rect 198608 999132 198614 999144
rect 203058 999132 203064 999144
rect 203116 999132 203122 999184
rect 258534 999132 258540 999184
rect 258592 999172 258598 999184
rect 262214 999172 262220 999184
rect 258592 999144 262220 999172
rect 258592 999132 258598 999144
rect 262214 999132 262220 999144
rect 262272 999132 262278 999184
rect 314286 999132 314292 999184
rect 314344 999172 314350 999184
rect 317506 999172 317512 999184
rect 314344 999144 317512 999172
rect 314344 999132 314350 999144
rect 317506 999132 317512 999144
rect 317564 999132 317570 999184
rect 357710 999132 357716 999184
rect 357768 999172 357774 999184
rect 365070 999172 365076 999184
rect 357768 999144 365076 999172
rect 357768 999132 357774 999144
rect 365070 999132 365076 999144
rect 365128 999132 365134 999184
rect 378042 999132 378048 999184
rect 378100 999172 378106 999184
rect 383194 999172 383200 999184
rect 378100 999144 383200 999172
rect 378100 999132 378106 999144
rect 383194 999132 383200 999144
rect 383252 999132 383258 999184
rect 400030 999132 400036 999184
rect 400088 999172 400094 999184
rect 400186 999172 400214 999824
rect 434622 999812 434628 999824
rect 434680 999812 434686 999864
rect 430850 999744 430856 999796
rect 430908 999784 430914 999796
rect 438118 999784 438124 999796
rect 430908 999756 438124 999784
rect 430908 999744 430914 999756
rect 438118 999744 438124 999756
rect 438176 999744 438182 999796
rect 508682 999744 508688 999796
rect 508740 999784 508746 999796
rect 515214 999784 515220 999796
rect 508740 999756 515220 999784
rect 508740 999744 508746 999756
rect 515214 999744 515220 999756
rect 515272 999744 515278 999796
rect 431678 999676 431684 999728
rect 431736 999716 431742 999728
rect 437934 999716 437940 999728
rect 431736 999688 437940 999716
rect 431736 999676 431742 999688
rect 437934 999676 437940 999688
rect 437992 999676 437998 999728
rect 506198 999676 506204 999728
rect 506256 999716 506262 999728
rect 511902 999716 511908 999728
rect 506256 999688 511908 999716
rect 506256 999676 506262 999688
rect 511902 999676 511908 999688
rect 511960 999676 511966 999728
rect 429194 999608 429200 999660
rect 429252 999648 429258 999660
rect 434714 999648 434720 999660
rect 429252 999620 434720 999648
rect 429252 999608 429258 999620
rect 434714 999608 434720 999620
rect 434772 999608 434778 999660
rect 507026 999608 507032 999660
rect 507084 999648 507090 999660
rect 512086 999648 512092 999660
rect 507084 999620 512092 999648
rect 507084 999608 507090 999620
rect 512086 999608 512092 999620
rect 512144 999608 512150 999660
rect 430022 999540 430028 999592
rect 430080 999580 430086 999592
rect 434806 999580 434812 999592
rect 430080 999552 434812 999580
rect 430080 999540 430086 999552
rect 434806 999540 434812 999552
rect 434864 999540 434870 999592
rect 508222 999540 508228 999592
rect 508280 999580 508286 999592
rect 513466 999580 513472 999592
rect 508280 999552 513472 999580
rect 508280 999540 508286 999552
rect 513466 999540 513472 999552
rect 513524 999540 513530 999592
rect 431218 999472 431224 999524
rect 431276 999512 431282 999524
rect 436186 999512 436192 999524
rect 431276 999484 436192 999512
rect 431276 999472 431282 999484
rect 436186 999472 436192 999484
rect 436244 999472 436250 999524
rect 507854 999472 507860 999524
rect 507912 999512 507918 999524
rect 512270 999512 512276 999524
rect 507912 999484 512276 999512
rect 507912 999472 507918 999484
rect 512270 999472 512276 999484
rect 512328 999472 512334 999524
rect 429654 999404 429660 999456
rect 429712 999444 429718 999456
rect 433426 999444 433432 999456
rect 429712 999416 433432 999444
rect 429712 999404 429718 999416
rect 433426 999404 433432 999416
rect 433484 999404 433490 999456
rect 506566 999404 506572 999456
rect 506624 999444 506630 999456
rect 510890 999444 510896 999456
rect 506624 999416 510896 999444
rect 506624 999404 506630 999416
rect 510890 999404 510896 999416
rect 510948 999404 510954 999456
rect 432506 999336 432512 999388
rect 432564 999376 432570 999388
rect 437382 999376 437388 999388
rect 432564 999348 437388 999376
rect 432564 999336 432570 999348
rect 437382 999336 437388 999348
rect 437440 999336 437446 999388
rect 500494 999336 500500 999388
rect 500552 999376 500558 999388
rect 508774 999376 508780 999388
rect 500552 999348 508780 999376
rect 500552 999336 500558 999348
rect 508774 999336 508780 999348
rect 508832 999336 508838 999388
rect 509050 999336 509056 999388
rect 509108 999376 509114 999388
rect 513650 999376 513656 999388
rect 509108 999348 513656 999376
rect 509108 999336 509114 999348
rect 513650 999336 513656 999348
rect 513708 999336 513714 999388
rect 432874 999268 432880 999320
rect 432932 999308 432938 999320
rect 437566 999308 437572 999320
rect 432932 999280 437572 999308
rect 432932 999268 432938 999280
rect 437566 999268 437572 999280
rect 437624 999268 437630 999320
rect 509510 999268 509516 999320
rect 509568 999308 509574 999320
rect 514846 999308 514852 999320
rect 509568 999280 514852 999308
rect 509568 999268 509574 999280
rect 514846 999268 514852 999280
rect 514904 999268 514910 999320
rect 432046 999200 432052 999252
rect 432104 999240 432110 999252
rect 436094 999240 436100 999252
rect 432104 999212 436100 999240
rect 432104 999200 432110 999212
rect 436094 999200 436100 999212
rect 436152 999200 436158 999252
rect 500862 999200 500868 999252
rect 500920 999240 500926 999252
rect 500920 999212 505784 999240
rect 500920 999200 500926 999212
rect 400088 999144 400214 999172
rect 400088 999132 400094 999144
rect 430390 999132 430396 999184
rect 430448 999172 430454 999184
rect 433334 999172 433340 999184
rect 430448 999144 433340 999172
rect 430448 999132 430454 999144
rect 433334 999132 433340 999144
rect 433392 999132 433398 999184
rect 465258 999132 465264 999184
rect 465316 999172 465322 999184
rect 472434 999172 472440 999184
rect 465316 999144 472440 999172
rect 465316 999132 465322 999144
rect 472434 999132 472440 999144
rect 472492 999132 472498 999184
rect 488902 999132 488908 999184
rect 488960 999172 488966 999184
rect 505646 999172 505652 999184
rect 488960 999144 505652 999172
rect 488960 999132 488966 999144
rect 505646 999132 505652 999144
rect 505704 999132 505710 999184
rect 505756 999172 505784 999212
rect 507394 999200 507400 999252
rect 507452 999240 507458 999252
rect 510706 999240 510712 999252
rect 507452 999212 510712 999240
rect 507452 999200 507458 999212
rect 510706 999200 510712 999212
rect 510764 999200 510770 999252
rect 540330 999200 540336 999252
rect 540388 999240 540394 999252
rect 546466 999240 546494 1000028
rect 566550 1000016 566556 1000028
rect 566608 1000016 566614 1000068
rect 560846 999744 560852 999796
rect 560904 999784 560910 999796
rect 567102 999784 567108 999796
rect 560904 999756 567108 999784
rect 560904 999744 560910 999756
rect 567102 999744 567108 999756
rect 567160 999744 567166 999796
rect 560478 999608 560484 999660
rect 560536 999648 560542 999660
rect 565814 999648 565820 999660
rect 560536 999620 565820 999648
rect 560536 999608 560542 999620
rect 565814 999608 565820 999620
rect 565872 999608 565878 999660
rect 590654 999472 590660 999524
rect 590712 999512 590718 999524
rect 625798 999512 625804 999524
rect 590712 999484 625804 999512
rect 590712 999472 590718 999484
rect 625798 999472 625804 999484
rect 625856 999472 625862 999524
rect 610066 999404 610072 999456
rect 610124 999444 610130 999456
rect 625706 999444 625712 999456
rect 610124 999416 625712 999444
rect 610124 999404 610130 999416
rect 625706 999404 625712 999416
rect 625764 999404 625770 999456
rect 609974 999336 609980 999388
rect 610032 999376 610038 999388
rect 625614 999376 625620 999388
rect 610032 999348 625620 999376
rect 610032 999336 610038 999348
rect 625614 999336 625620 999348
rect 625672 999336 625678 999388
rect 601602 999268 601608 999320
rect 601660 999308 601666 999320
rect 625798 999308 625804 999320
rect 601660 999280 625804 999308
rect 601660 999268 601666 999280
rect 625798 999268 625804 999280
rect 625856 999268 625862 999320
rect 540388 999212 546494 999240
rect 540388 999200 540394 999212
rect 593414 999200 593420 999252
rect 593472 999240 593478 999252
rect 625522 999240 625528 999252
rect 593472 999212 625528 999240
rect 593472 999200 593478 999212
rect 625522 999200 625528 999212
rect 625580 999200 625586 999252
rect 509510 999172 509516 999184
rect 505756 999144 509516 999172
rect 509510 999132 509516 999144
rect 509568 999132 509574 999184
rect 509878 999132 509884 999184
rect 509936 999172 509942 999184
rect 514662 999172 514668 999184
rect 509936 999144 514668 999172
rect 509936 999132 509942 999144
rect 514662 999132 514668 999144
rect 514720 999132 514726 999184
rect 552290 999132 552296 999184
rect 552348 999172 552354 999184
rect 558914 999172 558920 999184
rect 552348 999144 558920 999172
rect 552348 999132 552354 999144
rect 558914 999132 558920 999144
rect 558972 999132 558978 999184
rect 144270 999064 144276 999116
rect 144328 999104 144334 999116
rect 158254 999104 158260 999116
rect 144328 999076 158260 999104
rect 144328 999064 144334 999076
rect 158254 999064 158260 999076
rect 158312 999064 158318 999116
rect 246574 999064 246580 999116
rect 246632 999104 246638 999116
rect 265158 999104 265164 999116
rect 246632 999076 265164 999104
rect 246632 999064 246638 999076
rect 265158 999064 265164 999076
rect 265216 999064 265222 999116
rect 298738 999064 298744 999116
rect 298796 999104 298802 999116
rect 317598 999104 317604 999116
rect 298796 999076 317604 999104
rect 298796 999064 298802 999076
rect 317598 999064 317604 999076
rect 317656 999064 317662 999116
rect 399938 999064 399944 999116
rect 399996 999104 400002 999116
rect 436186 999104 436192 999116
rect 399996 999076 436192 999104
rect 399996 999064 400002 999076
rect 436186 999064 436192 999076
rect 436244 999064 436250 999116
rect 453942 999064 453948 999116
rect 454000 999104 454006 999116
rect 462590 999104 462596 999116
rect 454000 999076 462596 999104
rect 454000 999064 454006 999076
rect 462590 999064 462596 999076
rect 462648 999064 462654 999116
rect 489454 999064 489460 999116
rect 489512 999104 489518 999116
rect 513466 999104 513472 999116
rect 489512 999076 513472 999104
rect 489512 999064 489518 999076
rect 513466 999064 513472 999076
rect 513524 999064 513530 999116
rect 508774 998996 508780 999048
rect 508832 999036 508838 999048
rect 521286 999036 521292 999048
rect 508832 999008 521292 999036
rect 508832 998996 508838 999008
rect 521286 998996 521292 999008
rect 521344 998996 521350 999048
rect 509142 998928 509148 998980
rect 509200 998968 509206 998980
rect 521378 998968 521384 998980
rect 509200 998940 521384 998968
rect 509200 998928 509206 998940
rect 521378 998928 521384 998940
rect 521436 998928 521442 998980
rect 509234 998860 509240 998912
rect 509292 998900 509298 998912
rect 520550 998900 520556 998912
rect 509292 998872 520556 998900
rect 509292 998860 509298 998872
rect 520550 998860 520556 998872
rect 520608 998860 520614 998912
rect 509510 998792 509516 998844
rect 509568 998832 509574 998844
rect 521470 998832 521476 998844
rect 509568 998804 521476 998832
rect 509568 998792 509574 998804
rect 521470 998792 521476 998804
rect 521528 998792 521534 998844
rect 364886 998452 364892 998504
rect 364944 998492 364950 998504
rect 374546 998492 374552 998504
rect 364944 998464 374552 998492
rect 364944 998452 364950 998464
rect 374546 998452 374552 998464
rect 374604 998452 374610 998504
rect 467834 998316 467840 998368
rect 467892 998356 467898 998368
rect 469214 998356 469220 998368
rect 467892 998328 469220 998356
rect 467892 998316 467898 998328
rect 469214 998316 469220 998328
rect 469272 998316 469278 998368
rect 467926 998180 467932 998232
rect 467984 998220 467990 998232
rect 471054 998220 471060 998232
rect 467984 998192 471060 998220
rect 467984 998180 467990 998192
rect 471054 998180 471060 998192
rect 471112 998180 471118 998232
rect 518894 998180 518900 998232
rect 518952 998220 518958 998232
rect 521654 998220 521660 998232
rect 518952 998192 521660 998220
rect 518952 998180 518958 998192
rect 521654 998180 521660 998192
rect 521712 998180 521718 998232
rect 467742 998044 467748 998096
rect 467800 998084 467806 998096
rect 469306 998084 469312 998096
rect 467800 998056 469312 998084
rect 467800 998044 467806 998056
rect 469306 998044 469312 998056
rect 469364 998044 469370 998096
rect 558914 997908 558920 997960
rect 558972 997948 558978 997960
rect 568666 997948 568672 997960
rect 558972 997920 568672 997948
rect 558972 997908 558978 997920
rect 568666 997908 568672 997920
rect 568724 997908 568730 997960
rect 365070 997772 365076 997824
rect 365128 997812 365134 997824
rect 374454 997812 374460 997824
rect 365128 997784 374460 997812
rect 365128 997772 365134 997784
rect 374454 997772 374460 997784
rect 374512 997772 374518 997824
rect 143810 997704 143816 997756
rect 143868 997744 143874 997756
rect 156138 997744 156144 997756
rect 143868 997716 156144 997744
rect 143868 997704 143874 997716
rect 156138 997704 156144 997716
rect 156196 997704 156202 997756
rect 501322 997704 501328 997756
rect 501380 997744 501386 997756
rect 521562 997744 521568 997756
rect 501380 997716 521568 997744
rect 501380 997704 501386 997716
rect 521562 997704 521568 997716
rect 521620 997704 521626 997756
rect 553486 997704 553492 997756
rect 553544 997744 553550 997756
rect 568574 997744 568580 997756
rect 553544 997716 568580 997744
rect 553544 997704 553550 997716
rect 568574 997704 568580 997716
rect 568632 997704 568638 997756
rect 569862 997704 569868 997756
rect 569920 997744 569926 997756
rect 623774 997744 623780 997756
rect 569920 997716 623780 997744
rect 569920 997704 569926 997716
rect 623774 997704 623780 997716
rect 623832 997704 623838 997756
rect 556338 997636 556344 997688
rect 556396 997676 556402 997688
rect 601602 997676 601608 997688
rect 556396 997648 601608 997676
rect 556396 997636 556402 997648
rect 601602 997636 601608 997648
rect 601660 997636 601666 997688
rect 571334 997568 571340 997620
rect 571392 997608 571398 997620
rect 609974 997608 609980 997620
rect 571392 997580 609980 997608
rect 571392 997568 571398 997580
rect 609974 997568 609980 997580
rect 610032 997568 610038 997620
rect 569954 997500 569960 997552
rect 570012 997540 570018 997552
rect 610066 997540 610072 997552
rect 570012 997512 610072 997540
rect 570012 997500 570018 997512
rect 610066 997500 610072 997512
rect 610124 997500 610130 997552
rect 557166 997432 557172 997484
rect 557224 997472 557230 997484
rect 620922 997472 620928 997484
rect 557224 997444 620928 997472
rect 557224 997432 557230 997444
rect 620922 997432 620928 997444
rect 620980 997432 620986 997484
rect 571426 997364 571432 997416
rect 571484 997404 571490 997416
rect 590654 997404 590660 997416
rect 571484 997376 590660 997404
rect 571484 997364 571490 997376
rect 590654 997364 590660 997376
rect 590712 997364 590718 997416
rect 572622 997296 572628 997348
rect 572680 997336 572686 997348
rect 593414 997336 593420 997348
rect 572680 997308 593420 997336
rect 572680 997296 572686 997308
rect 593414 997296 593420 997308
rect 593472 997296 593478 997348
rect 107654 997160 107660 997212
rect 107712 997200 107718 997212
rect 115934 997200 115940 997212
rect 107712 997172 115940 997200
rect 107712 997160 107718 997172
rect 115934 997160 115940 997172
rect 115992 997160 115998 997212
rect 210418 997160 210424 997212
rect 210476 997200 210482 997212
rect 215294 997200 215300 997212
rect 210476 997172 215300 997200
rect 210476 997160 210482 997172
rect 215294 997160 215300 997172
rect 215352 997160 215358 997212
rect 363414 997160 363420 997212
rect 363472 997200 363478 997212
rect 367094 997200 367100 997212
rect 363472 997172 367100 997200
rect 363472 997160 363478 997172
rect 367094 997160 367100 997172
rect 367152 997160 367158 997212
rect 96522 996412 96528 996464
rect 96580 996452 96586 996464
rect 101122 996452 101128 996464
rect 96580 996424 101128 996452
rect 96580 996412 96586 996424
rect 101122 996412 101128 996424
rect 101180 996412 101186 996464
rect 148870 996412 148876 996464
rect 148928 996452 148934 996464
rect 154114 996452 154120 996464
rect 148928 996424 154120 996452
rect 148928 996412 148934 996424
rect 154114 996412 154120 996424
rect 154172 996412 154178 996464
rect 146202 996344 146208 996396
rect 146260 996384 146266 996396
rect 151722 996384 151728 996396
rect 146260 996356 151728 996384
rect 146260 996344 146266 996356
rect 151722 996344 151728 996356
rect 151780 996344 151786 996396
rect 301774 996276 301780 996328
rect 301832 996316 301838 996328
rect 308122 996316 308128 996328
rect 301832 996288 308128 996316
rect 301832 996276 301838 996288
rect 308122 996276 308128 996288
rect 308180 996276 308186 996328
rect 146110 996208 146116 996260
rect 146168 996248 146174 996260
rect 153746 996248 153752 996260
rect 146168 996220 153752 996248
rect 146168 996208 146174 996220
rect 153746 996208 153752 996220
rect 153804 996208 153810 996260
rect 211246 996248 211252 996260
rect 198706 996220 211252 996248
rect 125686 996140 125692 996192
rect 125744 996180 125750 996192
rect 159450 996180 159456 996192
rect 125744 996152 159456 996180
rect 125744 996140 125750 996152
rect 159450 996140 159456 996152
rect 159508 996140 159514 996192
rect 173894 996140 173900 996192
rect 173952 996180 173958 996192
rect 198706 996180 198734 996220
rect 211246 996208 211252 996220
rect 211304 996208 211310 996260
rect 300210 996208 300216 996260
rect 300268 996248 300274 996260
rect 308950 996248 308956 996260
rect 300268 996220 308956 996248
rect 300268 996208 300274 996220
rect 308950 996208 308956 996220
rect 309008 996208 309014 996260
rect 365438 996208 365444 996260
rect 365496 996248 365502 996260
rect 371142 996248 371148 996260
rect 365496 996220 371148 996248
rect 365496 996208 365502 996220
rect 371142 996208 371148 996220
rect 371200 996208 371206 996260
rect 208762 996180 208768 996192
rect 173952 996152 198734 996180
rect 204088 996152 208768 996180
rect 173952 996140 173958 996152
rect 96522 996072 96528 996124
rect 96580 996112 96586 996124
rect 100294 996112 100300 996124
rect 96580 996084 100300 996112
rect 96580 996072 96586 996084
rect 100294 996072 100300 996084
rect 100352 996072 100358 996124
rect 108850 996072 108856 996124
rect 108908 996112 108914 996124
rect 113266 996112 113272 996124
rect 108908 996084 113272 996112
rect 108908 996072 108914 996084
rect 113266 996072 113272 996084
rect 113324 996072 113330 996124
rect 125778 996072 125784 996124
rect 125836 996112 125842 996124
rect 157794 996112 157800 996124
rect 125836 996084 157800 996112
rect 125836 996072 125842 996084
rect 157794 996072 157800 996084
rect 157852 996072 157858 996124
rect 173986 996072 173992 996124
rect 174044 996112 174050 996124
rect 204088 996112 204116 996152
rect 208762 996140 208768 996152
rect 208820 996180 208826 996192
rect 212810 996180 212816 996192
rect 208820 996152 212816 996180
rect 208820 996140 208826 996152
rect 212810 996140 212816 996152
rect 212868 996140 212874 996192
rect 227898 996140 227904 996192
rect 227956 996180 227962 996192
rect 267826 996180 267832 996192
rect 227956 996152 267832 996180
rect 227956 996140 227962 996152
rect 267826 996140 267832 996152
rect 267884 996180 267890 996192
rect 270402 996180 270408 996192
rect 267884 996152 270408 996180
rect 267884 996140 267890 996152
rect 270402 996140 270408 996152
rect 270460 996140 270466 996192
rect 280154 996140 280160 996192
rect 280212 996180 280218 996192
rect 317414 996180 317420 996192
rect 280212 996152 317420 996180
rect 280212 996140 280218 996152
rect 317414 996140 317420 996152
rect 317472 996140 317478 996192
rect 364242 996140 364248 996192
rect 364300 996180 364306 996192
rect 367278 996180 367284 996192
rect 364300 996152 367284 996180
rect 364300 996140 364306 996152
rect 367278 996140 367284 996152
rect 367336 996140 367342 996192
rect 512270 996140 512276 996192
rect 512328 996180 512334 996192
rect 559282 996180 559288 996192
rect 512328 996152 559288 996180
rect 512328 996140 512334 996152
rect 559282 996140 559288 996152
rect 559340 996140 559346 996192
rect 174044 996084 204116 996112
rect 174044 996072 174050 996084
rect 204162 996072 204168 996124
rect 204220 996112 204226 996124
rect 211614 996112 211620 996124
rect 204220 996084 211620 996112
rect 204220 996072 204226 996084
rect 211614 996072 211620 996084
rect 211672 996072 211678 996124
rect 227806 996072 227812 996124
rect 227864 996112 227870 996124
rect 265066 996112 265072 996124
rect 227864 996084 265072 996112
rect 227864 996072 227870 996084
rect 265066 996072 265072 996084
rect 265124 996112 265130 996124
rect 267642 996112 267648 996124
rect 265124 996084 267648 996112
rect 265124 996072 265130 996084
rect 267642 996072 267648 996084
rect 267700 996072 267706 996124
rect 280338 996072 280344 996124
rect 280396 996112 280402 996124
rect 317506 996112 317512 996124
rect 280396 996084 317512 996112
rect 280396 996072 280402 996084
rect 317506 996072 317512 996084
rect 317564 996072 317570 996124
rect 364702 996072 364708 996124
rect 364760 996112 364766 996124
rect 369854 996112 369860 996124
rect 364760 996084 369860 996112
rect 364760 996072 364766 996084
rect 369854 996072 369860 996084
rect 369912 996072 369918 996124
rect 558454 996072 558460 996124
rect 558512 996112 558518 996124
rect 564434 996112 564440 996124
rect 558512 996084 564440 996112
rect 558512 996072 558518 996084
rect 564434 996072 564440 996084
rect 564492 996072 564498 996124
rect 96430 996004 96436 996056
rect 96488 996044 96494 996056
rect 101490 996044 101496 996056
rect 96488 996016 101496 996044
rect 96488 996004 96494 996016
rect 101490 996004 101496 996016
rect 101548 996004 101554 996056
rect 108482 996004 108488 996056
rect 108540 996044 108546 996056
rect 113174 996044 113180 996056
rect 108540 996016 113180 996044
rect 108540 996004 108546 996016
rect 113174 996004 113180 996016
rect 113232 996004 113238 996056
rect 125594 996004 125600 996056
rect 125652 996044 125658 996056
rect 156966 996044 156972 996056
rect 125652 996016 156972 996044
rect 125652 996004 125658 996016
rect 156966 996004 156972 996016
rect 157024 996044 157030 996056
rect 160186 996044 160192 996056
rect 157024 996016 160192 996044
rect 157024 996004 157030 996016
rect 160186 996004 160192 996016
rect 160244 996004 160250 996056
rect 174078 996004 174084 996056
rect 174136 996044 174142 996056
rect 209590 996044 209596 996056
rect 174136 996016 209596 996044
rect 174136 996004 174142 996016
rect 209590 996004 209596 996016
rect 209648 996044 209654 996056
rect 212626 996044 212632 996056
rect 209648 996016 212632 996044
rect 209648 996004 209654 996016
rect 212626 996004 212632 996016
rect 212684 996004 212690 996056
rect 227714 996004 227720 996056
rect 227772 996044 227778 996056
rect 265250 996044 265256 996056
rect 227772 996016 265256 996044
rect 227772 996004 227778 996016
rect 265250 996004 265256 996016
rect 265308 996044 265314 996056
rect 267550 996044 267556 996056
rect 265308 996016 267556 996044
rect 265308 996004 265314 996016
rect 267550 996004 267556 996016
rect 267608 996004 267614 996056
rect 280246 996004 280252 996056
rect 280304 996044 280310 996056
rect 315114 996044 315120 996056
rect 280304 996016 315120 996044
rect 280304 996004 280310 996016
rect 315114 996004 315120 996016
rect 315172 996004 315178 996056
rect 365070 996004 365076 996056
rect 365128 996044 365134 996056
rect 371326 996044 371332 996056
rect 365128 996016 371332 996044
rect 365128 996004 365134 996016
rect 371326 996004 371332 996016
rect 371384 996004 371390 996056
rect 625522 996004 625528 996056
rect 625580 996044 625586 996056
rect 625580 996016 631226 996044
rect 625580 996004 625586 996016
rect 154574 995976 154580 995988
rect 136468 995948 154580 995976
rect 86034 995800 86040 995852
rect 86092 995840 86098 995852
rect 100754 995840 100760 995852
rect 86092 995812 100760 995840
rect 86092 995800 86098 995812
rect 100754 995800 100760 995812
rect 100812 995800 100818 995852
rect 136266 995800 136272 995852
rect 136324 995840 136330 995852
rect 136468 995840 136496 995948
rect 154574 995936 154580 995948
rect 154632 995936 154638 995988
rect 211246 995936 211252 995988
rect 211304 995976 211310 995988
rect 215478 995976 215484 995988
rect 211304 995948 215484 995976
rect 211304 995936 211310 995948
rect 215478 995936 215484 995948
rect 215536 995936 215542 995988
rect 307754 995976 307760 995988
rect 286796 995948 307760 995976
rect 151262 995908 151268 995920
rect 136836 995880 151268 995908
rect 136836 995852 136864 995880
rect 151262 995868 151268 995880
rect 151320 995868 151326 995920
rect 198458 995908 198464 995920
rect 188080 995880 198464 995908
rect 136324 995812 136496 995840
rect 136324 995800 136330 995812
rect 136818 995800 136824 995852
rect 136876 995800 136882 995852
rect 137922 995800 137928 995852
rect 137980 995840 137986 995852
rect 150894 995840 150900 995852
rect 137980 995812 150900 995840
rect 137980 995800 137986 995812
rect 150894 995800 150900 995812
rect 150952 995800 150958 995852
rect 91554 995732 91560 995784
rect 91612 995772 91618 995784
rect 92290 995772 92296 995784
rect 91612 995744 92296 995772
rect 91612 995732 91618 995744
rect 92290 995732 92296 995744
rect 92348 995732 92354 995784
rect 139210 995732 139216 995784
rect 139268 995772 139274 995784
rect 152550 995772 152556 995784
rect 139268 995744 152556 995772
rect 139268 995732 139274 995744
rect 152550 995732 152556 995744
rect 152608 995732 152614 995784
rect 184474 995732 184480 995784
rect 184532 995772 184538 995784
rect 188080 995772 188108 995880
rect 198458 995868 198464 995880
rect 198516 995868 198522 995920
rect 246482 995908 246488 995920
rect 239048 995880 246488 995908
rect 239048 995852 239076 995880
rect 246482 995868 246488 995880
rect 246540 995868 246546 995920
rect 286796 995852 286824 995948
rect 307754 995936 307760 995948
rect 307812 995936 307818 995988
rect 362586 995936 362592 995988
rect 362644 995976 362650 995988
rect 367370 995976 367376 995988
rect 362644 995948 367376 995976
rect 362644 995936 362650 995948
rect 367370 995936 367376 995948
rect 367428 995936 367434 995988
rect 383470 995936 383476 995988
rect 383528 995976 383534 995988
rect 383528 995948 391934 995976
rect 383528 995936 383534 995948
rect 306926 995908 306932 995920
rect 293604 995880 306932 995908
rect 293604 995852 293632 995880
rect 306926 995868 306932 995880
rect 306984 995868 306990 995920
rect 383194 995868 383200 995920
rect 383252 995908 383258 995920
rect 383252 995880 389404 995908
rect 383252 995868 383258 995880
rect 188154 995800 188160 995852
rect 188212 995840 188218 995852
rect 198642 995840 198648 995852
rect 188212 995812 198648 995840
rect 188212 995800 188218 995812
rect 198642 995800 198648 995812
rect 198700 995800 198706 995852
rect 239030 995800 239036 995852
rect 239088 995800 239094 995852
rect 239582 995800 239588 995852
rect 239640 995840 239646 995852
rect 254118 995840 254124 995852
rect 239640 995812 254124 995840
rect 239640 995800 239646 995812
rect 254118 995800 254124 995812
rect 254176 995800 254182 995852
rect 286778 995800 286784 995852
rect 286836 995800 286842 995852
rect 293586 995800 293592 995852
rect 293644 995800 293650 995852
rect 295058 995800 295064 995852
rect 295116 995840 295122 995852
rect 310146 995840 310152 995852
rect 295116 995812 310152 995840
rect 295116 995800 295122 995812
rect 310146 995800 310152 995812
rect 310204 995800 310210 995852
rect 389376 995784 389404 995880
rect 391906 995852 391934 995948
rect 566550 995936 566556 995988
rect 566608 995976 566614 995988
rect 576302 995976 576308 995988
rect 566608 995948 576308 995976
rect 566608 995936 566614 995948
rect 576302 995936 576308 995948
rect 576360 995936 576366 995988
rect 625614 995936 625620 995988
rect 625672 995976 625678 995988
rect 625672 995948 630168 995976
rect 625672 995936 625678 995948
rect 472434 995868 472440 995920
rect 472492 995908 472498 995920
rect 472492 995880 474780 995908
rect 472492 995868 472498 995880
rect 474752 995852 474780 995880
rect 523034 995868 523040 995920
rect 523092 995908 523098 995920
rect 523092 995880 528508 995908
rect 523092 995868 523098 995880
rect 528480 995852 528508 995880
rect 625706 995868 625712 995920
rect 625764 995908 625770 995920
rect 625764 995880 627224 995908
rect 625764 995868 625770 995880
rect 627196 995852 627224 995880
rect 391906 995812 391940 995852
rect 391934 995800 391940 995812
rect 391992 995800 391998 995852
rect 396626 995800 396632 995852
rect 396684 995840 396690 995852
rect 400030 995840 400036 995852
rect 396684 995812 400036 995840
rect 396684 995800 396690 995812
rect 400030 995800 400036 995812
rect 400088 995800 400094 995852
rect 472526 995800 472532 995852
rect 472584 995840 472590 995852
rect 473998 995840 474004 995852
rect 472584 995812 474004 995840
rect 472584 995800 472590 995812
rect 473998 995800 474004 995812
rect 474056 995800 474062 995852
rect 474734 995800 474740 995852
rect 474792 995800 474798 995852
rect 485682 995800 485688 995852
rect 485740 995840 485746 995852
rect 488902 995840 488908 995852
rect 485740 995812 488908 995840
rect 485740 995800 485746 995812
rect 488902 995800 488908 995812
rect 488960 995800 488966 995852
rect 523954 995800 523960 995852
rect 524012 995840 524018 995852
rect 524782 995840 524788 995852
rect 524012 995812 524788 995840
rect 524012 995800 524018 995812
rect 524782 995800 524788 995812
rect 524840 995800 524846 995852
rect 528462 995800 528468 995852
rect 528520 995800 528526 995852
rect 537018 995800 537024 995852
rect 537076 995840 537082 995852
rect 540330 995840 540336 995852
rect 537076 995812 540336 995840
rect 537076 995800 537082 995812
rect 540330 995800 540336 995812
rect 540388 995800 540394 995852
rect 625798 995800 625804 995852
rect 625856 995840 625862 995852
rect 626534 995840 626540 995852
rect 625856 995812 626540 995840
rect 625856 995800 625862 995812
rect 626534 995800 626540 995812
rect 626592 995800 626598 995852
rect 627178 995800 627184 995852
rect 627236 995800 627242 995852
rect 630140 995840 630168 995948
rect 630214 995840 630220 995852
rect 630140 995812 630220 995840
rect 630214 995800 630220 995812
rect 630272 995800 630278 995852
rect 631198 995840 631226 996016
rect 631502 995840 631508 995852
rect 631198 995812 631508 995840
rect 631502 995800 631508 995812
rect 631560 995800 631566 995852
rect 184532 995744 188108 995772
rect 184532 995732 184538 995744
rect 194318 995732 194324 995784
rect 194376 995772 194382 995784
rect 195238 995772 195244 995784
rect 194376 995744 195244 995772
rect 194376 995732 194382 995744
rect 195238 995732 195244 995744
rect 195296 995732 195302 995784
rect 245562 995732 245568 995784
rect 245620 995772 245626 995784
rect 246666 995772 246672 995784
rect 245620 995744 246672 995772
rect 245620 995732 245626 995744
rect 246666 995732 246672 995744
rect 246724 995732 246730 995784
rect 383654 995732 383660 995784
rect 383712 995772 383718 995784
rect 384942 995772 384948 995784
rect 383712 995744 384948 995772
rect 383712 995732 383718 995744
rect 384942 995732 384948 995744
rect 385000 995732 385006 995784
rect 389358 995732 389364 995784
rect 389416 995732 389422 995784
rect 472618 995732 472624 995784
rect 472676 995772 472682 995784
rect 473262 995772 473268 995784
rect 472676 995744 473268 995772
rect 472676 995732 472682 995744
rect 473262 995732 473268 995744
rect 473320 995732 473326 995784
rect 524046 995732 524052 995784
rect 524104 995772 524110 995784
rect 525334 995772 525340 995784
rect 524104 995744 525340 995772
rect 524104 995732 524110 995744
rect 525334 995732 525340 995744
rect 525392 995732 525398 995784
rect 620922 995732 620928 995784
rect 620980 995772 620986 995784
rect 627822 995772 627828 995784
rect 620980 995744 627828 995772
rect 620980 995732 620986 995744
rect 627822 995732 627828 995744
rect 627880 995732 627886 995784
rect 89714 995664 89720 995716
rect 89772 995704 89778 995716
rect 92474 995704 92480 995716
rect 89772 995676 92480 995704
rect 89772 995664 89778 995676
rect 92474 995664 92480 995676
rect 92532 995664 92538 995716
rect 190638 995664 190644 995716
rect 190696 995704 190702 995716
rect 195422 995704 195428 995716
rect 190696 995676 195428 995704
rect 190696 995664 190702 995676
rect 195422 995664 195428 995676
rect 195480 995664 195486 995716
rect 243906 995664 243912 995716
rect 243964 995704 243970 995716
rect 246758 995704 246764 995716
rect 243964 995676 246764 995704
rect 243964 995664 243970 995676
rect 246758 995664 246764 995676
rect 246816 995664 246822 995716
rect 291746 995664 291752 995716
rect 291804 995704 291810 995716
rect 306466 995704 306472 995716
rect 291804 995676 306472 995704
rect 291804 995664 291810 995676
rect 306466 995664 306472 995676
rect 306524 995664 306530 995716
rect 383746 995664 383752 995716
rect 383804 995704 383810 995716
rect 384390 995704 384396 995716
rect 383804 995676 384396 995704
rect 383804 995664 383810 995676
rect 384390 995664 384396 995676
rect 384448 995664 384454 995716
rect 472342 995664 472348 995716
rect 472400 995704 472406 995716
rect 476942 995704 476948 995716
rect 472400 995676 476948 995704
rect 472400 995664 472406 995676
rect 476942 995664 476948 995676
rect 477000 995664 477006 995716
rect 523218 995664 523224 995716
rect 523276 995704 523282 995716
rect 529014 995704 529020 995716
rect 523276 995676 529020 995704
rect 523276 995664 523282 995676
rect 529014 995664 529020 995676
rect 529072 995664 529078 995716
rect 625890 995664 625896 995716
rect 625948 995704 625954 995716
rect 630858 995704 630864 995716
rect 625948 995676 630864 995704
rect 625948 995664 625954 995676
rect 630858 995664 630864 995676
rect 630916 995664 630922 995716
rect 77938 995596 77944 995648
rect 77996 995636 78002 995648
rect 92382 995636 92388 995648
rect 77996 995608 92388 995636
rect 77996 995596 78002 995608
rect 92382 995596 92388 995608
rect 92440 995596 92446 995648
rect 133138 995596 133144 995648
rect 133196 995636 133202 995648
rect 152918 995636 152924 995648
rect 133196 995608 152924 995636
rect 133196 995596 133202 995608
rect 152918 995596 152924 995608
rect 152976 995596 152982 995648
rect 189442 995596 189448 995648
rect 189500 995636 189506 995648
rect 195514 995636 195520 995648
rect 189500 995608 195520 995636
rect 189500 995596 189506 995608
rect 195514 995596 195520 995608
rect 195572 995596 195578 995648
rect 240870 995596 240876 995648
rect 240928 995636 240934 995648
rect 253658 995636 253664 995648
rect 240928 995608 253664 995636
rect 240928 995596 240934 995608
rect 253658 995596 253664 995608
rect 253716 995596 253722 995648
rect 287514 995596 287520 995648
rect 287572 995636 287578 995648
rect 307294 995636 307300 995648
rect 287572 995608 307300 995636
rect 287572 995596 287578 995608
rect 307294 995596 307300 995608
rect 307352 995596 307358 995648
rect 383378 995596 383384 995648
rect 383436 995636 383442 995648
rect 385678 995636 385684 995648
rect 383436 995608 385684 995636
rect 383436 995596 383442 995608
rect 385678 995596 385684 995608
rect 385736 995596 385742 995648
rect 469214 995596 469220 995648
rect 469272 995636 469278 995648
rect 481910 995636 481916 995648
rect 469272 995608 481916 995636
rect 469272 995596 469278 995608
rect 481910 995596 481916 995608
rect 481968 995596 481974 995648
rect 521470 995596 521476 995648
rect 521528 995636 521534 995648
rect 532694 995636 532700 995648
rect 521528 995608 532700 995636
rect 521528 995596 521534 995608
rect 532694 995596 532700 995608
rect 532752 995596 532758 995648
rect 623774 995596 623780 995648
rect 623832 995636 623838 995648
rect 635826 995636 635832 995648
rect 623832 995608 635832 995636
rect 623832 995596 623838 995608
rect 635826 995596 635832 995608
rect 635884 995596 635890 995648
rect 88978 995528 88984 995580
rect 89036 995568 89042 995580
rect 92566 995568 92572 995580
rect 89036 995540 92572 995568
rect 89036 995528 89042 995540
rect 92566 995528 92572 995540
rect 92624 995528 92630 995580
rect 132402 995528 132408 995580
rect 132460 995568 132466 995580
rect 153378 995568 153384 995580
rect 132460 995540 153384 995568
rect 132460 995528 132466 995540
rect 153378 995528 153384 995540
rect 153436 995528 153442 995580
rect 184658 995528 184664 995580
rect 184716 995568 184722 995580
rect 198550 995568 198556 995580
rect 184716 995540 198556 995568
rect 184716 995528 184722 995540
rect 198550 995528 198556 995540
rect 198608 995528 198614 995580
rect 383562 995528 383568 995580
rect 383620 995568 383626 995580
rect 387518 995568 387524 995580
rect 383620 995540 387524 995568
rect 383620 995528 383626 995540
rect 387518 995528 387524 995540
rect 387576 995528 387582 995580
rect 469306 995528 469312 995580
rect 469364 995568 469370 995580
rect 482646 995568 482652 995580
rect 469364 995540 482652 995568
rect 469364 995528 469370 995540
rect 482646 995528 482652 995540
rect 482704 995528 482710 995580
rect 521378 995528 521384 995580
rect 521436 995568 521442 995580
rect 533430 995568 533436 995580
rect 521436 995540 533436 995568
rect 521436 995528 521442 995540
rect 533430 995528 533436 995540
rect 533488 995528 533494 995580
rect 130010 995460 130016 995512
rect 130068 995500 130074 995512
rect 143810 995500 143816 995512
rect 130068 995472 143816 995500
rect 130068 995460 130074 995472
rect 143810 995460 143816 995472
rect 143868 995460 143874 995512
rect 188798 995460 188804 995512
rect 188856 995500 188862 995512
rect 195606 995500 195612 995512
rect 188856 995472 195612 995500
rect 188856 995460 188862 995472
rect 195606 995460 195612 995472
rect 195664 995460 195670 995512
rect 383286 995460 383292 995512
rect 383344 995500 383350 995512
rect 388622 995500 388628 995512
rect 383344 995472 388628 995500
rect 383344 995460 383350 995472
rect 388622 995460 388628 995472
rect 388680 995460 388686 995512
rect 393590 995500 393596 995512
rect 391906 995472 393596 995500
rect 131850 995392 131856 995444
rect 131908 995432 131914 995444
rect 146018 995432 146024 995444
rect 131908 995404 146024 995432
rect 131908 995392 131914 995404
rect 146018 995392 146024 995404
rect 146076 995392 146082 995444
rect 183830 995392 183836 995444
rect 183888 995432 183894 995444
rect 198366 995432 198372 995444
rect 183888 995404 198372 995432
rect 183888 995392 183894 995404
rect 198366 995392 198372 995404
rect 198424 995392 198430 995444
rect 381262 995392 381268 995444
rect 381320 995432 381326 995444
rect 391906 995432 391934 995472
rect 393590 995460 393596 995472
rect 393648 995460 393654 995512
rect 381320 995404 391934 995432
rect 381320 995392 381326 995404
rect 183278 995324 183284 995376
rect 183336 995364 183342 995376
rect 195974 995364 195980 995376
rect 183336 995336 195980 995364
rect 183336 995324 183342 995336
rect 195974 995324 195980 995336
rect 196032 995324 196038 995376
rect 180472 995256 180478 995308
rect 180530 995296 180536 995308
rect 195698 995296 195704 995308
rect 180530 995268 195704 995296
rect 180530 995256 180536 995268
rect 195698 995256 195704 995268
rect 195756 995256 195762 995308
rect 303522 994720 303528 994772
rect 303580 994720 303586 994772
rect 283466 993828 283472 993880
rect 283524 993868 283530 993880
rect 301774 993868 301780 993880
rect 283524 993840 301780 993868
rect 283524 993828 283530 993840
rect 301774 993828 301780 993840
rect 301832 993828 301838 993880
rect 378318 993828 378324 993880
rect 378376 993868 378382 993880
rect 392670 993868 392676 993880
rect 378376 993840 392676 993868
rect 378376 993828 378382 993840
rect 392670 993828 392676 993840
rect 392728 993828 392734 993880
rect 146110 993800 146116 993812
rect 129706 993772 146116 993800
rect 129090 993692 129096 993744
rect 129148 993732 129154 993744
rect 129706 993732 129734 993772
rect 146110 993760 146116 993772
rect 146168 993760 146174 993812
rect 285950 993760 285956 993812
rect 286008 993800 286014 993812
rect 314838 993800 314844 993812
rect 286008 993772 314844 993800
rect 286008 993760 286014 993772
rect 314838 993760 314844 993772
rect 314896 993760 314902 993812
rect 469766 993760 469772 993812
rect 469824 993800 469830 993812
rect 487798 993800 487804 993812
rect 469824 993772 487804 993800
rect 469824 993760 469830 993772
rect 487798 993760 487804 993772
rect 487856 993760 487862 993812
rect 520550 993760 520556 993812
rect 520608 993800 520614 993812
rect 535546 993800 535552 993812
rect 520608 993772 535552 993800
rect 520608 993760 520614 993772
rect 535546 993760 535552 993772
rect 535604 993760 535610 993812
rect 129148 993704 129734 993732
rect 129148 993692 129154 993704
rect 140498 993692 140504 993744
rect 140556 993732 140562 993744
rect 151814 993732 151820 993744
rect 140556 993704 151820 993732
rect 140556 993692 140562 993704
rect 151814 993692 151820 993704
rect 151872 993692 151878 993744
rect 180150 993692 180156 993744
rect 180208 993732 180214 993744
rect 207014 993732 207020 993744
rect 180208 993704 207020 993732
rect 180208 993692 180214 993704
rect 207014 993692 207020 993704
rect 207072 993692 207078 993744
rect 284110 993692 284116 993744
rect 284168 993732 284174 993744
rect 315022 993732 315028 993744
rect 284168 993704 315028 993732
rect 284168 993692 284174 993704
rect 315022 993692 315028 993704
rect 315080 993692 315086 993744
rect 374546 993692 374552 993744
rect 374604 993732 374610 993744
rect 393314 993732 393320 993744
rect 374604 993704 393320 993732
rect 374604 993692 374610 993704
rect 393314 993692 393320 993704
rect 393372 993692 393378 993744
rect 471054 993692 471060 993744
rect 471112 993732 471118 993744
rect 484118 993732 484124 993744
rect 471112 993704 484124 993732
rect 471112 993692 471118 993704
rect 484118 993692 484124 993704
rect 484176 993692 484182 993744
rect 574094 993692 574100 993744
rect 574152 993732 574158 993744
rect 633986 993732 633992 993744
rect 574152 993704 633992 993732
rect 574152 993692 574158 993704
rect 633986 993692 633992 993704
rect 634044 993692 634050 993744
rect 77018 993624 77024 993676
rect 77076 993664 77082 993676
rect 104158 993664 104164 993676
rect 77076 993636 104164 993664
rect 77076 993624 77082 993636
rect 104158 993624 104164 993636
rect 104216 993624 104222 993676
rect 128446 993624 128452 993676
rect 128504 993664 128510 993676
rect 160278 993664 160284 993676
rect 128504 993636 160284 993664
rect 128504 993624 128510 993636
rect 160278 993624 160284 993636
rect 160336 993624 160342 993676
rect 181438 993624 181444 993676
rect 181496 993664 181502 993676
rect 207750 993664 207756 993676
rect 181496 993636 207756 993664
rect 181496 993624 181502 993636
rect 207750 993624 207756 993636
rect 207808 993624 207814 993676
rect 231578 993624 231584 993676
rect 231636 993664 231642 993676
rect 262214 993664 262220 993676
rect 231636 993636 262220 993664
rect 231636 993624 231642 993636
rect 262214 993624 262220 993636
rect 262272 993624 262278 993676
rect 282822 993624 282828 993676
rect 282880 993664 282886 993676
rect 314930 993664 314936 993676
rect 282880 993636 314936 993664
rect 282880 993624 282886 993636
rect 314930 993624 314936 993636
rect 314988 993624 314994 993676
rect 359182 993624 359188 993676
rect 359240 993664 359246 993676
rect 398834 993664 398840 993676
rect 359240 993636 398840 993664
rect 359240 993624 359246 993636
rect 398834 993624 398840 993636
rect 398892 993624 398898 993676
rect 462590 993624 462596 993676
rect 462648 993664 462654 993676
rect 485958 993664 485964 993676
rect 462648 993636 485964 993664
rect 462648 993624 462654 993636
rect 485958 993624 485964 993636
rect 486016 993624 486022 993676
rect 503622 993624 503628 993676
rect 503680 993664 503686 993676
rect 539226 993664 539232 993676
rect 503680 993636 539232 993664
rect 503680 993624 503686 993636
rect 539226 993624 539232 993636
rect 539284 993624 539290 993676
rect 555050 993624 555056 993676
rect 555108 993664 555114 993676
rect 640702 993664 640708 993676
rect 555108 993636 640708 993664
rect 555108 993624 555114 993636
rect 640702 993624 640708 993636
rect 640760 993624 640766 993676
rect 433518 993556 433524 993608
rect 433576 993596 433582 993608
rect 434714 993596 434720 993608
rect 433576 993568 434720 993596
rect 433576 993556 433582 993568
rect 434714 993556 434720 993568
rect 434772 993596 434778 993608
rect 510890 993596 510896 993608
rect 434772 993568 510896 993596
rect 434772 993556 434778 993568
rect 510890 993556 510896 993568
rect 510948 993556 510954 993608
rect 510982 993556 510988 993608
rect 511040 993596 511046 993608
rect 512086 993596 512092 993608
rect 511040 993568 512092 993596
rect 511040 993556 511046 993568
rect 512086 993556 512092 993568
rect 512144 993596 512150 993608
rect 558546 993596 558552 993608
rect 512144 993568 558552 993596
rect 512144 993556 512150 993568
rect 558546 993556 558552 993568
rect 558604 993556 558610 993608
rect 367370 993488 367376 993540
rect 367428 993528 367434 993540
rect 368566 993528 368572 993540
rect 367428 993500 368572 993528
rect 367428 993488 367434 993500
rect 368566 993488 368572 993500
rect 368624 993528 368630 993540
rect 433334 993528 433340 993540
rect 368624 993500 433340 993528
rect 368624 993488 368630 993500
rect 433334 993488 433340 993500
rect 433392 993488 433398 993540
rect 433610 993488 433616 993540
rect 433668 993528 433674 993540
rect 434806 993528 434812 993540
rect 433668 993500 434812 993528
rect 433668 993488 433674 993500
rect 434806 993488 434812 993500
rect 434864 993528 434870 993540
rect 510706 993528 510712 993540
rect 434864 993500 510712 993528
rect 434864 993488 434870 993500
rect 510706 993488 510712 993500
rect 510764 993488 510770 993540
rect 510798 993488 510804 993540
rect 510856 993528 510862 993540
rect 511902 993528 511908 993540
rect 510856 993500 511908 993528
rect 510856 993488 510862 993500
rect 511902 993488 511908 993500
rect 511960 993528 511966 993540
rect 557718 993528 557724 993540
rect 511960 993500 557724 993528
rect 511960 993488 511966 993500
rect 557718 993488 557724 993500
rect 557776 993488 557782 993540
rect 367278 993420 367284 993472
rect 367336 993460 367342 993472
rect 368382 993460 368388 993472
rect 367336 993432 368388 993460
rect 367336 993420 367342 993432
rect 368382 993420 368388 993432
rect 368440 993420 368446 993472
rect 368750 993420 368756 993472
rect 368808 993460 368814 993472
rect 433426 993460 433432 993472
rect 368808 993432 433432 993460
rect 368808 993420 368814 993432
rect 433426 993420 433432 993432
rect 433484 993420 433490 993472
rect 436186 993420 436192 993472
rect 436244 993460 436250 993472
rect 437934 993460 437940 993472
rect 436244 993432 437940 993460
rect 436244 993420 436250 993432
rect 437934 993420 437940 993432
rect 437992 993460 437998 993472
rect 513650 993460 513656 993472
rect 437992 993432 513656 993460
rect 437992 993420 437998 993432
rect 513650 993420 513656 993432
rect 513708 993420 513714 993472
rect 513742 993420 513748 993472
rect 513800 993460 513806 993472
rect 515214 993460 515220 993472
rect 513800 993432 515220 993460
rect 513800 993420 513806 993432
rect 515214 993420 515220 993432
rect 515272 993460 515278 993472
rect 565814 993460 565820 993472
rect 515272 993432 565820 993460
rect 515272 993420 515278 993432
rect 565814 993420 565820 993432
rect 565872 993420 565878 993472
rect 368400 993392 368428 993420
rect 436094 993392 436100 993404
rect 368400 993364 436100 993392
rect 436094 993352 436100 993364
rect 436152 993352 436158 993404
rect 367462 992536 367468 992588
rect 367520 992576 367526 992588
rect 368750 992576 368756 992588
rect 367520 992548 368756 992576
rect 367520 992536 367526 992548
rect 368750 992536 368756 992548
rect 368808 992536 368814 992588
rect 116026 990836 116032 990888
rect 116084 990876 116090 990888
rect 116084 990848 121408 990876
rect 116084 990836 116090 990848
rect 121380 990808 121408 990848
rect 122098 990808 122104 990820
rect 121380 990780 122104 990808
rect 122098 990768 122104 990780
rect 122156 990768 122162 990820
rect 168374 990632 168380 990684
rect 168432 990672 168438 990684
rect 170398 990672 170404 990684
rect 168432 990644 170404 990672
rect 168432 990632 168438 990644
rect 170398 990632 170404 990644
rect 170456 990632 170462 990684
rect 203150 990632 203156 990684
rect 203208 990672 203214 990684
rect 204162 990672 204168 990684
rect 203208 990644 204168 990672
rect 203208 990632 203214 990644
rect 204162 990632 204168 990644
rect 204220 990632 204226 990684
rect 331214 990632 331220 990684
rect 331272 990672 331278 990684
rect 332686 990672 332692 990684
rect 331272 990644 332692 990672
rect 331272 990632 331278 990644
rect 332686 990632 332692 990644
rect 332744 990632 332750 990684
rect 89622 990088 89628 990140
rect 89680 990128 89686 990140
rect 92474 990128 92480 990140
rect 89680 990100 92480 990128
rect 89680 990088 89686 990100
rect 92474 990088 92480 990100
rect 92532 990088 92538 990140
rect 366174 989680 366180 989732
rect 366232 989720 366238 989732
rect 381630 989720 381636 989732
rect 366232 989692 381636 989720
rect 366232 989680 366238 989692
rect 381630 989680 381636 989692
rect 381688 989680 381694 989732
rect 434622 989680 434628 989732
rect 434680 989720 434686 989732
rect 446490 989720 446496 989732
rect 434680 989692 446496 989720
rect 434680 989680 434686 989692
rect 446490 989680 446496 989692
rect 446548 989680 446554 989732
rect 371142 989612 371148 989664
rect 371200 989652 371206 989664
rect 397822 989652 397828 989664
rect 371200 989624 397828 989652
rect 371200 989612 371206 989624
rect 397822 989612 397828 989624
rect 397880 989612 397886 989664
rect 437566 989612 437572 989664
rect 437624 989652 437630 989664
rect 462774 989652 462780 989664
rect 437624 989624 462780 989652
rect 437624 989612 437630 989624
rect 462774 989612 462780 989624
rect 462832 989612 462838 989664
rect 514662 989612 514668 989664
rect 514720 989652 514726 989664
rect 527634 989652 527640 989664
rect 514720 989624 527640 989652
rect 514720 989612 514726 989624
rect 527634 989612 527640 989624
rect 527692 989612 527698 989664
rect 567470 989612 567476 989664
rect 567528 989652 567534 989664
rect 592494 989652 592500 989664
rect 567528 989624 592500 989652
rect 567528 989612 567534 989624
rect 592494 989612 592500 989624
rect 592552 989612 592558 989664
rect 321462 989544 321468 989596
rect 321520 989584 321526 989596
rect 349154 989584 349160 989596
rect 321520 989556 349160 989584
rect 321520 989544 321526 989556
rect 349154 989544 349160 989556
rect 349212 989544 349218 989596
rect 371510 989544 371516 989596
rect 371568 989584 371574 989596
rect 414106 989584 414112 989596
rect 371568 989556 414112 989584
rect 371568 989544 371574 989556
rect 414106 989544 414112 989556
rect 414164 989544 414170 989596
rect 437750 989544 437756 989596
rect 437808 989584 437814 989596
rect 478966 989584 478972 989596
rect 437808 989556 478972 989584
rect 437808 989544 437814 989556
rect 478966 989544 478972 989556
rect 479024 989544 479030 989596
rect 515030 989544 515036 989596
rect 515088 989584 515094 989596
rect 543826 989584 543832 989596
rect 515088 989556 543832 989584
rect 515088 989544 515094 989556
rect 543826 989544 543832 989556
rect 543884 989544 543890 989596
rect 567286 989544 567292 989596
rect 567344 989584 567350 989596
rect 608778 989584 608784 989596
rect 567344 989556 608784 989584
rect 567344 989544 567350 989556
rect 608778 989544 608784 989556
rect 608836 989544 608842 989596
rect 269206 989476 269212 989528
rect 269264 989516 269270 989528
rect 300486 989516 300492 989528
rect 269264 989488 300492 989516
rect 269264 989476 269270 989488
rect 300486 989476 300492 989488
rect 300544 989476 300550 989528
rect 319070 989476 319076 989528
rect 319128 989516 319134 989528
rect 365438 989516 365444 989528
rect 319128 989488 365444 989516
rect 319128 989476 319134 989488
rect 365438 989476 365444 989488
rect 365496 989476 365502 989528
rect 371326 989476 371332 989528
rect 371384 989516 371390 989528
rect 430298 989516 430304 989528
rect 371384 989488 430304 989516
rect 371384 989476 371390 989488
rect 430298 989476 430304 989488
rect 430356 989476 430362 989528
rect 437382 989476 437388 989528
rect 437440 989516 437446 989528
rect 495158 989516 495164 989528
rect 437440 989488 495164 989516
rect 437440 989476 437446 989488
rect 495158 989476 495164 989488
rect 495216 989476 495222 989528
rect 514846 989476 514852 989528
rect 514904 989516 514910 989528
rect 560110 989516 560116 989528
rect 514904 989488 560116 989516
rect 514904 989476 514910 989488
rect 560110 989476 560116 989488
rect 560168 989476 560174 989528
rect 567102 989476 567108 989528
rect 567160 989516 567166 989528
rect 624970 989516 624976 989528
rect 567160 989488 624976 989516
rect 567160 989476 567166 989488
rect 624970 989476 624976 989488
rect 625028 989476 625034 989528
rect 73430 989408 73436 989460
rect 73488 989448 73494 989460
rect 92934 989448 92940 989460
rect 73488 989420 92940 989448
rect 73488 989408 73494 989420
rect 92934 989408 92940 989420
rect 92992 989408 92998 989460
rect 105814 989408 105820 989460
rect 105872 989448 105878 989460
rect 113266 989448 113272 989460
rect 105872 989420 113272 989448
rect 105872 989408 105878 989420
rect 113266 989408 113272 989420
rect 113324 989408 113330 989460
rect 151814 989408 151820 989460
rect 151872 989448 151878 989460
rect 186958 989448 186964 989460
rect 151872 989420 186964 989448
rect 151872 989408 151878 989420
rect 186958 989408 186964 989420
rect 187016 989408 187022 989460
rect 216582 989408 216588 989460
rect 216640 989448 216646 989460
rect 235626 989448 235632 989460
rect 216640 989420 235632 989448
rect 216640 989408 216646 989420
rect 235626 989408 235632 989420
rect 235684 989408 235690 989460
rect 269022 989408 269028 989460
rect 269080 989448 269086 989460
rect 284294 989448 284300 989460
rect 269080 989420 284300 989448
rect 269080 989408 269086 989420
rect 284294 989408 284300 989420
rect 284352 989408 284358 989460
rect 303522 989408 303528 989460
rect 303580 989448 303586 989460
rect 666554 989448 666560 989460
rect 303580 989420 666560 989448
rect 303580 989408 303586 989420
rect 666554 989408 666560 989420
rect 666612 989408 666618 989460
rect 138290 988728 138296 988780
rect 138348 988768 138354 988780
rect 144822 988768 144828 988780
rect 138348 988740 144828 988768
rect 138348 988728 138354 988740
rect 144822 988728 144828 988740
rect 144880 988728 144886 988780
rect 505646 988252 505652 988304
rect 505704 988292 505710 988304
rect 511442 988292 511448 988304
rect 505704 988264 511448 988292
rect 505704 988252 505710 988264
rect 511442 988252 511448 988264
rect 511500 988252 511506 988304
rect 248322 988116 248328 988168
rect 248380 988156 248386 988168
rect 251818 988156 251824 988168
rect 248380 988128 251824 988156
rect 248380 988116 248386 988128
rect 251818 988116 251824 988128
rect 251876 988116 251882 988168
rect 45462 987980 45468 988032
rect 45520 988020 45526 988032
rect 367186 988020 367192 988032
rect 45520 987992 367192 988020
rect 45520 987980 45526 987992
rect 367186 987980 367192 987992
rect 367244 987980 367250 988032
rect 45738 987912 45744 987964
rect 45796 987952 45802 987964
rect 368750 987952 368756 987964
rect 45796 987924 368756 987952
rect 45796 987912 45802 987924
rect 368750 987912 368756 987924
rect 368808 987912 368814 987964
rect 45554 987844 45560 987896
rect 45612 987884 45618 987896
rect 369854 987884 369860 987896
rect 45612 987856 369860 987884
rect 45612 987844 45618 987856
rect 369854 987844 369860 987856
rect 369912 987844 369918 987896
rect 318886 987776 318892 987828
rect 318944 987816 318950 987828
rect 666646 987816 666652 987828
rect 318944 987788 666652 987816
rect 318944 987776 318950 987788
rect 666646 987776 666652 987788
rect 666704 987776 666710 987828
rect 317506 987708 317512 987760
rect 317564 987748 317570 987760
rect 666922 987748 666928 987760
rect 317564 987720 666928 987748
rect 317564 987708 317570 987720
rect 666922 987708 666928 987720
rect 666980 987708 666986 987760
rect 318702 987640 318708 987692
rect 318760 987680 318766 987692
rect 669222 987680 669228 987692
rect 318760 987652 669228 987680
rect 318760 987640 318766 987652
rect 669222 987640 669228 987652
rect 669280 987640 669286 987692
rect 315114 987572 315120 987624
rect 315172 987612 315178 987624
rect 666738 987612 666744 987624
rect 315172 987584 666744 987612
rect 315172 987572 315178 987584
rect 666738 987572 666744 987584
rect 666796 987572 666802 987624
rect 280062 987504 280068 987556
rect 280120 987544 280126 987556
rect 651374 987544 651380 987556
rect 280120 987516 651380 987544
rect 280120 987504 280126 987516
rect 651374 987504 651380 987516
rect 651432 987504 651438 987556
rect 270402 987436 270408 987488
rect 270460 987476 270466 987488
rect 652846 987476 652852 987488
rect 270460 987448 652852 987476
rect 270460 987436 270466 987448
rect 652846 987436 652852 987448
rect 652904 987436 652910 987488
rect 267642 987368 267648 987420
rect 267700 987408 267706 987420
rect 652662 987408 652668 987420
rect 267700 987380 652668 987408
rect 267700 987368 267706 987380
rect 652662 987368 652668 987380
rect 652720 987368 652726 987420
rect 48222 987300 48228 987352
rect 48280 987340 48286 987352
rect 433518 987340 433524 987352
rect 48280 987312 433524 987340
rect 48280 987300 48286 987312
rect 433518 987300 433524 987312
rect 433576 987300 433582 987352
rect 267550 987232 267556 987284
rect 267608 987272 267614 987284
rect 652754 987272 652760 987284
rect 267608 987244 652760 987272
rect 267608 987232 267614 987244
rect 652754 987232 652760 987244
rect 652812 987232 652818 987284
rect 227622 987164 227628 987216
rect 227680 987204 227686 987216
rect 651558 987204 651564 987216
rect 227680 987176 651564 987204
rect 227680 987164 227686 987176
rect 651558 987164 651564 987176
rect 651616 987164 651622 987216
rect 215478 987096 215484 987148
rect 215536 987136 215542 987148
rect 658274 987136 658280 987148
rect 215536 987108 658280 987136
rect 215536 987096 215542 987108
rect 658274 987096 658280 987108
rect 658332 987096 658338 987148
rect 212810 987028 212816 987080
rect 212868 987068 212874 987080
rect 658182 987068 658188 987080
rect 212868 987040 658188 987068
rect 212868 987028 212874 987040
rect 658182 987028 658188 987040
rect 658240 987028 658246 987080
rect 175182 986960 175188 987012
rect 175240 987000 175246 987012
rect 651650 987000 651656 987012
rect 175240 986972 651656 987000
rect 175240 986960 175246 986972
rect 651650 986960 651656 986972
rect 651708 986960 651714 987012
rect 125502 986892 125508 986944
rect 125560 986932 125566 986944
rect 651466 986932 651472 986944
rect 125560 986904 651472 986932
rect 125560 986892 125566 986904
rect 651466 986892 651472 986904
rect 651524 986892 651530 986944
rect 62666 986824 62672 986876
rect 62724 986864 62730 986876
rect 113174 986864 113180 986876
rect 62724 986836 113180 986864
rect 62724 986824 62730 986836
rect 113174 986824 113180 986836
rect 113232 986864 113238 986876
rect 669498 986864 669504 986876
rect 113232 986836 669504 986864
rect 113232 986824 113238 986836
rect 669498 986824 669504 986836
rect 669556 986824 669562 986876
rect 62298 986756 62304 986808
rect 62356 986796 62362 986808
rect 110598 986796 110604 986808
rect 62356 986768 110604 986796
rect 62356 986756 62362 986768
rect 110598 986756 110604 986768
rect 110656 986796 110662 986808
rect 669406 986796 669412 986808
rect 110656 986768 669412 986796
rect 110656 986756 110662 986768
rect 669406 986756 669412 986768
rect 669464 986756 669470 986808
rect 62482 986688 62488 986740
rect 62540 986728 62546 986740
rect 110782 986728 110788 986740
rect 62540 986700 110788 986728
rect 62540 986688 62546 986700
rect 110782 986688 110788 986700
rect 110840 986728 110846 986740
rect 669314 986728 669320 986740
rect 110840 986700 669320 986728
rect 110840 986688 110846 986700
rect 669314 986688 669320 986700
rect 669372 986688 669378 986740
rect 564526 985532 564532 985584
rect 564584 985572 564590 985584
rect 564710 985572 564716 985584
rect 564584 985544 564716 985572
rect 564584 985532 564590 985544
rect 564710 985532 564716 985544
rect 564768 985572 564774 985584
rect 675662 985572 675668 985584
rect 564768 985544 675668 985572
rect 564768 985532 564774 985544
rect 675662 985532 675668 985544
rect 675720 985532 675726 985584
rect 62850 985464 62856 985516
rect 62908 985504 62914 985516
rect 669590 985504 669596 985516
rect 62908 985476 669596 985504
rect 62908 985464 62914 985476
rect 669590 985464 669596 985476
rect 669648 985464 669654 985516
rect 62574 985396 62580 985448
rect 62632 985436 62638 985448
rect 670418 985436 670424 985448
rect 62632 985408 670424 985436
rect 62632 985396 62638 985408
rect 670418 985396 670424 985408
rect 670476 985396 670482 985448
rect 46474 985328 46480 985380
rect 46532 985368 46538 985380
rect 668762 985368 668768 985380
rect 46532 985340 668768 985368
rect 46532 985328 46538 985340
rect 668762 985328 668768 985340
rect 668820 985328 668826 985380
rect 350258 985124 350264 985176
rect 350316 985164 350322 985176
rect 670970 985164 670976 985176
rect 350316 985136 670976 985164
rect 350316 985124 350322 985136
rect 670970 985124 670976 985136
rect 671028 985124 671034 985176
rect 45646 985056 45652 985108
rect 45704 985096 45710 985108
rect 367094 985096 367100 985108
rect 45704 985068 367100 985096
rect 45704 985056 45710 985068
rect 367094 985056 367100 985068
rect 367152 985056 367158 985108
rect 45922 984988 45928 985040
rect 45980 985028 45986 985040
rect 368566 985028 368572 985040
rect 45980 985000 368572 985028
rect 45980 984988 45986 985000
rect 368566 984988 368572 985000
rect 368624 984988 368630 985040
rect 45830 984920 45836 984972
rect 45888 984960 45894 984972
rect 368382 984960 368388 984972
rect 45888 984932 368388 984960
rect 45888 984920 45894 984932
rect 368382 984920 368388 984932
rect 368440 984920 368446 984972
rect 419442 984920 419448 984972
rect 419500 984960 419506 984972
rect 670878 984960 670884 984972
rect 419500 984932 670884 984960
rect 419500 984920 419506 984932
rect 670878 984920 670884 984932
rect 670936 984920 670942 984972
rect 317414 984852 317420 984904
rect 317472 984892 317478 984904
rect 666830 984892 666836 984904
rect 317472 984864 666836 984892
rect 317472 984852 317478 984864
rect 666830 984852 666836 984864
rect 666888 984852 666894 984904
rect 315942 984784 315948 984836
rect 316000 984824 316006 984836
rect 671982 984824 671988 984836
rect 316000 984796 671988 984824
rect 316000 984784 316006 984796
rect 671982 984784 671988 984796
rect 672040 984784 672046 984836
rect 300762 984716 300768 984768
rect 300820 984756 300826 984768
rect 671062 984756 671068 984768
rect 300820 984728 671068 984756
rect 300820 984716 300826 984728
rect 671062 984716 671068 984728
rect 671120 984716 671126 984768
rect 46106 984648 46112 984700
rect 46164 984688 46170 984700
rect 433610 984688 433616 984700
rect 46164 984660 433616 984688
rect 46164 984648 46170 984660
rect 433610 984648 433616 984660
rect 433668 984648 433674 984700
rect 48314 984580 48320 984632
rect 48372 984620 48378 984632
rect 436186 984620 436192 984632
rect 48372 984592 436192 984620
rect 48372 984580 48378 984592
rect 436186 984580 436192 984592
rect 436244 984580 436250 984632
rect 496722 984580 496728 984632
rect 496780 984620 496786 984632
rect 670786 984620 670792 984632
rect 496780 984592 670792 984620
rect 496780 984580 496786 984592
rect 670786 984580 670792 984592
rect 670844 984580 670850 984632
rect 212626 984512 212632 984564
rect 212684 984552 212690 984564
rect 652938 984552 652944 984564
rect 212684 984524 652944 984552
rect 212684 984512 212690 984524
rect 652938 984512 652944 984524
rect 652996 984512 653002 984564
rect 46382 984444 46388 984496
rect 46440 984484 46446 984496
rect 510982 984484 510988 984496
rect 46440 984456 510988 984484
rect 46440 984444 46446 984456
rect 510982 984444 510988 984456
rect 511040 984444 511046 984496
rect 46198 984376 46204 984428
rect 46256 984416 46262 984428
rect 510798 984416 510804 984428
rect 46256 984388 510804 984416
rect 46256 984376 46262 984388
rect 510798 984376 510804 984388
rect 510856 984376 510862 984428
rect 48406 984308 48412 984360
rect 48464 984348 48470 984360
rect 513742 984348 513748 984360
rect 48464 984320 513748 984348
rect 48464 984308 48470 984320
rect 513742 984308 513748 984320
rect 513800 984308 513806 984360
rect 546310 984308 546316 984360
rect 546368 984348 546374 984360
rect 670694 984348 670700 984360
rect 546368 984320 670700 984348
rect 546368 984308 546374 984320
rect 670694 984308 670700 984320
rect 670752 984308 670758 984360
rect 162854 984240 162860 984292
rect 162912 984280 162918 984292
rect 655422 984280 655428 984292
rect 162912 984252 655428 984280
rect 162912 984240 162918 984252
rect 655422 984240 655428 984252
rect 655480 984240 655486 984292
rect 162946 984172 162952 984224
rect 163004 984212 163010 984224
rect 658458 984212 658464 984224
rect 163004 984184 658464 984212
rect 163004 984172 163010 984184
rect 658458 984172 658464 984184
rect 658516 984172 658522 984224
rect 46014 984104 46020 984156
rect 46072 984144 46078 984156
rect 110414 984144 110420 984156
rect 46072 984116 110420 984144
rect 46072 984104 46078 984116
rect 110414 984104 110420 984116
rect 110472 984104 110478 984156
rect 160186 984104 160192 984156
rect 160244 984144 160250 984156
rect 658366 984144 658372 984156
rect 160244 984116 658372 984144
rect 160244 984104 160250 984116
rect 658366 984104 658372 984116
rect 658424 984104 658430 984156
rect 62022 984036 62028 984088
rect 62080 984076 62086 984088
rect 561674 984076 561680 984088
rect 62080 984048 561680 984076
rect 62080 984036 62086 984048
rect 561674 984036 561680 984048
rect 561732 984036 561738 984088
rect 564342 984036 564348 984088
rect 564400 984076 564406 984088
rect 649902 984076 649908 984088
rect 564400 984048 649908 984076
rect 564400 984036 564406 984048
rect 649902 984036 649908 984048
rect 649960 984036 649966 984088
rect 62114 983968 62120 984020
rect 62172 984008 62178 984020
rect 564526 984008 564532 984020
rect 62172 983980 564532 984008
rect 62172 983968 62178 983980
rect 564526 983968 564532 983980
rect 564584 983968 564590 984020
rect 62206 983900 62212 983952
rect 62264 983940 62270 983952
rect 564434 983940 564440 983952
rect 62264 983912 564440 983940
rect 62264 983900 62270 983912
rect 564434 983900 564440 983912
rect 564492 983900 564498 983952
rect 62390 982948 62396 983000
rect 62448 982988 62454 983000
rect 669038 982988 669044 983000
rect 62448 982960 669044 982988
rect 62448 982948 62454 982960
rect 669038 982948 669044 982960
rect 669096 982948 669102 983000
rect 62758 982880 62764 982932
rect 62816 982920 62822 982932
rect 668670 982920 668676 982932
rect 62816 982892 668676 982920
rect 62816 982880 62822 982892
rect 668670 982880 668676 982892
rect 668728 982880 668734 982932
rect 42334 972884 42340 972936
rect 42392 972924 42398 972936
rect 58434 972924 58440 972936
rect 42392 972896 58440 972924
rect 42392 972884 42398 972896
rect 58434 972884 58440 972896
rect 58492 972884 58498 972936
rect 674834 970096 674840 970148
rect 674892 970136 674898 970148
rect 675662 970136 675668 970148
rect 674892 970108 675668 970136
rect 674892 970096 674898 970108
rect 675662 970096 675668 970108
rect 675720 970096 675726 970148
rect 42150 967240 42156 967292
rect 42208 967280 42214 967292
rect 42334 967280 42340 967292
rect 42208 967252 42340 967280
rect 42208 967240 42214 967252
rect 42334 967240 42340 967252
rect 42392 967240 42398 967292
rect 42058 967036 42064 967088
rect 42116 967076 42122 967088
rect 42794 967076 42800 967088
rect 42116 967048 42800 967076
rect 42116 967036 42122 967048
rect 42794 967036 42800 967048
rect 42852 967036 42858 967088
rect 674742 966152 674748 966204
rect 674800 966192 674806 966204
rect 675386 966192 675392 966204
rect 674800 966164 675392 966192
rect 674800 966152 674806 966164
rect 675386 966152 675392 966164
rect 675444 966152 675450 966204
rect 673546 965744 673552 965796
rect 673604 965784 673610 965796
rect 675386 965784 675392 965796
rect 673604 965756 675392 965784
rect 673604 965744 673610 965756
rect 675386 965744 675392 965756
rect 675444 965744 675450 965796
rect 673730 964996 673736 965048
rect 673788 965036 673794 965048
rect 675478 965036 675484 965048
rect 673788 965008 675484 965036
rect 673788 964996 673794 965008
rect 675478 964996 675484 965008
rect 675536 964996 675542 965048
rect 42150 963976 42156 964028
rect 42208 964016 42214 964028
rect 42978 964016 42984 964028
rect 42208 963988 42984 964016
rect 42208 963976 42214 963988
rect 42978 963976 42984 963988
rect 43036 963976 43042 964028
rect 673914 963160 673920 963212
rect 673972 963200 673978 963212
rect 675386 963200 675392 963212
rect 673972 963172 675392 963200
rect 673972 963160 673978 963172
rect 675386 963160 675392 963172
rect 675444 963160 675450 963212
rect 42150 962616 42156 962668
rect 42208 962656 42214 962668
rect 42886 962656 42892 962668
rect 42208 962628 42892 962656
rect 42208 962616 42214 962628
rect 42886 962616 42892 962628
rect 42944 962616 42950 962668
rect 673638 962480 673644 962532
rect 673696 962520 673702 962532
rect 675478 962520 675484 962532
rect 673696 962492 675484 962520
rect 673696 962480 673702 962492
rect 675478 962480 675484 962492
rect 675536 962480 675542 962532
rect 42150 962072 42156 962124
rect 42208 962112 42214 962124
rect 43070 962112 43076 962124
rect 42208 962084 43076 962112
rect 42208 962072 42214 962084
rect 43070 962072 43076 962084
rect 43128 962072 43134 962124
rect 673454 962004 673460 962056
rect 673512 962044 673518 962056
rect 675386 962044 675392 962056
rect 673512 962016 675392 962044
rect 673512 962004 673518 962016
rect 675386 962004 675392 962016
rect 675444 962004 675450 962056
rect 673822 961324 673828 961376
rect 673880 961364 673886 961376
rect 675386 961364 675392 961376
rect 673880 961336 675392 961364
rect 673880 961324 673886 961336
rect 675386 961324 675392 961336
rect 675444 961324 675450 961376
rect 48498 960508 48504 960560
rect 48556 960548 48562 960560
rect 57974 960548 57980 960560
rect 48556 960520 57980 960548
rect 48556 960508 48562 960520
rect 57974 960508 57980 960520
rect 58032 960508 58038 960560
rect 655606 960508 655612 960560
rect 655664 960548 655670 960560
rect 675018 960548 675024 960560
rect 655664 960520 675024 960548
rect 655664 960508 655670 960520
rect 675018 960508 675024 960520
rect 675076 960508 675082 960560
rect 42886 959624 42892 959676
rect 42944 959664 42950 959676
rect 43622 959664 43628 959676
rect 42944 959636 43628 959664
rect 42944 959624 42950 959636
rect 43622 959624 43628 959636
rect 43680 959624 43686 959676
rect 42058 959488 42064 959540
rect 42116 959528 42122 959540
rect 42886 959528 42892 959540
rect 42116 959500 42892 959528
rect 42116 959488 42122 959500
rect 42886 959488 42892 959500
rect 42944 959488 42950 959540
rect 42150 959080 42156 959132
rect 42208 959120 42214 959132
rect 43346 959120 43352 959132
rect 42208 959092 43352 959120
rect 42208 959080 42214 959092
rect 43346 959080 43352 959092
rect 43404 959080 43410 959132
rect 674650 958808 674656 958860
rect 674708 958848 674714 958860
rect 675386 958848 675392 958860
rect 674708 958820 675392 958848
rect 674708 958808 674714 958820
rect 675386 958808 675392 958820
rect 675444 958808 675450 958860
rect 42058 958332 42064 958384
rect 42116 958372 42122 958384
rect 43162 958372 43168 958384
rect 42116 958344 43168 958372
rect 42116 958332 42122 958344
rect 43162 958332 43168 958344
rect 43220 958332 43226 958384
rect 674282 958332 674288 958384
rect 674340 958372 674346 958384
rect 675386 958372 675392 958384
rect 674340 958344 675392 958372
rect 674340 958332 674346 958344
rect 675386 958332 675392 958344
rect 675444 958332 675450 958384
rect 42058 957720 42064 957772
rect 42116 957760 42122 957772
rect 43254 957760 43260 957772
rect 42116 957732 43260 957760
rect 42116 957720 42122 957732
rect 43254 957720 43260 957732
rect 43312 957720 43318 957772
rect 674374 957720 674380 957772
rect 674432 957760 674438 957772
rect 675478 957760 675484 957772
rect 674432 957732 675484 957760
rect 674432 957720 674438 957732
rect 675478 957720 675484 957732
rect 675536 957720 675542 957772
rect 674558 956972 674564 957024
rect 674616 957012 674622 957024
rect 675386 957012 675392 957024
rect 674616 956984 675392 957012
rect 674616 956972 674622 956984
rect 675386 956972 675392 956984
rect 675444 956972 675450 957024
rect 674466 955680 674472 955732
rect 674524 955720 674530 955732
rect 675478 955720 675484 955732
rect 674524 955692 675484 955720
rect 674524 955680 674530 955692
rect 675478 955680 675484 955692
rect 675536 955680 675542 955732
rect 675018 955476 675024 955528
rect 675076 955516 675082 955528
rect 675478 955516 675484 955528
rect 675076 955488 675484 955516
rect 675076 955476 675082 955488
rect 675478 955476 675484 955488
rect 675536 955476 675542 955528
rect 42150 955340 42156 955392
rect 42208 955380 42214 955392
rect 42702 955380 42708 955392
rect 42208 955352 42708 955380
rect 42208 955340 42214 955352
rect 42702 955340 42708 955352
rect 42760 955340 42766 955392
rect 674006 953980 674012 954032
rect 674064 954020 674070 954032
rect 674742 954020 674748 954032
rect 674064 953992 674748 954020
rect 674064 953980 674070 953992
rect 674742 953980 674748 953992
rect 674800 953980 674806 954032
rect 674742 953844 674748 953896
rect 674800 953884 674806 953896
rect 675386 953884 675392 953896
rect 674800 953856 675392 953884
rect 674800 953844 674806 953856
rect 675386 953844 675392 953856
rect 675444 953844 675450 953896
rect 674834 952144 674840 952196
rect 674892 952184 674898 952196
rect 674892 952156 675708 952184
rect 674892 952144 674898 952156
rect 674834 952008 674840 952060
rect 674892 952048 674898 952060
rect 675386 952048 675392 952060
rect 674892 952020 675392 952048
rect 674892 952008 674898 952020
rect 675386 952008 675392 952020
rect 675444 952008 675450 952060
rect 675680 951788 675708 952156
rect 675662 951736 675668 951788
rect 675720 951736 675726 951788
rect 674006 951056 674012 951108
rect 674064 951096 674070 951108
rect 675754 951096 675760 951108
rect 674064 951068 675760 951096
rect 674064 951056 674070 951068
rect 675754 951056 675760 951068
rect 675812 951056 675818 951108
rect 673730 950920 673736 950972
rect 673788 950960 673794 950972
rect 674006 950960 674012 950972
rect 673788 950932 674012 950960
rect 673788 950920 673794 950932
rect 674006 950920 674012 950932
rect 674064 950920 674070 950972
rect 673454 950716 673460 950768
rect 673512 950756 673518 950768
rect 673638 950756 673644 950768
rect 673512 950728 673644 950756
rect 673512 950716 673518 950728
rect 673638 950716 673644 950728
rect 673696 950716 673702 950768
rect 35618 949560 35624 949612
rect 35676 949600 35682 949612
rect 43622 949600 43628 949612
rect 35676 949572 43628 949600
rect 35676 949560 35682 949572
rect 43622 949560 43628 949572
rect 43680 949560 43686 949612
rect 35710 949492 35716 949544
rect 35768 949532 35774 949544
rect 42886 949532 42892 949544
rect 35768 949504 42892 949532
rect 35768 949492 35774 949504
rect 42886 949492 42892 949504
rect 42944 949492 42950 949544
rect 41506 949424 41512 949476
rect 41564 949464 41570 949476
rect 58434 949464 58440 949476
rect 41564 949436 58440 949464
rect 41564 949424 41570 949436
rect 58434 949424 58440 949436
rect 58492 949424 58498 949476
rect 41966 943236 41972 943288
rect 42024 943276 42030 943288
rect 62666 943276 62672 943288
rect 42024 943248 62672 943276
rect 42024 943236 42030 943248
rect 62666 943236 62672 943248
rect 62724 943236 62730 943288
rect 41782 943032 41788 943084
rect 41840 943072 41846 943084
rect 49694 943072 49700 943084
rect 41840 943044 49700 943072
rect 41840 943032 41846 943044
rect 49694 943032 49700 943044
rect 49752 943032 49758 943084
rect 703446 942896 703452 942948
rect 703504 942936 703510 942948
rect 709334 942936 709340 942948
rect 703504 942908 709340 942936
rect 703504 942896 703510 942908
rect 709334 942896 709340 942908
rect 709392 942896 709398 942948
rect 41782 942692 41788 942744
rect 41840 942732 41846 942744
rect 48498 942732 48504 942744
rect 41840 942704 48504 942732
rect 41840 942692 41846 942704
rect 48498 942692 48504 942704
rect 48556 942692 48562 942744
rect 41782 941468 41788 941520
rect 41840 941508 41846 941520
rect 46014 941508 46020 941520
rect 41840 941480 46020 941508
rect 41840 941468 41846 941480
rect 46014 941468 46020 941480
rect 46072 941468 46078 941520
rect 41782 941332 41788 941384
rect 41840 941372 41846 941384
rect 42702 941372 42708 941384
rect 41840 941344 42708 941372
rect 41840 941332 41846 941344
rect 42702 941332 42708 941344
rect 42760 941332 42766 941384
rect 41874 941196 41880 941248
rect 41932 941236 41938 941248
rect 42702 941236 42708 941248
rect 41932 941208 42708 941236
rect 41932 941196 41938 941208
rect 42702 941196 42708 941208
rect 42760 941196 42766 941248
rect 703538 940856 703544 940908
rect 703596 940896 703602 940908
rect 708874 940896 708880 940908
rect 703596 940868 708880 940896
rect 703596 940856 703602 940868
rect 708874 940856 708880 940868
rect 708932 940856 708938 940908
rect 708046 940828 708052 940840
rect 704844 940800 708052 940828
rect 704844 940704 704872 940800
rect 708046 940788 708052 940800
rect 708104 940788 708110 940840
rect 704918 940720 704924 940772
rect 704976 940760 704982 940772
rect 707954 940760 707960 940772
rect 704976 940732 707960 940760
rect 704976 940720 704982 940732
rect 707954 940720 707960 940732
rect 708012 940720 708018 940772
rect 704826 940652 704832 940704
rect 704884 940652 704890 940704
rect 707034 940692 707040 940704
rect 705764 940664 707040 940692
rect 705764 940568 705792 940664
rect 707034 940652 707040 940664
rect 707092 940652 707098 940704
rect 706666 940624 706672 940636
rect 706224 940596 706672 940624
rect 706224 940568 706252 940596
rect 706666 940584 706672 940596
rect 706724 940584 706730 940636
rect 705746 940516 705752 940568
rect 705804 940516 705810 940568
rect 706206 940516 706212 940568
rect 706264 940516 706270 940568
rect 706298 940516 706304 940568
rect 706356 940556 706362 940568
rect 706574 940556 706580 940568
rect 706356 940528 706580 940556
rect 706356 940516 706362 940528
rect 706574 940516 706580 940528
rect 706632 940516 706638 940568
rect 705838 940448 705844 940500
rect 705896 940488 705902 940500
rect 707034 940488 707040 940500
rect 705896 940460 707040 940488
rect 705896 940448 705902 940460
rect 707034 940448 707040 940460
rect 707092 940448 707098 940500
rect 707586 940448 707592 940500
rect 707644 940448 707650 940500
rect 705378 940380 705384 940432
rect 705436 940420 705442 940432
rect 707494 940420 707500 940432
rect 705436 940392 707500 940420
rect 705436 940380 705442 940392
rect 707494 940380 707500 940392
rect 707552 940380 707558 940432
rect 705286 940312 705292 940364
rect 705344 940352 705350 940364
rect 707604 940352 707632 940448
rect 705344 940324 707632 940352
rect 705344 940312 705350 940324
rect 708506 940312 708512 940364
rect 708564 940312 708570 940364
rect 704458 940244 704464 940296
rect 704516 940284 704522 940296
rect 708414 940284 708420 940296
rect 704516 940256 708420 940284
rect 704516 940244 704522 940256
rect 708414 940244 708420 940256
rect 708472 940244 708478 940296
rect 704366 940176 704372 940228
rect 704424 940216 704430 940228
rect 708524 940216 708552 940312
rect 704424 940188 708552 940216
rect 704424 940176 704430 940188
rect 655790 938816 655796 938868
rect 655848 938856 655854 938868
rect 676214 938856 676220 938868
rect 655848 938828 676220 938856
rect 655848 938816 655854 938828
rect 676214 938816 676220 938828
rect 676272 938816 676278 938868
rect 655698 938680 655704 938732
rect 655756 938720 655762 938732
rect 676306 938720 676312 938732
rect 655756 938692 676312 938720
rect 655756 938680 655762 938692
rect 676306 938680 676312 938692
rect 676364 938680 676370 938732
rect 655514 938544 655520 938596
rect 655572 938584 655578 938596
rect 676122 938584 676128 938596
rect 655572 938556 676128 938584
rect 655572 938544 655578 938556
rect 676122 938544 676128 938556
rect 676180 938544 676186 938596
rect 49694 938340 49700 938392
rect 49752 938380 49758 938392
rect 58434 938380 58440 938392
rect 49752 938352 58440 938380
rect 49752 938340 49758 938352
rect 58434 938340 58440 938352
rect 58492 938340 58498 938392
rect 41138 936504 41144 936556
rect 41196 936544 41202 936556
rect 41690 936544 41696 936556
rect 41196 936516 41696 936544
rect 41196 936504 41202 936516
rect 41690 936504 41696 936516
rect 41748 936504 41754 936556
rect 670326 935756 670332 935808
rect 670384 935796 670390 935808
rect 676030 935796 676036 935808
rect 670384 935768 676036 935796
rect 670384 935756 670390 935768
rect 676030 935756 676036 935768
rect 676088 935756 676094 935808
rect 670142 935688 670148 935740
rect 670200 935728 670206 935740
rect 676214 935728 676220 935740
rect 670200 935700 676220 935728
rect 670200 935688 670206 935700
rect 676214 935688 676220 935700
rect 676272 935688 676278 935740
rect 649902 935620 649908 935672
rect 649960 935660 649966 935672
rect 678974 935660 678980 935672
rect 649960 935632 678980 935660
rect 649960 935620 649966 935632
rect 678974 935620 678980 935632
rect 679032 935620 679038 935672
rect 674742 935552 674748 935604
rect 674800 935592 674806 935604
rect 676030 935592 676036 935604
rect 674800 935564 676036 935592
rect 674800 935552 674806 935564
rect 676030 935552 676036 935564
rect 676088 935552 676094 935604
rect 674650 935484 674656 935536
rect 674708 935524 674714 935536
rect 676122 935524 676128 935536
rect 674708 935496 676128 935524
rect 674708 935484 674714 935496
rect 676122 935484 676128 935496
rect 676180 935484 676186 935536
rect 674006 935416 674012 935468
rect 674064 935456 674070 935468
rect 675938 935456 675944 935468
rect 674064 935428 675944 935456
rect 674064 935416 674070 935428
rect 675938 935416 675944 935428
rect 675996 935416 676002 935468
rect 673914 935280 673920 935332
rect 673972 935320 673978 935332
rect 675938 935320 675944 935332
rect 673972 935292 675944 935320
rect 673972 935280 673978 935292
rect 675938 935280 675944 935292
rect 675996 935280 676002 935332
rect 674834 934940 674840 934992
rect 674892 934980 674898 934992
rect 676030 934980 676036 934992
rect 674892 934952 676036 934980
rect 674892 934940 674898 934952
rect 676030 934940 676036 934952
rect 676088 934940 676094 934992
rect 673546 933308 673552 933360
rect 673604 933348 673610 933360
rect 676030 933348 676036 933360
rect 673604 933320 676036 933348
rect 673604 933308 673610 933320
rect 676030 933308 676036 933320
rect 676088 933308 676094 933360
rect 674466 932832 674472 932884
rect 674524 932872 674530 932884
rect 676030 932872 676036 932884
rect 674524 932844 676036 932872
rect 674524 932832 674530 932844
rect 676030 932832 676036 932844
rect 676088 932832 676094 932884
rect 673730 932764 673736 932816
rect 673788 932804 673794 932816
rect 676122 932804 676128 932816
rect 673788 932776 676128 932804
rect 673788 932764 673794 932776
rect 676122 932764 676128 932776
rect 676180 932764 676186 932816
rect 673638 932696 673644 932748
rect 673696 932736 673702 932748
rect 675938 932736 675944 932748
rect 673696 932708 675944 932736
rect 673696 932696 673702 932708
rect 675938 932696 675944 932708
rect 675996 932696 676002 932748
rect 674282 932628 674288 932680
rect 674340 932668 674346 932680
rect 676122 932668 676128 932680
rect 674340 932640 676128 932668
rect 674340 932628 674346 932640
rect 676122 932628 676128 932640
rect 676180 932628 676186 932680
rect 41782 932424 41788 932476
rect 41840 932464 41846 932476
rect 46014 932464 46020 932476
rect 41840 932436 46020 932464
rect 41840 932424 41846 932436
rect 46014 932424 46020 932436
rect 46072 932424 46078 932476
rect 673822 932084 673828 932136
rect 673880 932124 673886 932136
rect 675938 932124 675944 932136
rect 673880 932096 675944 932124
rect 673880 932084 673886 932096
rect 675938 932084 675944 932096
rect 675996 932084 676002 932136
rect 674374 931676 674380 931728
rect 674432 931716 674438 931728
rect 676030 931716 676036 931728
rect 674432 931688 676036 931716
rect 674432 931676 674438 931688
rect 676030 931676 676036 931688
rect 676088 931676 676094 931728
rect 674558 931268 674564 931320
rect 674616 931308 674622 931320
rect 676030 931308 676036 931320
rect 674616 931280 676036 931308
rect 674616 931268 674622 931280
rect 676030 931268 676036 931280
rect 676088 931268 676094 931320
rect 672074 927392 672080 927444
rect 672132 927432 672138 927444
rect 678974 927432 678980 927444
rect 672132 927404 678980 927432
rect 672132 927392 672138 927404
rect 678974 927392 678980 927404
rect 679032 927392 679038 927444
rect 654686 922224 654692 922276
rect 654744 922264 654750 922276
rect 669866 922264 669872 922276
rect 654744 922236 669872 922264
rect 654744 922224 654750 922236
rect 669866 922224 669872 922236
rect 669924 922224 669930 922276
rect 48498 921816 48504 921868
rect 48556 921856 48562 921868
rect 58434 921856 58440 921868
rect 48556 921828 58440 921856
rect 48556 921816 48562 921828
rect 58434 921816 58440 921828
rect 58492 921816 58498 921868
rect 53834 908080 53840 908132
rect 53892 908120 53898 908132
rect 58066 908120 58072 908132
rect 53892 908092 58072 908120
rect 53892 908080 53898 908092
rect 58066 908080 58072 908092
rect 58124 908080 58130 908132
rect 654870 908080 654876 908132
rect 654928 908120 654934 908132
rect 663794 908120 663800 908132
rect 654928 908092 663800 908120
rect 654928 908080 654934 908092
rect 663794 908080 663800 908092
rect 663852 908080 663858 908132
rect 53926 896996 53932 897048
rect 53984 897036 53990 897048
rect 58526 897036 58532 897048
rect 53984 897008 58532 897036
rect 53984 896996 53990 897008
rect 58526 896996 58532 897008
rect 58584 896996 58590 897048
rect 654686 895364 654692 895416
rect 654744 895404 654750 895416
rect 660942 895404 660948 895416
rect 654744 895376 660948 895404
rect 654744 895364 654750 895376
rect 660942 895364 660948 895376
rect 661000 895364 661006 895416
rect 51074 883192 51080 883244
rect 51132 883232 51138 883244
rect 58434 883232 58440 883244
rect 51132 883204 58440 883232
rect 51132 883192 51138 883204
rect 58434 883192 58440 883204
rect 58492 883192 58498 883244
rect 673546 873468 673552 873520
rect 673604 873508 673610 873520
rect 675386 873508 675392 873520
rect 673604 873480 675392 873508
rect 673604 873468 673610 873480
rect 675386 873468 675392 873480
rect 675444 873468 675450 873520
rect 674742 872652 674748 872704
rect 674800 872692 674806 872704
rect 675386 872692 675392 872704
rect 674800 872664 675392 872692
rect 674800 872652 674806 872664
rect 675386 872652 675392 872664
rect 675444 872652 675450 872704
rect 655146 870748 655152 870800
rect 655204 870788 655210 870800
rect 674926 870788 674932 870800
rect 655204 870760 674932 870788
rect 655204 870748 655210 870760
rect 674926 870748 674932 870760
rect 674984 870748 674990 870800
rect 673638 869796 673644 869848
rect 673696 869836 673702 869848
rect 675386 869836 675392 869848
rect 673696 869808 675392 869836
rect 673696 869796 673702 869808
rect 675386 869796 675392 869808
rect 675444 869796 675450 869848
rect 656802 869592 656808 869644
rect 656860 869632 656866 869644
rect 663702 869632 663708 869644
rect 656860 869604 663708 869632
rect 656860 869592 656866 869604
rect 663702 869592 663708 869604
rect 663760 869592 663766 869644
rect 50982 869388 50988 869440
rect 51040 869428 51046 869440
rect 58434 869428 58440 869440
rect 51040 869400 58440 869428
rect 51040 869388 51046 869400
rect 58434 869388 58440 869400
rect 58492 869388 58498 869440
rect 674190 868980 674196 869032
rect 674248 869020 674254 869032
rect 675386 869020 675392 869032
rect 674248 868992 675392 869020
rect 674248 868980 674254 868992
rect 675386 868980 675392 868992
rect 675444 868980 675450 869032
rect 673730 868504 673736 868556
rect 673788 868544 673794 868556
rect 675386 868544 675392 868556
rect 673788 868516 675392 868544
rect 673788 868504 673794 868516
rect 675386 868504 675392 868516
rect 675444 868504 675450 868556
rect 674282 867756 674288 867808
rect 674340 867796 674346 867808
rect 675386 867796 675392 867808
rect 674340 867768 675392 867796
rect 674340 867756 674346 867768
rect 675386 867756 675392 867768
rect 675444 867756 675450 867808
rect 673822 866464 673828 866516
rect 673880 866504 673886 866516
rect 675386 866504 675392 866516
rect 673880 866476 675392 866504
rect 673880 866464 673886 866476
rect 675386 866464 675392 866476
rect 675444 866464 675450 866516
rect 674926 866260 674932 866312
rect 674984 866300 674990 866312
rect 675386 866300 675392 866312
rect 674984 866272 675392 866300
rect 674984 866260 674990 866272
rect 675386 866260 675392 866272
rect 675444 866260 675450 866312
rect 674006 864628 674012 864680
rect 674064 864668 674070 864680
rect 675386 864668 675392 864680
rect 674064 864640 675392 864668
rect 674064 864628 674070 864640
rect 675386 864628 675392 864640
rect 675444 864628 675450 864680
rect 673914 862792 673920 862844
rect 673972 862832 673978 862844
rect 675478 862832 675484 862844
rect 673972 862804 675484 862832
rect 673972 862792 673978 862804
rect 675478 862792 675484 862804
rect 675536 862792 675542 862844
rect 48590 858372 48596 858424
rect 48648 858412 48654 858424
rect 58434 858412 58440 858424
rect 48648 858384 58440 858412
rect 48648 858372 48654 858384
rect 58434 858372 58440 858384
rect 58492 858372 58498 858424
rect 655238 855584 655244 855636
rect 655296 855624 655302 855636
rect 666462 855624 666468 855636
rect 655296 855596 666468 855624
rect 655296 855584 655302 855596
rect 666462 855584 666468 855596
rect 666520 855584 666526 855636
rect 674742 854224 674748 854276
rect 674800 854264 674806 854276
rect 675570 854264 675576 854276
rect 674800 854236 675576 854264
rect 674800 854224 674806 854236
rect 675570 854224 675576 854236
rect 675628 854224 675634 854276
rect 48682 844568 48688 844620
rect 48740 844608 48746 844620
rect 58434 844608 58440 844620
rect 48740 844580 58440 844608
rect 48740 844568 48746 844580
rect 58434 844568 58440 844580
rect 58492 844568 58498 844620
rect 654870 841780 654876 841832
rect 654928 841820 654934 841832
rect 667106 841820 667112 841832
rect 654928 841792 667112 841820
rect 654928 841780 654934 841792
rect 667106 841780 667112 841792
rect 667164 841780 667170 841832
rect 54018 830764 54024 830816
rect 54076 830804 54082 830816
rect 57974 830804 57980 830816
rect 54076 830776 57980 830804
rect 54076 830764 54082 830776
rect 57974 830764 57980 830776
rect 58032 830764 58038 830816
rect 41138 819748 41144 819800
rect 41196 819788 41202 819800
rect 62298 819788 62304 819800
rect 41196 819760 62304 819788
rect 41196 819748 41202 819760
rect 62298 819748 62304 819760
rect 62356 819748 62362 819800
rect 41782 817436 41788 817488
rect 41840 817476 41846 817488
rect 53926 817476 53932 817488
rect 41840 817448 53932 817476
rect 41840 817436 41846 817448
rect 53926 817436 53932 817448
rect 53984 817436 53990 817488
rect 41782 817300 41788 817352
rect 41840 817340 41846 817352
rect 51074 817340 51080 817352
rect 41840 817312 51080 817340
rect 41840 817300 41846 817312
rect 51074 817300 51080 817312
rect 51132 817300 51138 817352
rect 53742 817028 53748 817080
rect 53800 817068 53806 817080
rect 59170 817068 59176 817080
rect 53800 817040 59176 817068
rect 53800 817028 53806 817040
rect 59170 817028 59176 817040
rect 59228 817028 59234 817080
rect 42702 816960 42708 817012
rect 42760 817000 42766 817012
rect 62482 817000 62488 817012
rect 42760 816972 62488 817000
rect 42760 816960 42766 816972
rect 62482 816960 62488 816972
rect 62540 816960 62546 817012
rect 655054 815600 655060 815652
rect 655112 815640 655118 815652
rect 668946 815640 668952 815652
rect 655112 815612 668952 815640
rect 655112 815600 655118 815612
rect 668946 815600 668952 815612
rect 669004 815600 669010 815652
rect 41782 814240 41788 814292
rect 41840 814280 41846 814292
rect 42886 814280 42892 814292
rect 41840 814252 42892 814280
rect 41840 814240 41846 814252
rect 42886 814240 42892 814252
rect 42944 814280 42950 814292
rect 62666 814280 62672 814292
rect 42944 814252 62672 814280
rect 42944 814240 42950 814252
rect 62666 814240 62672 814252
rect 62724 814240 62730 814292
rect 41782 810024 41788 810076
rect 41840 810064 41846 810076
rect 43714 810064 43720 810076
rect 41840 810036 43720 810064
rect 41840 810024 41846 810036
rect 43714 810024 43720 810036
rect 43772 810024 43778 810076
rect 41874 807848 41880 807900
rect 41932 807888 41938 807900
rect 43162 807888 43168 807900
rect 41932 807860 43168 807888
rect 41932 807848 41938 807860
rect 43162 807848 43168 807860
rect 43220 807848 43226 807900
rect 41782 807576 41788 807628
rect 41840 807616 41846 807628
rect 42702 807616 42708 807628
rect 41840 807588 42708 807616
rect 41840 807576 41846 807588
rect 42702 807576 42708 807588
rect 42760 807576 42766 807628
rect 41782 806624 41788 806676
rect 41840 806664 41846 806676
rect 46290 806664 46296 806676
rect 41840 806636 46296 806664
rect 41840 806624 41846 806636
rect 46290 806624 46296 806636
rect 46348 806624 46354 806676
rect 51074 805944 51080 805996
rect 51132 805984 51138 805996
rect 58434 805984 58440 805996
rect 51132 805956 58440 805984
rect 51132 805944 51138 805956
rect 58434 805944 58440 805956
rect 58492 805944 58498 805996
rect 656158 803224 656164 803276
rect 656216 803264 656222 803276
rect 661034 803264 661040 803276
rect 656216 803236 661040 803264
rect 656216 803224 656222 803236
rect 661034 803224 661040 803236
rect 661092 803224 661098 803276
rect 44266 800436 44272 800488
rect 44324 800476 44330 800488
rect 48498 800476 48504 800488
rect 44324 800448 48504 800476
rect 44324 800436 44330 800448
rect 48498 800436 48504 800448
rect 48556 800436 48562 800488
rect 41966 800164 41972 800216
rect 42024 800164 42030 800216
rect 41984 800012 42012 800164
rect 41966 799960 41972 800012
rect 42024 799960 42030 800012
rect 43806 799756 43812 799808
rect 43864 799796 43870 799808
rect 44082 799796 44088 799808
rect 43864 799768 44088 799796
rect 43864 799756 43870 799768
rect 44082 799756 44088 799768
rect 44140 799756 44146 799808
rect 42334 799688 42340 799740
rect 42392 799728 42398 799740
rect 42392 799700 43852 799728
rect 42392 799688 42398 799700
rect 43824 799672 43852 799700
rect 43806 799620 43812 799672
rect 43864 799620 43870 799672
rect 42150 798124 42156 798176
rect 42208 798164 42214 798176
rect 42886 798164 42892 798176
rect 42208 798136 42892 798164
rect 42208 798124 42214 798136
rect 42886 798124 42892 798136
rect 42944 798124 42950 798176
rect 43806 798164 43812 798176
rect 43732 798136 43812 798164
rect 42702 797920 42708 797972
rect 42760 797920 42766 797972
rect 43438 797920 43444 797972
rect 43496 797920 43502 797972
rect 42426 797580 42432 797632
rect 42484 797620 42490 797632
rect 42720 797620 42748 797920
rect 42978 797852 42984 797904
rect 43036 797892 43042 797904
rect 43456 797892 43484 797920
rect 43036 797864 43484 797892
rect 43036 797852 43042 797864
rect 43530 797648 43536 797700
rect 43588 797688 43594 797700
rect 43732 797688 43760 798136
rect 43806 798124 43812 798136
rect 43864 798124 43870 798176
rect 43806 797988 43812 798040
rect 43864 798028 43870 798040
rect 44174 798028 44180 798040
rect 43864 798000 44180 798028
rect 43864 797988 43870 798000
rect 44174 797988 44180 798000
rect 44232 797988 44238 798040
rect 43588 797660 43760 797688
rect 43588 797648 43594 797660
rect 42484 797592 42748 797620
rect 42484 797580 42490 797592
rect 42150 797240 42156 797292
rect 42208 797280 42214 797292
rect 44266 797280 44272 797292
rect 42208 797252 44272 797280
rect 42208 797240 42214 797252
rect 44266 797240 44272 797252
rect 44324 797240 44330 797292
rect 42150 796288 42156 796340
rect 42208 796328 42214 796340
rect 42702 796328 42708 796340
rect 42208 796300 42708 796328
rect 42208 796288 42214 796300
rect 42702 796288 42708 796300
rect 42760 796288 42766 796340
rect 674558 796220 674564 796272
rect 674616 796260 674622 796272
rect 675570 796260 675576 796272
rect 674616 796232 675576 796260
rect 674616 796220 674622 796232
rect 675570 796220 675576 796232
rect 675628 796220 675634 796272
rect 42150 794996 42156 795048
rect 42208 795036 42214 795048
rect 43162 795036 43168 795048
rect 42208 795008 43168 795036
rect 42208 794996 42214 795008
rect 43162 794996 43168 795008
rect 43220 794996 43226 795048
rect 42150 794248 42156 794300
rect 42208 794288 42214 794300
rect 43254 794288 43260 794300
rect 42208 794260 43260 794288
rect 42208 794248 42214 794260
rect 43254 794248 43260 794260
rect 43312 794248 43318 794300
rect 42150 793772 42156 793824
rect 42208 793812 42214 793824
rect 42426 793812 42432 793824
rect 42208 793784 42432 793812
rect 42208 793772 42214 793784
rect 42426 793772 42432 793784
rect 42484 793772 42490 793824
rect 42150 792956 42156 793008
rect 42208 792996 42214 793008
rect 43714 792996 43720 793008
rect 42208 792968 43720 792996
rect 42208 792956 42214 792968
rect 43714 792956 43720 792968
rect 43772 792956 43778 793008
rect 51166 792140 51172 792192
rect 51224 792180 51230 792192
rect 58066 792180 58072 792192
rect 51224 792152 58072 792180
rect 51224 792140 51230 792152
rect 58066 792140 58072 792152
rect 58124 792140 58130 792192
rect 42150 790644 42156 790696
rect 42208 790684 42214 790696
rect 43622 790684 43628 790696
rect 42208 790656 43628 790684
rect 42208 790644 42214 790656
rect 43622 790644 43628 790656
rect 43680 790644 43686 790696
rect 42150 790100 42156 790152
rect 42208 790140 42214 790152
rect 43898 790140 43904 790152
rect 42208 790112 43904 790140
rect 42208 790100 42214 790112
rect 43898 790100 43904 790112
rect 43956 790100 43962 790152
rect 655054 789352 655060 789404
rect 655112 789392 655118 789404
rect 663886 789392 663892 789404
rect 655112 789364 663892 789392
rect 655112 789352 655118 789364
rect 663886 789352 663892 789364
rect 663944 789352 663950 789404
rect 42150 789284 42156 789336
rect 42208 789324 42214 789336
rect 43806 789324 43812 789336
rect 42208 789296 43812 789324
rect 42208 789284 42214 789296
rect 43806 789284 43812 789296
rect 43864 789284 43870 789336
rect 42150 788808 42156 788860
rect 42208 788848 42214 788860
rect 43070 788848 43076 788860
rect 42208 788820 43076 788848
rect 42208 788808 42214 788820
rect 43070 788808 43076 788820
rect 43128 788808 43134 788860
rect 42150 786972 42156 787024
rect 42208 787012 42214 787024
rect 43346 787012 43352 787024
rect 42208 786984 43352 787012
rect 42208 786972 42214 786984
rect 43346 786972 43352 786984
rect 43404 786972 43410 787024
rect 42058 786224 42064 786276
rect 42116 786264 42122 786276
rect 44082 786264 44088 786276
rect 42116 786236 44088 786264
rect 42116 786224 42122 786236
rect 44082 786224 44088 786236
rect 44140 786224 44146 786276
rect 42150 785748 42156 785800
rect 42208 785788 42214 785800
rect 42886 785788 42892 785800
rect 42208 785760 42892 785788
rect 42208 785748 42214 785760
rect 42886 785748 42892 785760
rect 42944 785748 42950 785800
rect 674374 784932 674380 784984
rect 674432 784972 674438 784984
rect 675386 784972 675392 784984
rect 674432 784944 675392 784972
rect 674432 784932 674438 784944
rect 675386 784932 675392 784944
rect 675444 784932 675450 784984
rect 673454 782892 673460 782944
rect 673512 782932 673518 782944
rect 675478 782932 675484 782944
rect 673512 782904 675484 782932
rect 673512 782892 673518 782904
rect 675478 782892 675484 782904
rect 675536 782892 675542 782944
rect 655514 782416 655520 782468
rect 655572 782456 655578 782468
rect 674650 782456 674656 782468
rect 655572 782428 674656 782456
rect 655572 782416 655578 782428
rect 674650 782416 674656 782428
rect 674708 782416 674714 782468
rect 674282 780580 674288 780632
rect 674340 780620 674346 780632
rect 675478 780620 675484 780632
rect 674340 780592 675484 780620
rect 674340 780580 674346 780592
rect 675478 780580 675484 780592
rect 675536 780580 675542 780632
rect 674466 779764 674472 779816
rect 674524 779804 674530 779816
rect 675478 779804 675484 779816
rect 674524 779776 675484 779804
rect 674524 779764 674530 779776
rect 675478 779764 675484 779776
rect 675536 779764 675542 779816
rect 674190 779288 674196 779340
rect 674248 779328 674254 779340
rect 675386 779328 675392 779340
rect 674248 779300 675392 779328
rect 674248 779288 674254 779300
rect 675386 779288 675392 779300
rect 675444 779288 675450 779340
rect 674742 778608 674748 778660
rect 674800 778648 674806 778660
rect 675478 778648 675484 778660
rect 674800 778620 675484 778648
rect 674800 778608 674806 778620
rect 675478 778608 675484 778620
rect 675536 778608 675542 778660
rect 48866 778336 48872 778388
rect 48924 778376 48930 778388
rect 58434 778376 58440 778388
rect 48924 778348 58440 778376
rect 48924 778336 48930 778348
rect 58434 778336 58440 778348
rect 58492 778336 58498 778388
rect 674374 777316 674380 777368
rect 674432 777356 674438 777368
rect 675386 777356 675392 777368
rect 674432 777328 675392 777356
rect 674432 777316 674438 777328
rect 675386 777316 675392 777328
rect 675444 777316 675450 777368
rect 674650 777044 674656 777096
rect 674708 777084 674714 777096
rect 675386 777084 675392 777096
rect 674708 777056 675392 777084
rect 674708 777044 674714 777056
rect 675386 777044 675392 777056
rect 675444 777044 675450 777096
rect 674558 775480 674564 775532
rect 674616 775520 674622 775532
rect 675386 775520 675392 775532
rect 674616 775492 675392 775520
rect 674616 775480 674622 775492
rect 675386 775480 675392 775492
rect 675444 775480 675450 775532
rect 41506 774732 41512 774784
rect 41564 774772 41570 774784
rect 48682 774772 48688 774784
rect 41564 774744 48688 774772
rect 41564 774732 41570 774744
rect 48682 774732 48688 774744
rect 48740 774732 48746 774784
rect 41782 774188 41788 774240
rect 41840 774228 41846 774240
rect 54018 774228 54024 774240
rect 41840 774200 54024 774228
rect 41840 774188 41846 774200
rect 54018 774188 54024 774200
rect 54076 774188 54082 774240
rect 41506 773916 41512 773968
rect 41564 773956 41570 773968
rect 48590 773956 48596 773968
rect 41564 773928 48596 773956
rect 41564 773916 41570 773928
rect 48590 773916 48596 773928
rect 48648 773916 48654 773968
rect 674650 773848 674656 773900
rect 674708 773888 674714 773900
rect 675202 773888 675208 773900
rect 674708 773860 675208 773888
rect 674708 773848 674714 773860
rect 675202 773848 675208 773860
rect 675260 773848 675266 773900
rect 41506 773576 41512 773628
rect 41564 773616 41570 773628
rect 43346 773616 43352 773628
rect 41564 773588 43352 773616
rect 41564 773576 41570 773588
rect 43346 773576 43352 773588
rect 43404 773616 43410 773628
rect 43990 773616 43996 773628
rect 43404 773588 43996 773616
rect 43404 773576 43410 773588
rect 43990 773576 43996 773588
rect 44048 773576 44054 773628
rect 674650 773576 674656 773628
rect 674708 773616 674714 773628
rect 675478 773616 675484 773628
rect 674708 773588 675484 773616
rect 674708 773576 674714 773588
rect 675478 773576 675484 773588
rect 675536 773576 675542 773628
rect 674466 773372 674472 773424
rect 674524 773412 674530 773424
rect 675662 773412 675668 773424
rect 674524 773384 675668 773412
rect 674524 773372 674530 773384
rect 675662 773372 675668 773384
rect 675720 773372 675726 773424
rect 675202 773304 675208 773356
rect 675260 773344 675266 773356
rect 675570 773344 675576 773356
rect 675260 773316 675576 773344
rect 675260 773304 675266 773316
rect 675570 773304 675576 773316
rect 675628 773304 675634 773356
rect 674742 773100 674748 773152
rect 674800 773140 674806 773152
rect 675478 773140 675484 773152
rect 674800 773112 675484 773140
rect 674800 773100 674806 773112
rect 675478 773100 675484 773112
rect 675536 773100 675542 773152
rect 42886 772828 42892 772880
rect 42944 772868 42950 772880
rect 62850 772868 62856 772880
rect 42944 772840 62856 772868
rect 42944 772828 42950 772840
rect 62850 772828 62856 772840
rect 62908 772828 62914 772880
rect 674282 770516 674288 770568
rect 674340 770556 674346 770568
rect 674558 770556 674564 770568
rect 674340 770528 674564 770556
rect 674340 770516 674346 770528
rect 674558 770516 674564 770528
rect 674616 770516 674622 770568
rect 673454 770244 673460 770296
rect 673512 770284 673518 770296
rect 674282 770284 674288 770296
rect 673512 770256 674288 770284
rect 673512 770244 673518 770256
rect 674282 770244 674288 770256
rect 674340 770244 674346 770296
rect 48774 767320 48780 767372
rect 48832 767360 48838 767372
rect 58434 767360 58440 767372
rect 48832 767332 58440 767360
rect 48832 767320 48838 767332
rect 58434 767320 58440 767332
rect 58492 767320 58498 767372
rect 43162 766368 43168 766420
rect 43220 766408 43226 766420
rect 43806 766408 43812 766420
rect 43220 766380 43812 766408
rect 43220 766368 43226 766380
rect 43806 766368 43812 766380
rect 43864 766368 43870 766420
rect 41506 763240 41512 763292
rect 41564 763280 41570 763292
rect 48498 763280 48504 763292
rect 41564 763252 48504 763280
rect 41564 763240 41570 763252
rect 48498 763240 48504 763252
rect 48556 763240 48562 763292
rect 708506 762532 708512 762544
rect 704384 762504 708512 762532
rect 704384 762408 704412 762504
rect 708506 762492 708512 762504
rect 708564 762492 708570 762544
rect 704458 762424 704464 762476
rect 704516 762464 704522 762476
rect 708414 762464 708420 762476
rect 704516 762436 708420 762464
rect 704516 762424 704522 762436
rect 708414 762424 708420 762436
rect 708472 762424 708478 762476
rect 704366 762356 704372 762408
rect 704424 762356 704430 762408
rect 707494 762396 707500 762408
rect 705304 762368 707500 762396
rect 705304 762272 705332 762368
rect 707494 762356 707500 762368
rect 707552 762356 707558 762408
rect 707034 762328 707040 762340
rect 705764 762300 707040 762328
rect 705764 762272 705792 762300
rect 707034 762288 707040 762300
rect 707092 762288 707098 762340
rect 705286 762220 705292 762272
rect 705344 762220 705350 762272
rect 705746 762220 705752 762272
rect 705804 762220 705810 762272
rect 706206 762220 706212 762272
rect 706264 762260 706270 762272
rect 706574 762260 706580 762272
rect 706264 762232 706580 762260
rect 706264 762220 706270 762232
rect 706574 762220 706580 762232
rect 706632 762220 706638 762272
rect 705838 762152 705844 762204
rect 705896 762192 705902 762204
rect 707034 762192 707040 762204
rect 705896 762164 707040 762192
rect 705896 762152 705902 762164
rect 707034 762152 707040 762164
rect 707092 762152 707098 762204
rect 706298 762084 706304 762136
rect 706356 762124 706362 762136
rect 706574 762124 706580 762136
rect 706356 762096 706580 762124
rect 706356 762084 706362 762096
rect 706574 762084 706580 762096
rect 706632 762084 706638 762136
rect 705378 762016 705384 762068
rect 705436 762056 705442 762068
rect 707494 762056 707500 762068
rect 705436 762028 707500 762056
rect 705436 762016 705442 762028
rect 707494 762016 707500 762028
rect 707552 762016 707558 762068
rect 708046 762016 708052 762068
rect 708104 762016 708110 762068
rect 704918 761948 704924 762000
rect 704976 761988 704982 762000
rect 707954 761988 707960 762000
rect 704976 761960 707960 761988
rect 704976 761948 704982 761960
rect 707954 761948 707960 761960
rect 708012 761948 708018 762000
rect 704826 761880 704832 761932
rect 704884 761920 704890 761932
rect 708064 761920 708092 762016
rect 704884 761892 708092 761920
rect 704884 761880 704890 761892
rect 708966 761880 708972 761932
rect 709024 761880 709030 761932
rect 703538 761812 703544 761864
rect 703596 761852 703602 761864
rect 708874 761852 708880 761864
rect 703596 761824 708880 761852
rect 703596 761812 703602 761824
rect 708874 761812 708880 761824
rect 708932 761812 708938 761864
rect 654686 761744 654692 761796
rect 654744 761784 654750 761796
rect 667014 761784 667020 761796
rect 654744 761756 667020 761784
rect 654744 761744 654750 761756
rect 667014 761744 667020 761756
rect 667072 761744 667078 761796
rect 703998 761744 704004 761796
rect 704056 761784 704062 761796
rect 708984 761784 709012 761880
rect 704056 761756 709012 761784
rect 704056 761744 704062 761756
rect 41966 760520 41972 760572
rect 42024 760560 42030 760572
rect 50982 760560 50988 760572
rect 42024 760532 50988 760560
rect 42024 760520 42030 760532
rect 50982 760520 50988 760532
rect 51040 760520 51046 760572
rect 669866 759568 669872 759620
rect 669924 759608 669930 759620
rect 676214 759608 676220 759620
rect 669924 759580 676220 759608
rect 669924 759568 669930 759580
rect 676214 759568 676220 759580
rect 676272 759568 676278 759620
rect 663794 759432 663800 759484
rect 663852 759472 663858 759484
rect 678974 759472 678980 759484
rect 663852 759444 678980 759472
rect 663852 759432 663858 759444
rect 678974 759432 678980 759444
rect 679032 759432 679038 759484
rect 660942 759296 660948 759348
rect 661000 759336 661006 759348
rect 676122 759336 676128 759348
rect 661000 759308 676128 759336
rect 661000 759296 661006 759308
rect 676122 759296 676128 759308
rect 676180 759296 676186 759348
rect 673362 759092 673368 759144
rect 673420 759132 673426 759144
rect 676030 759132 676036 759144
rect 673420 759104 676036 759132
rect 673420 759092 673426 759104
rect 676030 759092 676036 759104
rect 676088 759092 676094 759144
rect 670510 759024 670516 759076
rect 670568 759064 670574 759076
rect 676306 759064 676312 759076
rect 670568 759036 676312 759064
rect 670568 759024 670574 759036
rect 676306 759024 676312 759036
rect 676364 759024 676370 759076
rect 674006 758956 674012 759008
rect 674064 758996 674070 759008
rect 676030 758996 676036 759008
rect 674064 758968 676036 758996
rect 674064 758956 674070 758968
rect 676030 758956 676036 758968
rect 676088 758956 676094 759008
rect 42426 757596 42432 757648
rect 42484 757636 42490 757648
rect 42978 757636 42984 757648
rect 42484 757608 42984 757636
rect 42484 757596 42490 757608
rect 42978 757596 42984 757608
rect 43036 757596 43042 757648
rect 43254 757596 43260 757648
rect 43312 757636 43318 757648
rect 43622 757636 43628 757648
rect 43312 757608 43628 757636
rect 43312 757596 43318 757608
rect 43622 757596 43628 757608
rect 43680 757596 43686 757648
rect 42150 757460 42156 757512
rect 42208 757500 42214 757512
rect 43254 757500 43260 757512
rect 42208 757472 43260 757500
rect 42208 757460 42214 757472
rect 43254 757460 43260 757472
rect 43312 757460 43318 757512
rect 42058 757392 42064 757444
rect 42116 757432 42122 757444
rect 42426 757432 42432 757444
rect 42116 757404 42432 757432
rect 42116 757392 42122 757404
rect 42426 757392 42432 757404
rect 42484 757392 42490 757444
rect 41874 756984 41880 757036
rect 41932 756984 41938 757036
rect 41892 756764 41920 756984
rect 41874 756712 41880 756764
rect 41932 756712 41938 756764
rect 42702 756508 42708 756560
rect 42760 756548 42766 756560
rect 44174 756548 44180 756560
rect 42760 756520 44180 756548
rect 42760 756508 42766 756520
rect 44174 756508 44180 756520
rect 44232 756508 44238 756560
rect 670602 756440 670608 756492
rect 670660 756480 670666 756492
rect 676122 756480 676128 756492
rect 670660 756452 676128 756480
rect 670660 756440 670666 756452
rect 676122 756440 676128 756452
rect 676180 756440 676186 756492
rect 668578 756372 668584 756424
rect 668636 756412 668642 756424
rect 676214 756412 676220 756424
rect 668636 756384 676220 756412
rect 668636 756372 668642 756384
rect 676214 756372 676220 756384
rect 676272 756372 676278 756424
rect 669958 756304 669964 756356
rect 670016 756344 670022 756356
rect 670326 756344 670332 756356
rect 670016 756316 670332 756344
rect 670016 756304 670022 756316
rect 670326 756304 670332 756316
rect 670384 756344 670390 756356
rect 676306 756344 676312 756356
rect 670384 756316 676312 756344
rect 670384 756304 670390 756316
rect 676306 756304 676312 756316
rect 676364 756304 676370 756356
rect 669866 756236 669872 756288
rect 669924 756276 669930 756288
rect 670142 756276 670148 756288
rect 669924 756248 670148 756276
rect 669924 756236 669930 756248
rect 670142 756236 670148 756248
rect 670200 756276 670206 756288
rect 678974 756276 678980 756288
rect 670200 756248 678980 756276
rect 670200 756236 670206 756248
rect 678974 756236 678980 756248
rect 679032 756236 679038 756288
rect 673914 756168 673920 756220
rect 673972 756208 673978 756220
rect 676030 756208 676036 756220
rect 673972 756180 676036 756208
rect 673972 756168 673978 756180
rect 676030 756168 676036 756180
rect 676088 756168 676094 756220
rect 673638 756100 673644 756152
rect 673696 756140 673702 756152
rect 676122 756140 676128 756152
rect 673696 756112 676128 756140
rect 673696 756100 673702 756112
rect 676122 756100 676128 756112
rect 676180 756100 676186 756152
rect 42426 755488 42432 755540
rect 42484 755528 42490 755540
rect 42484 755500 42748 755528
rect 42484 755488 42490 755500
rect 42720 755324 42748 755500
rect 42628 755296 42748 755324
rect 42628 755268 42656 755296
rect 42610 755216 42616 755268
rect 42668 755216 42674 755268
rect 42150 754876 42156 754928
rect 42208 754916 42214 754928
rect 43070 754916 43076 754928
rect 42208 754888 43076 754916
rect 42208 754876 42214 754888
rect 43070 754876 43076 754888
rect 43128 754876 43134 754928
rect 673546 754876 673552 754928
rect 673604 754916 673610 754928
rect 676030 754916 676036 754928
rect 673604 754888 676036 754916
rect 673604 754876 673610 754888
rect 676030 754876 676036 754888
rect 676088 754876 676094 754928
rect 43070 754740 43076 754792
rect 43128 754780 43134 754792
rect 43990 754780 43996 754792
rect 43128 754752 43996 754780
rect 43128 754740 43134 754752
rect 43990 754740 43996 754752
rect 44048 754740 44054 754792
rect 44082 754672 44088 754724
rect 44140 754672 44146 754724
rect 44100 754520 44128 754672
rect 44082 754468 44088 754520
rect 44140 754468 44146 754520
rect 53834 753516 53840 753568
rect 53892 753556 53898 753568
rect 58342 753556 58348 753568
rect 53892 753528 58348 753556
rect 53892 753516 53898 753528
rect 58342 753516 58348 753528
rect 58400 753516 58406 753568
rect 673822 753448 673828 753500
rect 673880 753488 673886 753500
rect 676030 753488 676036 753500
rect 673880 753460 676036 753488
rect 673880 753448 673886 753460
rect 676030 753448 676036 753460
rect 676088 753448 676094 753500
rect 673730 753244 673736 753296
rect 673788 753284 673794 753296
rect 676030 753284 676036 753296
rect 673788 753256 676036 753284
rect 673788 753244 673794 753256
rect 676030 753244 676036 753256
rect 676088 753244 676094 753296
rect 42150 753040 42156 753092
rect 42208 753080 42214 753092
rect 43162 753080 43168 753092
rect 42208 753052 43168 753080
rect 42208 753040 42214 753052
rect 43162 753040 43168 753052
rect 43220 753040 43226 753092
rect 42150 751748 42156 751800
rect 42208 751788 42214 751800
rect 42886 751788 42892 751800
rect 42208 751760 42892 751788
rect 42208 751748 42214 751760
rect 42886 751748 42892 751760
rect 42944 751748 42950 751800
rect 42150 751068 42156 751120
rect 42208 751108 42214 751120
rect 43530 751108 43536 751120
rect 42208 751080 43536 751108
rect 42208 751068 42214 751080
rect 43530 751068 43536 751080
rect 43588 751068 43594 751120
rect 42058 750592 42064 750644
rect 42116 750632 42122 750644
rect 43438 750632 43444 750644
rect 42116 750604 43444 750632
rect 42116 750592 42122 750604
rect 43438 750592 43444 750604
rect 43496 750592 43502 750644
rect 43438 750456 43444 750508
rect 43496 750496 43502 750508
rect 44082 750496 44088 750508
rect 43496 750468 44088 750496
rect 43496 750456 43502 750468
rect 44082 750456 44088 750468
rect 44140 750456 44146 750508
rect 672166 749912 672172 749964
rect 672224 749952 672230 749964
rect 679250 749952 679256 749964
rect 672224 749924 679256 749952
rect 672224 749912 672230 749924
rect 679250 749912 679256 749924
rect 679308 749912 679314 749964
rect 42150 749776 42156 749828
rect 42208 749816 42214 749828
rect 43806 749816 43812 749828
rect 42208 749788 43812 749816
rect 42208 749776 42214 749788
rect 43806 749776 43812 749788
rect 43864 749776 43870 749828
rect 43162 749096 43168 749148
rect 43220 749136 43226 749148
rect 43714 749136 43720 749148
rect 43220 749108 43720 749136
rect 43220 749096 43226 749108
rect 43714 749096 43720 749108
rect 43772 749096 43778 749148
rect 42610 748960 42616 749012
rect 42668 749000 42674 749012
rect 43714 749000 43720 749012
rect 42668 748972 43720 749000
rect 42668 748960 42674 748972
rect 43714 748960 43720 748972
rect 43772 748960 43778 749012
rect 654686 748960 654692 749012
rect 654744 749000 654750 749012
rect 668854 749000 668860 749012
rect 654744 748972 668860 749000
rect 654744 748960 654750 748972
rect 668854 748960 668860 748972
rect 668912 748960 668918 749012
rect 42150 746920 42156 746972
rect 42208 746960 42214 746972
rect 43070 746960 43076 746972
rect 42208 746932 43076 746960
rect 42208 746920 42214 746932
rect 43070 746920 43076 746932
rect 43128 746920 43134 746972
rect 42150 746716 42156 746768
rect 42208 746756 42214 746768
rect 43714 746756 43720 746768
rect 42208 746728 43720 746756
rect 42208 746716 42214 746728
rect 43714 746716 43720 746728
rect 43772 746716 43778 746768
rect 42150 746240 42156 746292
rect 42208 746280 42214 746292
rect 43438 746280 43444 746292
rect 42208 746252 43444 746280
rect 42208 746240 42214 746252
rect 43438 746240 43444 746252
rect 43496 746240 43502 746292
rect 42150 745424 42156 745476
rect 42208 745464 42214 745476
rect 43898 745464 43904 745476
rect 42208 745436 43904 745464
rect 42208 745424 42214 745436
rect 43898 745424 43904 745436
rect 43956 745424 43962 745476
rect 42150 743724 42156 743776
rect 42208 743764 42214 743776
rect 44082 743764 44088 743776
rect 42208 743736 44088 743764
rect 42208 743724 42214 743736
rect 44082 743724 44088 743736
rect 44140 743724 44146 743776
rect 42150 743248 42156 743300
rect 42208 743288 42214 743300
rect 43622 743288 43628 743300
rect 42208 743260 43628 743288
rect 42208 743248 42214 743260
rect 43622 743248 43628 743260
rect 43680 743248 43686 743300
rect 42150 742568 42156 742620
rect 42208 742608 42214 742620
rect 43162 742608 43168 742620
rect 42208 742580 43168 742608
rect 42208 742568 42214 742580
rect 43162 742568 43168 742580
rect 43220 742568 43226 742620
rect 48682 739712 48688 739764
rect 48740 739752 48746 739764
rect 58434 739752 58440 739764
rect 48740 739724 58440 739752
rect 48740 739712 48746 739724
rect 58434 739712 58440 739724
rect 58492 739712 58498 739764
rect 673914 738420 673920 738472
rect 673972 738460 673978 738472
rect 674650 738460 674656 738472
rect 673972 738432 674656 738460
rect 673972 738420 673978 738432
rect 674650 738420 674656 738432
rect 674708 738420 674714 738472
rect 655514 738284 655520 738336
rect 655572 738324 655578 738336
rect 674650 738324 674656 738336
rect 655572 738296 674656 738324
rect 655572 738284 655578 738296
rect 674650 738284 674656 738296
rect 674708 738284 674714 738336
rect 654134 736244 654140 736296
rect 654192 736284 654198 736296
rect 661126 736284 661132 736296
rect 654192 736256 661132 736284
rect 654192 736244 654198 736256
rect 661126 736244 661132 736256
rect 661184 736244 661190 736296
rect 674006 735428 674012 735480
rect 674064 735468 674070 735480
rect 675386 735468 675392 735480
rect 674064 735440 675392 735468
rect 674064 735428 674070 735440
rect 675386 735428 675392 735440
rect 675444 735428 675450 735480
rect 673730 734748 673736 734800
rect 673788 734788 673794 734800
rect 675386 734788 675392 734800
rect 673788 734760 675392 734788
rect 673788 734748 673794 734760
rect 675386 734748 675392 734760
rect 675444 734748 675450 734800
rect 673638 734340 673644 734392
rect 673696 734380 673702 734392
rect 675386 734380 675392 734392
rect 673696 734352 675392 734380
rect 673696 734340 673702 734352
rect 675386 734340 675392 734352
rect 675444 734340 675450 734392
rect 673546 733592 673552 733644
rect 673604 733632 673610 733644
rect 675386 733632 675392 733644
rect 673604 733604 675392 733632
rect 673604 733592 673610 733604
rect 675386 733592 675392 733604
rect 675444 733592 675450 733644
rect 673822 732300 673828 732352
rect 673880 732340 673886 732352
rect 675386 732340 675392 732352
rect 673880 732312 675392 732340
rect 673880 732300 673886 732312
rect 675386 732300 675392 732312
rect 675444 732300 675450 732352
rect 674650 732028 674656 732080
rect 674708 732068 674714 732080
rect 675386 732068 675392 732080
rect 674708 732040 675392 732068
rect 674708 732028 674714 732040
rect 675386 732028 675392 732040
rect 675444 732028 675450 732080
rect 674006 731892 674012 731944
rect 674064 731932 674070 731944
rect 674650 731932 674656 731944
rect 674064 731904 674656 731932
rect 674064 731892 674070 731904
rect 674650 731892 674656 731904
rect 674708 731892 674714 731944
rect 41782 731348 41788 731400
rect 41840 731388 41846 731400
rect 51166 731388 51172 731400
rect 41840 731360 51172 731388
rect 41840 731348 41846 731360
rect 51166 731348 51172 731360
rect 51224 731348 51230 731400
rect 41506 731076 41512 731128
rect 41564 731116 41570 731128
rect 48866 731116 48872 731128
rect 41564 731088 48872 731116
rect 41564 731076 41570 731088
rect 48866 731076 48872 731088
rect 48924 731076 48930 731128
rect 41506 730668 41512 730720
rect 41564 730708 41570 730720
rect 51074 730708 51080 730720
rect 41564 730680 51080 730708
rect 41564 730668 41570 730680
rect 51074 730668 51080 730680
rect 51132 730668 51138 730720
rect 41506 730464 41512 730516
rect 41564 730504 41570 730516
rect 43254 730504 43260 730516
rect 41564 730476 43260 730504
rect 41564 730464 41570 730476
rect 43254 730464 43260 730476
rect 43312 730464 43318 730516
rect 673730 730464 673736 730516
rect 673788 730504 673794 730516
rect 675386 730504 675392 730516
rect 673788 730476 675392 730504
rect 673788 730464 673794 730476
rect 675386 730464 675392 730476
rect 675444 730464 675450 730516
rect 42518 729240 42524 729292
rect 42576 729280 42582 729292
rect 42978 729280 42984 729292
rect 42576 729252 42984 729280
rect 42576 729240 42582 729252
rect 42978 729240 42984 729252
rect 43036 729240 43042 729292
rect 674834 728900 674840 728952
rect 674892 728940 674898 728952
rect 675478 728940 675484 728952
rect 674892 728912 675484 728940
rect 674892 728900 674898 728912
rect 675478 728900 675484 728912
rect 675536 728900 675542 728952
rect 41782 728832 41788 728884
rect 41840 728872 41846 728884
rect 44266 728872 44272 728884
rect 41840 728844 44272 728872
rect 41840 728832 41846 728844
rect 44266 728832 44272 728844
rect 44324 728832 44330 728884
rect 42518 728696 42524 728748
rect 42576 728736 42582 728748
rect 63034 728736 63040 728748
rect 42576 728708 63040 728736
rect 42576 728696 42582 728708
rect 63034 728696 63040 728708
rect 63092 728696 63098 728748
rect 51166 725908 51172 725960
rect 51224 725948 51230 725960
rect 58434 725948 58440 725960
rect 51224 725920 58440 725948
rect 51224 725908 51230 725920
rect 58434 725908 58440 725920
rect 58492 725908 58498 725960
rect 673362 723120 673368 723172
rect 673420 723160 673426 723172
rect 678974 723160 678980 723172
rect 673420 723132 678980 723160
rect 673420 723120 673426 723132
rect 678974 723120 678980 723132
rect 679032 723120 679038 723172
rect 673914 722848 673920 722900
rect 673972 722888 673978 722900
rect 675478 722888 675484 722900
rect 673972 722860 675484 722888
rect 673972 722848 673978 722860
rect 675478 722848 675484 722860
rect 675536 722848 675542 722900
rect 674190 721284 674196 721336
rect 674248 721324 674254 721336
rect 674926 721324 674932 721336
rect 674248 721296 674932 721324
rect 674248 721284 674254 721296
rect 674926 721284 674932 721296
rect 674984 721284 674990 721336
rect 674006 721148 674012 721200
rect 674064 721188 674070 721200
rect 674190 721188 674196 721200
rect 674064 721160 674196 721188
rect 674064 721148 674070 721160
rect 674190 721148 674196 721160
rect 674248 721148 674254 721200
rect 703446 720400 703452 720452
rect 703504 720440 703510 720452
rect 709242 720440 709248 720452
rect 703504 720412 709248 720440
rect 703504 720400 703510 720412
rect 709242 720400 709248 720412
rect 709300 720400 709306 720452
rect 41506 719992 41512 720044
rect 41564 720032 41570 720044
rect 48590 720032 48596 720044
rect 41564 720004 48596 720032
rect 41564 719992 41570 720004
rect 48590 719992 48596 720004
rect 48648 719992 48654 720044
rect 704476 717624 708460 717652
rect 41322 717544 41328 717596
rect 41380 717584 41386 717596
rect 43806 717584 43812 717596
rect 41380 717556 43812 717584
rect 41380 717544 41386 717556
rect 43806 717544 43812 717556
rect 43864 717544 43870 717596
rect 704476 717528 704504 717624
rect 708432 717528 708460 717624
rect 704458 717476 704464 717528
rect 704516 717476 704522 717528
rect 708414 717476 708420 717528
rect 708472 717476 708478 717528
rect 708506 717448 708512 717460
rect 704476 717420 708512 717448
rect 704476 717392 704504 717420
rect 708506 717408 708512 717420
rect 708564 717408 708570 717460
rect 704458 717340 704464 717392
rect 704516 717340 704522 717392
rect 705378 717340 705384 717392
rect 705436 717380 705442 717392
rect 707494 717380 707500 717392
rect 705436 717352 707500 717380
rect 705436 717340 705442 717352
rect 707494 717340 707500 717352
rect 707552 717340 707558 717392
rect 707034 717312 707040 717324
rect 705764 717284 707040 717312
rect 705764 717256 705792 717284
rect 707034 717272 707040 717284
rect 707092 717272 707098 717324
rect 705746 717204 705752 717256
rect 705804 717204 705810 717256
rect 706206 717204 706212 717256
rect 706264 717244 706270 717256
rect 706574 717244 706580 717256
rect 706264 717216 706580 717244
rect 706264 717204 706270 717216
rect 706574 717204 706580 717216
rect 706632 717204 706638 717256
rect 705838 717136 705844 717188
rect 705896 717176 705902 717188
rect 707034 717176 707040 717188
rect 705896 717148 707040 717176
rect 705896 717136 705902 717148
rect 707034 717136 707040 717148
rect 707092 717136 707098 717188
rect 707586 717136 707592 717188
rect 707644 717136 707650 717188
rect 706298 717068 706304 717120
rect 706356 717108 706362 717120
rect 706574 717108 706580 717120
rect 706356 717080 706580 717108
rect 706356 717068 706362 717080
rect 706574 717068 706580 717080
rect 706632 717068 706638 717120
rect 705378 717000 705384 717052
rect 705436 717040 705442 717052
rect 707604 717040 707632 717136
rect 705436 717012 707632 717040
rect 705436 717000 705442 717012
rect 708046 717000 708052 717052
rect 708104 717000 708110 717052
rect 704918 716932 704924 716984
rect 704976 716972 704982 716984
rect 707954 716972 707960 716984
rect 704976 716944 707960 716972
rect 704976 716932 704982 716944
rect 707954 716932 707960 716944
rect 708012 716932 708018 716984
rect 704826 716864 704832 716916
rect 704884 716904 704890 716916
rect 708064 716904 708092 717000
rect 704884 716876 708092 716904
rect 704884 716864 704890 716876
rect 703538 716796 703544 716848
rect 703596 716836 703602 716848
rect 708874 716836 708880 716848
rect 703596 716808 708880 716836
rect 703596 716796 703602 716808
rect 708874 716796 708880 716808
rect 708932 716796 708938 716848
rect 42518 716592 42524 716644
rect 42576 716632 42582 716644
rect 53742 716632 53748 716644
rect 42576 716604 53748 716632
rect 42576 716592 42582 716604
rect 53742 716592 53748 716604
rect 53800 716592 53806 716644
rect 666462 716524 666468 716576
rect 666520 716564 666526 716576
rect 676030 716564 676036 716576
rect 666520 716536 676036 716564
rect 666520 716524 666526 716536
rect 676030 716524 676036 716536
rect 676088 716524 676094 716576
rect 663702 716116 663708 716168
rect 663760 716156 663766 716168
rect 676030 716156 676036 716168
rect 663760 716128 676036 716156
rect 663760 716116 663766 716128
rect 676030 716116 676036 716128
rect 676088 716116 676094 716168
rect 667106 715708 667112 715760
rect 667164 715748 667170 715760
rect 676030 715748 676036 715760
rect 667164 715720 676036 715748
rect 667164 715708 667170 715720
rect 676030 715708 676036 715720
rect 676088 715708 676094 715760
rect 670510 715232 670516 715284
rect 670568 715272 670574 715284
rect 676030 715272 676036 715284
rect 670568 715244 676036 715272
rect 670568 715232 670574 715244
rect 676030 715232 676036 715244
rect 676088 715232 676094 715284
rect 670234 714892 670240 714944
rect 670292 714932 670298 714944
rect 676030 714932 676036 714944
rect 670292 714904 676036 714932
rect 670292 714892 670298 714904
rect 676030 714892 676036 714904
rect 676088 714892 676094 714944
rect 50982 714824 50988 714876
rect 51040 714864 51046 714876
rect 58434 714864 58440 714876
rect 51040 714836 58440 714864
rect 51040 714824 51046 714836
rect 58434 714824 58440 714836
rect 58492 714824 58498 714876
rect 670142 714824 670148 714876
rect 670200 714864 670206 714876
rect 670510 714864 670516 714876
rect 670200 714836 670516 714864
rect 670200 714824 670206 714836
rect 670510 714824 670516 714836
rect 670568 714824 670574 714876
rect 673822 714076 673828 714128
rect 673880 714116 673886 714128
rect 675662 714116 675668 714128
rect 673880 714088 675668 714116
rect 673880 714076 673886 714088
rect 675662 714076 675668 714088
rect 675720 714076 675726 714128
rect 673086 714008 673092 714060
rect 673144 714048 673150 714060
rect 676030 714048 676036 714060
rect 673144 714020 676036 714048
rect 673144 714008 673150 714020
rect 676030 714008 676036 714020
rect 676088 714008 676094 714060
rect 41874 713804 41880 713856
rect 41932 713804 41938 713856
rect 41892 713584 41920 713804
rect 670326 713600 670332 713652
rect 670384 713640 670390 713652
rect 670602 713640 670608 713652
rect 670384 713612 670608 713640
rect 670384 713600 670390 713612
rect 670602 713600 670608 713612
rect 670660 713640 670666 713652
rect 676030 713640 676036 713652
rect 670660 713612 676036 713640
rect 670660 713600 670666 713612
rect 676030 713600 676036 713612
rect 676088 713600 676094 713652
rect 41874 713532 41880 713584
rect 41932 713532 41938 713584
rect 669038 713192 669044 713244
rect 669096 713232 669102 713244
rect 670602 713232 670608 713244
rect 669096 713204 670608 713232
rect 669096 713192 669102 713204
rect 670602 713192 670608 713204
rect 670660 713232 670666 713244
rect 676030 713232 676036 713244
rect 670660 713204 676036 713232
rect 670660 713192 670666 713204
rect 676030 713192 676036 713204
rect 676088 713192 676094 713244
rect 668578 712852 668584 712904
rect 668636 712892 668642 712904
rect 676030 712892 676036 712904
rect 668636 712864 676036 712892
rect 668636 712852 668642 712864
rect 676030 712852 676036 712864
rect 676088 712852 676094 712904
rect 669130 712444 669136 712496
rect 669188 712484 669194 712496
rect 670510 712484 670516 712496
rect 669188 712456 670516 712484
rect 669188 712444 669194 712456
rect 670510 712444 670516 712456
rect 670568 712484 670574 712496
rect 676030 712484 676036 712496
rect 670568 712456 676036 712484
rect 670568 712444 670574 712456
rect 676030 712444 676036 712456
rect 676088 712444 676094 712496
rect 674926 712036 674932 712088
rect 674984 712076 674990 712088
rect 676030 712076 676036 712088
rect 674984 712048 676036 712076
rect 674984 712036 674990 712048
rect 676030 712036 676036 712048
rect 676088 712036 676094 712088
rect 674558 711968 674564 712020
rect 674616 712008 674622 712020
rect 675938 712008 675944 712020
rect 674616 711980 675944 712008
rect 674616 711968 674622 711980
rect 675938 711968 675944 711980
rect 675996 711968 676002 712020
rect 674190 711900 674196 711952
rect 674248 711940 674254 711952
rect 675846 711940 675852 711952
rect 674248 711912 675852 711940
rect 674248 711900 674254 711912
rect 675846 711900 675852 711912
rect 675904 711900 675910 711952
rect 42150 711628 42156 711680
rect 42208 711668 42214 711680
rect 43070 711668 43076 711680
rect 42208 711640 43076 711668
rect 42208 711628 42214 711640
rect 43070 711628 43076 711640
rect 43128 711628 43134 711680
rect 43070 711492 43076 711544
rect 43128 711532 43134 711544
rect 43346 711532 43352 711544
rect 43128 711504 43352 711532
rect 43128 711492 43134 711504
rect 43346 711492 43352 711504
rect 43404 711492 43410 711544
rect 42150 711084 42156 711136
rect 42208 711124 42214 711136
rect 42518 711124 42524 711136
rect 42208 711096 42524 711124
rect 42208 711084 42214 711096
rect 42518 711084 42524 711096
rect 42576 711084 42582 711136
rect 673546 710676 673552 710728
rect 673604 710716 673610 710728
rect 674006 710716 674012 710728
rect 673604 710688 674012 710716
rect 673604 710676 673610 710688
rect 674006 710676 674012 710688
rect 674064 710676 674070 710728
rect 674650 710676 674656 710728
rect 674708 710716 674714 710728
rect 675570 710716 675576 710728
rect 674708 710688 675576 710716
rect 674708 710676 674714 710688
rect 675570 710676 675576 710688
rect 675628 710676 675634 710728
rect 673730 710608 673736 710660
rect 673788 710648 673794 710660
rect 674834 710648 674840 710660
rect 673788 710620 674840 710648
rect 673788 710608 673794 710620
rect 674834 710608 674840 710620
rect 674892 710608 674898 710660
rect 674742 710540 674748 710592
rect 674800 710580 674806 710592
rect 676030 710580 676036 710592
rect 674800 710552 676036 710580
rect 674800 710540 674806 710552
rect 676030 710540 676036 710552
rect 676088 710540 676094 710592
rect 42150 709860 42156 709912
rect 42208 709900 42214 709912
rect 42794 709900 42800 709912
rect 42208 709872 42800 709900
rect 42208 709860 42214 709872
rect 42794 709860 42800 709872
rect 42852 709860 42858 709912
rect 42794 709724 42800 709776
rect 42852 709764 42858 709776
rect 43162 709764 43168 709776
rect 42852 709736 43168 709764
rect 42852 709724 42858 709736
rect 43162 709724 43168 709736
rect 43220 709724 43226 709776
rect 655974 709724 655980 709776
rect 656032 709764 656038 709776
rect 660942 709764 660948 709776
rect 656032 709736 660948 709764
rect 656032 709724 656038 709736
rect 660942 709724 660948 709736
rect 661000 709724 661006 709776
rect 43162 709588 43168 709640
rect 43220 709628 43226 709640
rect 43714 709628 43720 709640
rect 43220 709600 43720 709628
rect 43220 709588 43226 709600
rect 43714 709588 43720 709600
rect 43772 709588 43778 709640
rect 674466 709248 674472 709300
rect 674524 709288 674530 709300
rect 676030 709288 676036 709300
rect 674524 709260 676036 709288
rect 674524 709248 674530 709260
rect 676030 709248 676036 709260
rect 676088 709248 676094 709300
rect 42150 708432 42156 708484
rect 42208 708472 42214 708484
rect 43254 708472 43260 708484
rect 42208 708444 43260 708472
rect 42208 708432 42214 708444
rect 43254 708432 43260 708444
rect 43312 708432 43318 708484
rect 674374 708228 674380 708280
rect 674432 708268 674438 708280
rect 676030 708268 676036 708280
rect 674432 708240 676036 708268
rect 674432 708228 674438 708240
rect 676030 708228 676036 708240
rect 676088 708228 676094 708280
rect 42150 708024 42156 708076
rect 42208 708064 42214 708076
rect 43438 708064 43444 708076
rect 42208 708036 43444 708064
rect 42208 708024 42214 708036
rect 43438 708024 43444 708036
rect 43496 708024 43502 708076
rect 674282 707820 674288 707872
rect 674340 707860 674346 707872
rect 676030 707860 676036 707872
rect 674340 707832 676036 707860
rect 674340 707820 674346 707832
rect 676030 707820 676036 707832
rect 676088 707820 676094 707872
rect 676030 707412 676036 707464
rect 676088 707452 676094 707464
rect 676582 707452 676588 707464
rect 676088 707424 676588 707452
rect 676088 707412 676094 707424
rect 676582 707412 676588 707424
rect 676640 707412 676646 707464
rect 42150 707208 42156 707260
rect 42208 707248 42214 707260
rect 44082 707248 44088 707260
rect 42208 707220 44088 707248
rect 42208 707208 42214 707220
rect 44082 707208 44088 707220
rect 44140 707208 44146 707260
rect 42150 706732 42156 706784
rect 42208 706772 42214 706784
rect 43070 706772 43076 706784
rect 42208 706744 43076 706772
rect 42208 706732 42214 706744
rect 43070 706732 43076 706744
rect 43128 706732 43134 706784
rect 671798 705440 671804 705492
rect 671856 705480 671862 705492
rect 675938 705480 675944 705492
rect 671856 705452 675944 705480
rect 671856 705440 671862 705452
rect 675938 705440 675944 705452
rect 675996 705440 676002 705492
rect 42242 704828 42248 704880
rect 42300 704868 42306 704880
rect 42978 704868 42984 704880
rect 42300 704840 42984 704868
rect 42300 704828 42306 704840
rect 42978 704828 42984 704840
rect 43036 704828 43042 704880
rect 42058 704216 42064 704268
rect 42116 704256 42122 704268
rect 43898 704256 43904 704268
rect 42116 704228 43904 704256
rect 42116 704216 42122 704228
rect 43898 704216 43904 704228
rect 43956 704216 43962 704268
rect 42058 702856 42064 702908
rect 42116 702896 42122 702908
rect 43806 702896 43812 702908
rect 42116 702868 43812 702896
rect 42116 702856 42122 702868
rect 43806 702856 43812 702868
rect 43864 702856 43870 702908
rect 42058 702380 42064 702432
rect 42116 702420 42122 702432
rect 43530 702420 43536 702432
rect 42116 702392 43536 702420
rect 42116 702380 42122 702392
rect 43530 702380 43536 702392
rect 43588 702380 43594 702432
rect 53742 701020 53748 701072
rect 53800 701060 53806 701072
rect 58158 701060 58164 701072
rect 53800 701032 58164 701060
rect 53800 701020 53806 701032
rect 58158 701020 58164 701032
rect 58216 701020 58222 701072
rect 42150 700408 42156 700460
rect 42208 700448 42214 700460
rect 43622 700448 43628 700460
rect 42208 700420 43628 700448
rect 42208 700408 42214 700420
rect 43622 700408 43628 700420
rect 43680 700408 43686 700460
rect 42150 700000 42156 700052
rect 42208 700040 42214 700052
rect 42886 700040 42892 700052
rect 42208 700012 42892 700040
rect 42208 700000 42214 700012
rect 42886 700000 42892 700012
rect 42944 700000 42950 700052
rect 670510 699728 670516 699780
rect 670568 699728 670574 699780
rect 670528 699564 670556 699728
rect 674742 699660 674748 699712
rect 674800 699700 674806 699712
rect 675478 699700 675484 699712
rect 674800 699672 675484 699700
rect 674800 699660 674806 699672
rect 675478 699660 675484 699672
rect 675536 699660 675542 699712
rect 674650 699592 674656 699644
rect 674708 699632 674714 699644
rect 675570 699632 675576 699644
rect 674708 699604 675576 699632
rect 674708 699592 674714 699604
rect 675570 699592 675576 699604
rect 675628 699592 675634 699644
rect 670602 699564 670608 699576
rect 670528 699536 670608 699564
rect 670602 699524 670608 699536
rect 670660 699524 670666 699576
rect 42058 699388 42064 699440
rect 42116 699428 42122 699440
rect 42794 699428 42800 699440
rect 42116 699400 42800 699428
rect 42116 699388 42122 699400
rect 42794 699388 42800 699400
rect 42852 699388 42858 699440
rect 654870 696396 654876 696448
rect 654928 696436 654934 696448
rect 663794 696436 663800 696448
rect 654928 696408 663800 696436
rect 654928 696396 654934 696408
rect 663794 696396 663800 696408
rect 663852 696396 663858 696448
rect 655514 691364 655520 691416
rect 655572 691404 655578 691416
rect 674558 691404 674564 691416
rect 655572 691376 674564 691404
rect 655572 691364 655578 691376
rect 674558 691364 674564 691376
rect 674616 691364 674622 691416
rect 673638 690412 673644 690464
rect 673696 690452 673702 690464
rect 675386 690452 675392 690464
rect 673696 690424 675392 690452
rect 673696 690412 673702 690424
rect 675386 690412 675392 690424
rect 675444 690412 675450 690464
rect 673178 689120 673184 689172
rect 673236 689160 673242 689172
rect 675478 689160 675484 689172
rect 673236 689132 675484 689160
rect 673236 689120 673242 689132
rect 675478 689120 675484 689132
rect 675536 689120 675542 689172
rect 672994 688576 673000 688628
rect 673052 688616 673058 688628
rect 675386 688616 675392 688628
rect 673052 688588 675392 688616
rect 673052 688576 673058 688588
rect 675386 688576 675392 688588
rect 675444 688576 675450 688628
rect 41506 688372 41512 688424
rect 41564 688412 41570 688424
rect 48682 688412 48688 688424
rect 41564 688384 48688 688412
rect 41564 688372 41570 688384
rect 48682 688372 48688 688384
rect 48740 688372 48746 688424
rect 41690 687828 41696 687880
rect 41748 687868 41754 687880
rect 53834 687868 53840 687880
rect 41748 687840 53840 687868
rect 41748 687828 41754 687840
rect 53834 687828 53840 687840
rect 53892 687828 53898 687880
rect 41782 687692 41788 687744
rect 41840 687732 41846 687744
rect 51166 687732 51172 687744
rect 41840 687704 51172 687732
rect 41840 687692 41846 687704
rect 51166 687692 51172 687704
rect 51224 687692 51230 687744
rect 673270 687284 673276 687336
rect 673328 687324 673334 687336
rect 675386 687324 675392 687336
rect 673328 687296 675392 687324
rect 673328 687284 673334 687296
rect 675386 687284 675392 687296
rect 675444 687284 675450 687336
rect 51074 687216 51080 687268
rect 51132 687256 51138 687268
rect 58434 687256 58440 687268
rect 51132 687228 58440 687256
rect 51132 687216 51138 687228
rect 58434 687216 58440 687228
rect 58492 687216 58498 687268
rect 674558 687012 674564 687064
rect 674616 687052 674622 687064
rect 675478 687052 675484 687064
rect 674616 687024 675484 687052
rect 674616 687012 674622 687024
rect 675478 687012 675484 687024
rect 675536 687012 675542 687064
rect 674282 685448 674288 685500
rect 674340 685488 674346 685500
rect 675386 685488 675392 685500
rect 674340 685460 675392 685488
rect 674340 685448 674346 685460
rect 675386 685448 675392 685460
rect 675444 685448 675450 685500
rect 42794 684428 42800 684480
rect 42852 684468 42858 684480
rect 62758 684468 62764 684480
rect 42852 684440 62764 684468
rect 42852 684428 42858 684440
rect 62758 684428 62764 684440
rect 62816 684428 62822 684480
rect 673822 683612 673828 683664
rect 673880 683652 673886 683664
rect 675478 683652 675484 683664
rect 673880 683624 675484 683652
rect 673880 683612 673886 683624
rect 675478 683612 675484 683624
rect 675536 683612 675542 683664
rect 654134 683408 654140 683460
rect 654192 683448 654198 683460
rect 669130 683448 669136 683460
rect 654192 683420 669136 683448
rect 654192 683408 654198 683420
rect 669130 683408 669136 683420
rect 669188 683408 669194 683460
rect 673086 678988 673092 679040
rect 673144 679028 673150 679040
rect 678974 679028 678980 679040
rect 673144 679000 678980 679028
rect 673144 678988 673150 679000
rect 678974 678988 678980 679000
rect 679032 678988 679038 679040
rect 41782 678172 41788 678224
rect 41840 678212 41846 678224
rect 43254 678212 43260 678224
rect 41840 678184 43260 678212
rect 41840 678172 41846 678184
rect 43254 678172 43260 678184
rect 43312 678172 43318 678224
rect 41782 677016 41788 677068
rect 41840 677056 41846 677068
rect 48682 677056 48688 677068
rect 41840 677028 48688 677056
rect 41840 677016 41846 677028
rect 48682 677016 48688 677028
rect 48740 677016 48746 677068
rect 48866 673480 48872 673532
rect 48924 673520 48930 673532
rect 58434 673520 58440 673532
rect 48924 673492 58440 673520
rect 48924 673480 48930 673492
rect 58434 673480 58440 673492
rect 58492 673480 58498 673532
rect 41322 673412 41328 673464
rect 41380 673452 41386 673464
rect 43070 673452 43076 673464
rect 41380 673424 43076 673452
rect 41380 673412 41386 673424
rect 43070 673412 43076 673424
rect 43128 673412 43134 673464
rect 703446 672324 703452 672376
rect 703504 672364 703510 672376
rect 703504 672336 709012 672364
rect 703504 672324 703510 672336
rect 708984 672308 709012 672336
rect 703538 672256 703544 672308
rect 703596 672296 703602 672308
rect 708874 672296 708880 672308
rect 703596 672268 708880 672296
rect 703596 672256 703602 672268
rect 708874 672256 708880 672268
rect 708932 672256 708938 672308
rect 708966 672256 708972 672308
rect 709024 672256 709030 672308
rect 708046 672228 708052 672240
rect 704844 672200 708052 672228
rect 704844 672104 704872 672200
rect 708046 672188 708052 672200
rect 708104 672188 708110 672240
rect 704918 672120 704924 672172
rect 704976 672160 704982 672172
rect 707954 672160 707960 672172
rect 704976 672132 707960 672160
rect 704976 672120 704982 672132
rect 707954 672120 707960 672132
rect 708012 672120 708018 672172
rect 704826 672052 704832 672104
rect 704884 672052 704890 672104
rect 707034 672092 707040 672104
rect 705764 672064 707040 672092
rect 705764 671968 705792 672064
rect 707034 672052 707040 672064
rect 707092 672052 707098 672104
rect 706666 672024 706672 672036
rect 706224 671996 706672 672024
rect 706224 671968 706252 671996
rect 706666 671984 706672 671996
rect 706724 671984 706730 672036
rect 705746 671916 705752 671968
rect 705804 671916 705810 671968
rect 706206 671916 706212 671968
rect 706264 671916 706270 671968
rect 706298 671916 706304 671968
rect 706356 671956 706362 671968
rect 706574 671956 706580 671968
rect 706356 671928 706580 671956
rect 706356 671916 706362 671928
rect 706574 671916 706580 671928
rect 706632 671916 706638 671968
rect 705838 671848 705844 671900
rect 705896 671888 705902 671900
rect 707034 671888 707040 671900
rect 705896 671860 707040 671888
rect 705896 671848 705902 671860
rect 707034 671848 707040 671860
rect 707092 671848 707098 671900
rect 707586 671848 707592 671900
rect 707644 671848 707650 671900
rect 705378 671780 705384 671832
rect 705436 671820 705442 671832
rect 707494 671820 707500 671832
rect 705436 671792 707500 671820
rect 705436 671780 705442 671792
rect 707494 671780 707500 671792
rect 707552 671780 707558 671832
rect 705286 671712 705292 671764
rect 705344 671752 705350 671764
rect 707604 671752 707632 671848
rect 705344 671724 707632 671752
rect 705344 671712 705350 671724
rect 708506 671712 708512 671764
rect 708564 671712 708570 671764
rect 704458 671644 704464 671696
rect 704516 671684 704522 671696
rect 708414 671684 708420 671696
rect 704516 671656 708420 671684
rect 704516 671644 704522 671656
rect 708414 671644 708420 671656
rect 708472 671644 708478 671696
rect 704366 671576 704372 671628
rect 704424 671616 704430 671628
rect 708524 671616 708552 671712
rect 704424 671588 708552 671616
rect 704424 671576 704430 671588
rect 674742 671236 674748 671288
rect 674800 671276 674806 671288
rect 675202 671276 675208 671288
rect 674800 671248 675208 671276
rect 674800 671236 674806 671248
rect 675202 671236 675208 671248
rect 675260 671236 675266 671288
rect 668946 670964 668952 671016
rect 669004 671004 669010 671016
rect 676030 671004 676036 671016
rect 669004 670976 676036 671004
rect 669004 670964 669010 670976
rect 676030 670964 676036 670976
rect 676088 670964 676094 671016
rect 661034 670760 661040 670812
rect 661092 670800 661098 670812
rect 676214 670800 676220 670812
rect 661092 670772 676220 670800
rect 661092 670760 661098 670772
rect 676214 670760 676220 670772
rect 676272 670760 676278 670812
rect 44174 670692 44180 670744
rect 44232 670732 44238 670744
rect 48774 670732 48780 670744
rect 44232 670704 48780 670732
rect 44232 670692 44238 670704
rect 48774 670692 48780 670704
rect 48832 670692 48838 670744
rect 44082 670624 44088 670676
rect 44140 670624 44146 670676
rect 41874 670556 41880 670608
rect 41932 670556 41938 670608
rect 41966 670556 41972 670608
rect 42024 670596 42030 670608
rect 42702 670596 42708 670608
rect 42024 670568 42708 670596
rect 42024 670556 42030 670568
rect 42702 670556 42708 670568
rect 42760 670556 42766 670608
rect 41892 670404 41920 670556
rect 41874 670352 41880 670404
rect 41932 670352 41938 670404
rect 44100 670256 44128 670624
rect 663886 670556 663892 670608
rect 663944 670596 663950 670608
rect 676030 670596 676036 670608
rect 663944 670568 676036 670596
rect 663944 670556 663950 670568
rect 676030 670556 676036 670568
rect 676088 670556 676094 670608
rect 670234 670284 670240 670336
rect 670292 670324 670298 670336
rect 676214 670324 676220 670336
rect 670292 670296 676220 670324
rect 670292 670284 670298 670296
rect 676214 670284 676220 670296
rect 676272 670284 676278 670336
rect 44100 670228 44220 670256
rect 44192 670200 44220 670228
rect 44174 670148 44180 670200
rect 44232 670148 44238 670200
rect 674558 668992 674564 669044
rect 674616 669032 674622 669044
rect 676030 669032 676036 669044
rect 674616 669004 676036 669032
rect 674616 668992 674622 669004
rect 676030 668992 676036 669004
rect 676088 668992 676094 669044
rect 670510 668652 670516 668704
rect 670568 668692 670574 668704
rect 676214 668692 676220 668704
rect 670568 668664 676220 668692
rect 670568 668652 670574 668664
rect 676214 668652 676220 668664
rect 676272 668652 676278 668704
rect 42058 668448 42064 668500
rect 42116 668488 42122 668500
rect 43990 668488 43996 668500
rect 42116 668460 43996 668488
rect 42116 668448 42122 668460
rect 43990 668448 43996 668460
rect 44048 668448 44054 668500
rect 673086 668040 673092 668092
rect 673144 668080 673150 668092
rect 675938 668080 675944 668092
rect 673144 668052 675944 668080
rect 673144 668040 673150 668052
rect 675938 668040 675944 668052
rect 675996 668040 676002 668092
rect 674742 667904 674748 667956
rect 674800 667944 674806 667956
rect 676030 667944 676036 667956
rect 674800 667916 676036 667944
rect 674800 667904 674806 667916
rect 676030 667904 676036 667916
rect 676088 667904 676094 667956
rect 673914 667836 673920 667888
rect 673972 667876 673978 667888
rect 676122 667876 676128 667888
rect 673972 667848 676128 667876
rect 673972 667836 673978 667848
rect 676122 667836 676128 667848
rect 676180 667836 676186 667888
rect 674650 667768 674656 667820
rect 674708 667808 674714 667820
rect 676030 667808 676036 667820
rect 674708 667780 676036 667808
rect 674708 667768 674714 667780
rect 676030 667768 676036 667780
rect 676088 667768 676094 667820
rect 42150 667700 42156 667752
rect 42208 667740 42214 667752
rect 44082 667740 44088 667752
rect 42208 667712 44088 667740
rect 42208 667700 42214 667712
rect 44082 667700 44088 667712
rect 44140 667700 44146 667752
rect 670602 667700 670608 667752
rect 670660 667740 670666 667752
rect 675938 667740 675944 667752
rect 670660 667712 675944 667740
rect 670660 667700 670666 667712
rect 675938 667700 675944 667712
rect 675996 667700 676002 667752
rect 42150 666680 42156 666732
rect 42208 666720 42214 666732
rect 43898 666720 43904 666732
rect 42208 666692 43904 666720
rect 42208 666680 42214 666692
rect 43898 666680 43904 666692
rect 43956 666680 43962 666732
rect 42150 665388 42156 665440
rect 42208 665428 42214 665440
rect 42702 665428 42708 665440
rect 42208 665400 42708 665428
rect 42208 665388 42214 665400
rect 42702 665388 42708 665400
rect 42760 665388 42766 665440
rect 675202 665116 675208 665168
rect 675260 665156 675266 665168
rect 676030 665156 676036 665168
rect 675260 665128 676036 665156
rect 675260 665116 675266 665128
rect 676030 665116 676036 665128
rect 676088 665116 676094 665168
rect 673730 665048 673736 665100
rect 673788 665088 673794 665100
rect 676122 665088 676128 665100
rect 673788 665060 676128 665088
rect 673788 665048 673794 665060
rect 676122 665048 676128 665060
rect 676180 665048 676186 665100
rect 42150 664640 42156 664692
rect 42208 664680 42214 664692
rect 43530 664680 43536 664692
rect 42208 664652 43536 664680
rect 42208 664640 42214 664652
rect 43530 664640 43536 664652
rect 43588 664640 43594 664692
rect 42150 664164 42156 664216
rect 42208 664204 42214 664216
rect 43254 664204 43260 664216
rect 42208 664176 43260 664204
rect 42208 664164 42214 664176
rect 43254 664164 43260 664176
rect 43312 664164 43318 664216
rect 42150 663552 42156 663604
rect 42208 663592 42214 663604
rect 43070 663592 43076 663604
rect 42208 663564 43076 663592
rect 42208 663552 42214 663564
rect 43070 663552 43076 663564
rect 43128 663552 43134 663604
rect 48958 662396 48964 662448
rect 49016 662436 49022 662448
rect 58434 662436 58440 662448
rect 49016 662408 58440 662436
rect 49016 662396 49022 662408
rect 58434 662396 58440 662408
rect 58492 662396 58498 662448
rect 42150 661036 42156 661088
rect 42208 661076 42214 661088
rect 44082 661076 44088 661088
rect 42208 661048 44088 661076
rect 42208 661036 42214 661048
rect 44082 661036 44088 661048
rect 44140 661036 44146 661088
rect 42150 660492 42156 660544
rect 42208 660532 42214 660544
rect 43622 660532 43628 660544
rect 42208 660504 43628 660532
rect 42208 660492 42214 660504
rect 43622 660492 43628 660504
rect 43680 660492 43686 660544
rect 42150 659880 42156 659932
rect 42208 659920 42214 659932
rect 43162 659920 43168 659932
rect 42208 659892 43168 659920
rect 42208 659880 42214 659892
rect 43162 659880 43168 659892
rect 43220 659880 43226 659932
rect 672350 659676 672356 659728
rect 672408 659716 672414 659728
rect 678974 659716 678980 659728
rect 672408 659688 678980 659716
rect 672408 659676 672414 659688
rect 678974 659676 678980 659688
rect 679032 659676 679038 659728
rect 42150 658996 42156 659048
rect 42208 659036 42214 659048
rect 43806 659036 43812 659048
rect 42208 659008 43812 659036
rect 42208 658996 42214 659008
rect 43806 658996 43812 659008
rect 43864 658996 43870 659048
rect 42150 657228 42156 657280
rect 42208 657268 42214 657280
rect 43346 657268 43352 657280
rect 42208 657240 43352 657268
rect 42208 657228 42214 657240
rect 43346 657228 43352 657240
rect 43404 657228 43410 657280
rect 656802 657024 656808 657076
rect 656860 657064 656866 657076
rect 663702 657064 663708 657076
rect 656860 657036 663708 657064
rect 656860 657024 656866 657036
rect 663702 657024 663708 657036
rect 663760 657024 663766 657076
rect 42150 656820 42156 656872
rect 42208 656860 42214 656872
rect 43714 656860 43720 656872
rect 42208 656832 43720 656860
rect 42208 656820 42214 656832
rect 43714 656820 43720 656832
rect 43772 656820 43778 656872
rect 42150 656140 42156 656192
rect 42208 656180 42214 656192
rect 42978 656180 42984 656192
rect 42208 656152 42984 656180
rect 42208 656140 42214 656152
rect 42978 656140 42984 656152
rect 43036 656140 43042 656192
rect 674374 649544 674380 649596
rect 674432 649584 674438 649596
rect 675386 649584 675392 649596
rect 674432 649556 675392 649584
rect 674432 649544 674438 649556
rect 675386 649544 675392 649556
rect 675444 649544 675450 649596
rect 53834 648592 53840 648644
rect 53892 648632 53898 648644
rect 59170 648632 59176 648644
rect 53892 648604 59176 648632
rect 53892 648592 53898 648604
rect 59170 648592 59176 648604
rect 59228 648592 59234 648644
rect 673546 647708 673552 647760
rect 673604 647748 673610 647760
rect 675478 647748 675484 647760
rect 673604 647720 675484 647748
rect 673604 647708 673610 647720
rect 675478 647708 675484 647720
rect 675536 647708 675542 647760
rect 674466 647300 674472 647352
rect 674524 647340 674530 647352
rect 674742 647340 674748 647352
rect 674524 647312 674748 647340
rect 674524 647300 674530 647312
rect 674742 647300 674748 647312
rect 674800 647300 674806 647352
rect 655514 647164 655520 647216
rect 655572 647204 655578 647216
rect 674742 647204 674748 647216
rect 655572 647176 674748 647204
rect 655572 647164 655578 647176
rect 674742 647164 674748 647176
rect 674800 647164 674806 647216
rect 673730 645396 673736 645448
rect 673788 645436 673794 645448
rect 675386 645436 675392 645448
rect 673788 645408 675392 645436
rect 673788 645396 673794 645408
rect 675386 645396 675392 645408
rect 675444 645396 675450 645448
rect 41506 645124 41512 645176
rect 41564 645164 41570 645176
rect 51074 645164 51080 645176
rect 41564 645136 51080 645164
rect 41564 645124 41570 645136
rect 51074 645124 51080 645136
rect 51132 645124 51138 645176
rect 41506 644716 41512 644768
rect 41564 644756 41570 644768
rect 48866 644756 48872 644768
rect 41564 644728 48872 644756
rect 41564 644716 41570 644728
rect 48866 644716 48872 644728
rect 48924 644716 48930 644768
rect 41506 644580 41512 644632
rect 41564 644620 41570 644632
rect 53742 644620 53748 644632
rect 41564 644592 53748 644620
rect 41564 644580 41570 644592
rect 53742 644580 53748 644592
rect 53800 644580 53806 644632
rect 674650 644580 674656 644632
rect 674708 644620 674714 644632
rect 675386 644620 675392 644632
rect 674708 644592 675392 644620
rect 674708 644580 674714 644592
rect 675386 644580 675392 644592
rect 675444 644580 675450 644632
rect 673914 644104 673920 644156
rect 673972 644144 673978 644156
rect 675386 644144 675392 644156
rect 673972 644116 675392 644144
rect 673972 644104 673978 644116
rect 675386 644104 675392 644116
rect 675444 644104 675450 644156
rect 41506 643424 41512 643476
rect 41564 643464 41570 643476
rect 44358 643464 44364 643476
rect 41564 643436 44364 643464
rect 41564 643424 41570 643436
rect 44358 643424 44364 643436
rect 44416 643424 44422 643476
rect 674190 643356 674196 643408
rect 674248 643396 674254 643408
rect 675386 643396 675392 643408
rect 674248 643368 675392 643396
rect 674248 643356 674254 643368
rect 675386 643356 675392 643368
rect 675444 643356 675450 643408
rect 42886 643152 42892 643204
rect 42944 643192 42950 643204
rect 62574 643192 62580 643204
rect 42944 643164 62580 643192
rect 42944 643152 42950 643164
rect 62574 643152 62580 643164
rect 62632 643152 62638 643204
rect 654870 643084 654876 643136
rect 654928 643124 654934 643136
rect 666462 643124 666468 643136
rect 654928 643096 666468 643124
rect 654928 643084 654934 643096
rect 666462 643084 666468 643096
rect 666520 643084 666526 643136
rect 674006 642064 674012 642116
rect 674064 642104 674070 642116
rect 675386 642104 675392 642116
rect 674064 642076 675392 642104
rect 674064 642064 674070 642076
rect 675386 642064 675392 642076
rect 675444 642064 675450 642116
rect 674742 641860 674748 641912
rect 674800 641900 674806 641912
rect 675386 641900 675392 641912
rect 674800 641872 675392 641900
rect 674800 641860 674806 641872
rect 675386 641860 675392 641872
rect 675444 641860 675450 641912
rect 674466 641656 674472 641708
rect 674524 641696 674530 641708
rect 674742 641696 674748 641708
rect 674524 641668 674748 641696
rect 674524 641656 674530 641668
rect 674742 641656 674748 641668
rect 674800 641656 674806 641708
rect 674466 640228 674472 640280
rect 674524 640268 674530 640280
rect 675386 640268 675392 640280
rect 674524 640240 675392 640268
rect 674524 640228 674530 640240
rect 675386 640228 675392 640240
rect 675444 640228 675450 640280
rect 674742 638664 674748 638716
rect 674800 638704 674806 638716
rect 675202 638704 675208 638716
rect 674800 638676 675208 638704
rect 674800 638664 674806 638676
rect 675202 638664 675208 638676
rect 675260 638664 675266 638716
rect 674650 638392 674656 638444
rect 674708 638432 674714 638444
rect 675478 638432 675484 638444
rect 674708 638404 675484 638432
rect 674708 638392 674714 638404
rect 675478 638392 675484 638404
rect 675536 638392 675542 638444
rect 674742 638188 674748 638240
rect 674800 638228 674806 638240
rect 675478 638228 675484 638240
rect 674800 638200 675484 638228
rect 674800 638188 674806 638200
rect 675478 638188 675484 638200
rect 675536 638188 675542 638240
rect 674282 638160 674288 638172
rect 674208 638132 674288 638160
rect 674208 637968 674236 638132
rect 674282 638120 674288 638132
rect 674340 638120 674346 638172
rect 674374 638120 674380 638172
rect 674432 638160 674438 638172
rect 675662 638160 675668 638172
rect 674432 638132 675668 638160
rect 674432 638120 674438 638132
rect 675662 638120 675668 638132
rect 675720 638120 675726 638172
rect 674190 637916 674196 637968
rect 674248 637916 674254 637968
rect 673086 637848 673092 637900
rect 673144 637888 673150 637900
rect 679158 637888 679164 637900
rect 673144 637860 679164 637888
rect 673144 637848 673150 637860
rect 679158 637848 679164 637860
rect 679216 637848 679222 637900
rect 675202 637508 675208 637560
rect 675260 637548 675266 637560
rect 679066 637548 679072 637560
rect 675260 637520 679072 637548
rect 675260 637508 675266 637520
rect 679066 637508 679072 637520
rect 679124 637508 679130 637560
rect 674006 637304 674012 637356
rect 674064 637344 674070 637356
rect 674190 637344 674196 637356
rect 674064 637316 674196 637344
rect 674064 637304 674070 637316
rect 674190 637304 674196 637316
rect 674248 637304 674254 637356
rect 673730 637168 673736 637220
rect 673788 637208 673794 637220
rect 674006 637208 674012 637220
rect 673788 637180 674012 637208
rect 673788 637168 673794 637180
rect 674006 637168 674012 637180
rect 674064 637168 674070 637220
rect 48866 634788 48872 634840
rect 48924 634828 48930 634840
rect 58434 634828 58440 634840
rect 48924 634800 58440 634828
rect 48924 634788 48930 634800
rect 58434 634788 58440 634800
rect 58492 634788 58498 634840
rect 41506 633632 41512 633684
rect 41564 633672 41570 633684
rect 48774 633672 48780 633684
rect 41564 633644 48780 633672
rect 41564 633632 41570 633644
rect 48774 633632 48780 633644
rect 48832 633632 48838 633684
rect 43898 629280 43904 629332
rect 43956 629320 43962 629332
rect 50982 629320 50988 629332
rect 43956 629292 50988 629320
rect 43956 629280 43962 629292
rect 50982 629280 50988 629292
rect 51040 629280 51046 629332
rect 654134 629280 654140 629332
rect 654192 629320 654198 629332
rect 667198 629320 667204 629332
rect 654192 629292 667204 629320
rect 654192 629280 654198 629292
rect 667198 629280 667204 629292
rect 667256 629280 667262 629332
rect 33042 627852 33048 627904
rect 33100 627892 33106 627904
rect 42518 627892 42524 627904
rect 33100 627864 42524 627892
rect 33100 627852 33106 627864
rect 42518 627852 42524 627864
rect 42576 627852 42582 627904
rect 41782 627376 41788 627428
rect 41840 627376 41846 627428
rect 41800 627088 41828 627376
rect 708506 627348 708512 627360
rect 704384 627320 708512 627348
rect 704384 627224 704412 627320
rect 708506 627308 708512 627320
rect 708564 627308 708570 627360
rect 704458 627240 704464 627292
rect 704516 627280 704522 627292
rect 708414 627280 708420 627292
rect 704516 627252 708420 627280
rect 704516 627240 704522 627252
rect 708414 627240 708420 627252
rect 708472 627240 708478 627292
rect 704366 627172 704372 627224
rect 704424 627172 704430 627224
rect 707494 627212 707500 627224
rect 705488 627184 707500 627212
rect 41782 627036 41788 627088
rect 41840 627036 41846 627088
rect 705286 627036 705292 627088
rect 705344 627076 705350 627088
rect 705488 627076 705516 627184
rect 707494 627172 707500 627184
rect 707552 627172 707558 627224
rect 707034 627144 707040 627156
rect 705764 627116 707040 627144
rect 705764 627088 705792 627116
rect 707034 627104 707040 627116
rect 707092 627104 707098 627156
rect 705344 627048 705516 627076
rect 705344 627036 705350 627048
rect 705746 627036 705752 627088
rect 705804 627036 705810 627088
rect 706206 627036 706212 627088
rect 706264 627076 706270 627088
rect 706574 627076 706580 627088
rect 706264 627048 706580 627076
rect 706264 627036 706270 627048
rect 706574 627036 706580 627048
rect 706632 627036 706638 627088
rect 705838 626968 705844 627020
rect 705896 627008 705902 627020
rect 707034 627008 707040 627020
rect 705896 626980 707040 627008
rect 705896 626968 705902 626980
rect 707034 626968 707040 626980
rect 707092 626968 707098 627020
rect 706298 626900 706304 626952
rect 706356 626940 706362 626952
rect 706574 626940 706580 626952
rect 706356 626912 706580 626940
rect 706356 626900 706362 626912
rect 706574 626900 706580 626912
rect 706632 626900 706638 626952
rect 705378 626832 705384 626884
rect 705436 626872 705442 626884
rect 707494 626872 707500 626884
rect 705436 626844 707500 626872
rect 705436 626832 705442 626844
rect 707494 626832 707500 626844
rect 707552 626832 707558 626884
rect 708046 626832 708052 626884
rect 708104 626832 708110 626884
rect 704918 626764 704924 626816
rect 704976 626804 704982 626816
rect 707954 626804 707960 626816
rect 704976 626776 707960 626804
rect 704976 626764 704982 626776
rect 707954 626764 707960 626776
rect 708012 626764 708018 626816
rect 704826 626696 704832 626748
rect 704884 626736 704890 626748
rect 708064 626736 708092 626832
rect 704884 626708 708092 626736
rect 704884 626696 704890 626708
rect 708966 626696 708972 626748
rect 709024 626696 709030 626748
rect 703538 626628 703544 626680
rect 703596 626668 703602 626680
rect 708874 626668 708880 626680
rect 703596 626640 708880 626668
rect 703596 626628 703602 626640
rect 708874 626628 708880 626640
rect 708932 626628 708938 626680
rect 703998 626560 704004 626612
rect 704056 626600 704062 626612
rect 708984 626600 709012 626696
rect 704056 626572 709012 626600
rect 704056 626560 704062 626572
rect 42150 625268 42156 625320
rect 42208 625308 42214 625320
rect 43530 625308 43536 625320
rect 42208 625280 43536 625308
rect 42208 625268 42214 625280
rect 43530 625268 43536 625280
rect 43588 625268 43594 625320
rect 42150 624656 42156 624708
rect 42208 624696 42214 624708
rect 43898 624696 43904 624708
rect 42208 624668 43904 624696
rect 42208 624656 42214 624668
rect 43898 624656 43904 624668
rect 43956 624656 43962 624708
rect 670602 624248 670608 624300
rect 670660 624288 670666 624300
rect 674558 624288 674564 624300
rect 670660 624260 674564 624288
rect 670660 624248 670666 624260
rect 674558 624248 674564 624260
rect 674616 624288 674622 624300
rect 676030 624288 676036 624300
rect 674616 624260 676036 624288
rect 674616 624248 674622 624260
rect 676030 624248 676036 624260
rect 676088 624248 676094 624300
rect 668854 624112 668860 624164
rect 668912 624152 668918 624164
rect 678974 624152 678980 624164
rect 668912 624124 678980 624152
rect 668912 624112 668918 624124
rect 678974 624112 678980 624124
rect 679032 624112 679038 624164
rect 667014 623976 667020 624028
rect 667072 624016 667078 624028
rect 676122 624016 676128 624028
rect 667072 623988 676128 624016
rect 667072 623976 667078 623988
rect 676122 623976 676128 623988
rect 676180 623976 676186 624028
rect 673362 623908 673368 623960
rect 673420 623948 673426 623960
rect 676030 623948 676036 623960
rect 673420 623920 676036 623948
rect 673420 623908 673426 623920
rect 676030 623908 676036 623920
rect 676088 623908 676094 623960
rect 661126 623840 661132 623892
rect 661184 623880 661190 623892
rect 676306 623880 676312 623892
rect 661184 623852 676312 623880
rect 661184 623840 661190 623852
rect 676306 623840 676312 623852
rect 676364 623840 676370 623892
rect 51074 623772 51080 623824
rect 51132 623812 51138 623824
rect 58434 623812 58440 623824
rect 51132 623784 58440 623812
rect 51132 623772 51138 623784
rect 58434 623772 58440 623784
rect 58492 623772 58498 623824
rect 670234 623772 670240 623824
rect 670292 623812 670298 623824
rect 670418 623812 670424 623824
rect 670292 623784 670424 623812
rect 670292 623772 670298 623784
rect 670418 623772 670424 623784
rect 670476 623812 670482 623824
rect 676214 623812 676220 623824
rect 670476 623784 676220 623812
rect 670476 623772 670482 623784
rect 676214 623772 676220 623784
rect 676272 623772 676278 623824
rect 674282 623704 674288 623756
rect 674340 623744 674346 623756
rect 676030 623744 676036 623756
rect 674340 623716 676036 623744
rect 674340 623704 674346 623716
rect 676030 623704 676036 623716
rect 676088 623704 676094 623756
rect 42150 623432 42156 623484
rect 42208 623472 42214 623484
rect 42886 623472 42892 623484
rect 42208 623444 42892 623472
rect 42208 623432 42214 623444
rect 42886 623432 42892 623444
rect 42944 623432 42950 623484
rect 42058 622140 42064 622192
rect 42116 622180 42122 622192
rect 42518 622180 42524 622192
rect 42116 622152 42524 622180
rect 42116 622140 42122 622152
rect 42518 622140 42524 622152
rect 42576 622140 42582 622192
rect 42150 621460 42156 621512
rect 42208 621500 42214 621512
rect 43346 621500 43352 621512
rect 42208 621472 43352 621500
rect 42208 621460 42214 621472
rect 43346 621460 43352 621472
rect 43404 621460 43410 621512
rect 670510 621052 670516 621104
rect 670568 621092 670574 621104
rect 676214 621092 676220 621104
rect 670568 621064 676220 621092
rect 670568 621052 670574 621064
rect 676214 621052 676220 621064
rect 676272 621052 676278 621104
rect 42058 620984 42064 621036
rect 42116 621024 42122 621036
rect 43254 621024 43260 621036
rect 42116 620996 43260 621024
rect 42116 620984 42122 620996
rect 43254 620984 43260 620996
rect 43312 620984 43318 621036
rect 670418 620984 670424 621036
rect 670476 621024 670482 621036
rect 678974 621024 678980 621036
rect 670476 620996 678980 621024
rect 670476 620984 670482 620996
rect 678974 620984 678980 620996
rect 679032 620984 679038 621036
rect 673822 620916 673828 620968
rect 673880 620956 673886 620968
rect 676030 620956 676036 620968
rect 673880 620928 676036 620956
rect 673880 620916 673886 620928
rect 676030 620916 676036 620928
rect 676088 620916 676094 620968
rect 673638 620848 673644 620900
rect 673696 620888 673702 620900
rect 676122 620888 676128 620900
rect 673696 620860 676128 620888
rect 673696 620848 673702 620860
rect 676122 620848 676128 620860
rect 676180 620848 676186 620900
rect 42058 620168 42064 620220
rect 42116 620208 42122 620220
rect 43438 620208 43444 620220
rect 42116 620180 43444 620208
rect 42116 620168 42122 620180
rect 43438 620168 43444 620180
rect 43496 620168 43502 620220
rect 42242 619012 42248 619064
rect 42300 619052 42306 619064
rect 43162 619052 43168 619064
rect 42300 619024 43168 619052
rect 42300 619012 42306 619024
rect 43162 619012 43168 619024
rect 43220 619012 43226 619064
rect 673270 618196 673276 618248
rect 673328 618236 673334 618248
rect 676030 618236 676036 618248
rect 673328 618208 676036 618236
rect 673328 618196 673334 618208
rect 676030 618196 676036 618208
rect 676088 618196 676094 618248
rect 673178 617924 673184 617976
rect 673236 617964 673242 617976
rect 676214 617964 676220 617976
rect 673236 617936 676220 617964
rect 673236 617924 673242 617936
rect 676214 617924 676220 617936
rect 676272 617924 676278 617976
rect 42150 617856 42156 617908
rect 42208 617896 42214 617908
rect 43622 617896 43628 617908
rect 42208 617868 43628 617896
rect 42208 617856 42214 617868
rect 43622 617856 43628 617868
rect 43680 617856 43686 617908
rect 42058 617108 42064 617160
rect 42116 617148 42122 617160
rect 43806 617148 43812 617160
rect 42116 617120 43812 617148
rect 42116 617108 42122 617120
rect 43806 617108 43812 617120
rect 43864 617108 43870 617160
rect 672994 616700 673000 616752
rect 673052 616740 673058 616752
rect 676214 616740 676220 616752
rect 673052 616712 676220 616740
rect 673052 616700 673058 616712
rect 676214 616700 676220 616712
rect 676272 616700 676278 616752
rect 42150 616632 42156 616684
rect 42208 616672 42214 616684
rect 43714 616672 43720 616684
rect 42208 616644 43720 616672
rect 42208 616632 42214 616644
rect 43714 616632 43720 616644
rect 43772 616632 43778 616684
rect 672442 614728 672448 614780
rect 672500 614768 672506 614780
rect 679250 614768 679256 614780
rect 672500 614740 679256 614768
rect 672500 614728 672506 614740
rect 679250 614728 679256 614740
rect 679308 614728 679314 614780
rect 42150 614184 42156 614236
rect 42208 614224 42214 614236
rect 43070 614224 43076 614236
rect 42208 614196 43076 614224
rect 42208 614184 42214 614196
rect 43070 614184 43076 614196
rect 43128 614184 43134 614236
rect 42150 613640 42156 613692
rect 42208 613680 42214 613692
rect 42978 613680 42984 613692
rect 42208 613652 42984 613680
rect 42208 613640 42214 613652
rect 42978 613640 42984 613652
rect 43036 613640 43042 613692
rect 42150 612960 42156 613012
rect 42208 613000 42214 613012
rect 42794 613000 42800 613012
rect 42208 612972 42800 613000
rect 42208 612960 42214 612972
rect 42794 612960 42800 612972
rect 42852 612960 42858 613012
rect 50982 609968 50988 610020
rect 51040 610008 51046 610020
rect 58434 610008 58440 610020
rect 51040 609980 58440 610008
rect 51040 609968 51046 609980
rect 58434 609968 58440 609980
rect 58492 609968 58498 610020
rect 674374 608744 674380 608796
rect 674432 608784 674438 608796
rect 675662 608784 675668 608796
rect 674432 608756 675668 608784
rect 674432 608744 674438 608756
rect 675662 608744 675668 608756
rect 675720 608744 675726 608796
rect 654594 603032 654600 603084
rect 654652 603072 654658 603084
rect 674558 603072 674564 603084
rect 654652 603044 674564 603072
rect 654652 603032 654658 603044
rect 674558 603032 674564 603044
rect 674616 603032 674622 603084
rect 654318 602148 654324 602200
rect 654376 602188 654382 602200
rect 661034 602188 661040 602200
rect 654376 602160 661040 602188
rect 654376 602148 654382 602160
rect 661034 602148 661040 602160
rect 661092 602148 661098 602200
rect 41506 601876 41512 601928
rect 41564 601916 41570 601928
rect 48866 601916 48872 601928
rect 41564 601888 48872 601916
rect 41564 601876 41570 601888
rect 48866 601876 48872 601888
rect 48924 601876 48930 601928
rect 41506 601468 41512 601520
rect 41564 601508 41570 601520
rect 51074 601508 51080 601520
rect 41564 601480 51080 601508
rect 41564 601468 41570 601480
rect 51074 601468 51080 601480
rect 51132 601468 51138 601520
rect 674282 600380 674288 600432
rect 674340 600420 674346 600432
rect 675478 600420 675484 600432
rect 674340 600392 675484 600420
rect 674340 600380 674346 600392
rect 675478 600380 675484 600392
rect 675536 600380 675542 600432
rect 41506 599836 41512 599888
rect 41564 599876 41570 599888
rect 44450 599876 44456 599888
rect 41564 599848 44456 599876
rect 41564 599836 41570 599848
rect 44450 599836 44456 599848
rect 44508 599836 44514 599888
rect 674742 599564 674748 599616
rect 674800 599604 674806 599616
rect 675478 599604 675484 599616
rect 674800 599576 675484 599604
rect 674800 599564 674806 599576
rect 675478 599564 675484 599576
rect 675536 599564 675542 599616
rect 673730 599088 673736 599140
rect 673788 599128 673794 599140
rect 675386 599128 675392 599140
rect 673788 599100 675392 599128
rect 673788 599088 673794 599100
rect 675386 599088 675392 599100
rect 675444 599088 675450 599140
rect 41506 598952 41512 599004
rect 41564 598992 41570 599004
rect 43346 598992 43352 599004
rect 41564 598964 43352 598992
rect 41564 598952 41570 598964
rect 43346 598952 43352 598964
rect 43404 598952 43410 599004
rect 673638 598408 673644 598460
rect 673696 598448 673702 598460
rect 675478 598448 675484 598460
rect 673696 598420 675484 598448
rect 673696 598408 673702 598420
rect 675478 598408 675484 598420
rect 675536 598408 675542 598460
rect 673822 597116 673828 597168
rect 673880 597156 673886 597168
rect 675386 597156 675392 597168
rect 673880 597128 675392 597156
rect 673880 597116 673886 597128
rect 675386 597116 675392 597128
rect 675444 597116 675450 597168
rect 674558 596844 674564 596896
rect 674616 596884 674622 596896
rect 675386 596884 675392 596896
rect 674616 596856 675392 596884
rect 674616 596844 674622 596856
rect 675386 596844 675392 596856
rect 675444 596844 675450 596896
rect 674466 596776 674472 596828
rect 674524 596776 674530 596828
rect 674484 596624 674512 596776
rect 674466 596572 674472 596624
rect 674524 596572 674530 596624
rect 53742 596164 53748 596216
rect 53800 596204 53806 596216
rect 59170 596204 59176 596216
rect 53800 596176 59176 596204
rect 53800 596164 53806 596176
rect 59170 596164 59176 596176
rect 59228 596164 59234 596216
rect 674374 595280 674380 595332
rect 674432 595320 674438 595332
rect 675386 595320 675392 595332
rect 674432 595292 675392 595320
rect 674432 595280 674438 595292
rect 675386 595280 675392 595292
rect 675444 595280 675450 595332
rect 675202 593648 675208 593700
rect 675260 593688 675266 593700
rect 675478 593688 675484 593700
rect 675260 593660 675484 593688
rect 675260 593648 675266 593660
rect 675478 593648 675484 593660
rect 675536 593648 675542 593700
rect 674558 593036 674564 593088
rect 674616 593076 674622 593088
rect 675570 593076 675576 593088
rect 674616 593048 675576 593076
rect 674616 593036 674622 593048
rect 675570 593036 675576 593048
rect 675628 593036 675634 593088
rect 43438 592560 43444 592612
rect 43496 592600 43502 592612
rect 43990 592600 43996 592612
rect 43496 592572 43996 592600
rect 43496 592560 43502 592572
rect 43990 592560 43996 592572
rect 44048 592560 44054 592612
rect 43254 592424 43260 592476
rect 43312 592464 43318 592476
rect 43438 592464 43444 592476
rect 43312 592436 43444 592464
rect 43312 592424 43318 592436
rect 43438 592424 43444 592436
rect 43496 592424 43502 592476
rect 656802 590656 656808 590708
rect 656860 590696 656866 590708
rect 669038 590696 669044 590708
rect 656860 590668 669044 590696
rect 656860 590656 656866 590668
rect 669038 590656 669044 590668
rect 669096 590656 669102 590708
rect 673362 587868 673368 587920
rect 673420 587908 673426 587920
rect 678974 587908 678980 587920
rect 673420 587880 678980 587908
rect 673420 587868 673426 587880
rect 678974 587868 678980 587880
rect 679032 587868 679038 587920
rect 41322 585148 41328 585200
rect 41380 585188 41386 585200
rect 44082 585188 44088 585200
rect 41380 585160 44088 585188
rect 41380 585148 41386 585160
rect 44082 585148 44088 585160
rect 44140 585148 44146 585200
rect 44174 585148 44180 585200
rect 44232 585188 44238 585200
rect 48958 585188 48964 585200
rect 44232 585160 48964 585188
rect 44232 585148 44238 585160
rect 48958 585148 48964 585160
rect 49016 585148 49022 585200
rect 41874 584196 41880 584248
rect 41932 584196 41938 584248
rect 41892 583976 41920 584196
rect 703446 584128 703452 584180
rect 703504 584168 703510 584180
rect 709334 584168 709340 584180
rect 703504 584140 709340 584168
rect 703504 584128 703510 584140
rect 709334 584128 709340 584140
rect 709392 584128 709398 584180
rect 41874 583924 41880 583976
rect 41932 583924 41938 583976
rect 674374 583924 674380 583976
rect 674432 583964 674438 583976
rect 674558 583964 674564 583976
rect 674432 583936 674564 583964
rect 674432 583924 674438 583936
rect 674558 583924 674564 583936
rect 674616 583924 674622 583976
rect 674650 583924 674656 583976
rect 674708 583964 674714 583976
rect 675386 583964 675392 583976
rect 674708 583936 675392 583964
rect 674708 583924 674714 583936
rect 675386 583924 675392 583936
rect 675444 583924 675450 583976
rect 43162 583856 43168 583908
rect 43220 583896 43226 583908
rect 43438 583896 43444 583908
rect 43220 583868 43444 583896
rect 43220 583856 43226 583868
rect 43438 583856 43444 583868
rect 43496 583856 43502 583908
rect 673822 583856 673828 583908
rect 673880 583896 673886 583908
rect 673880 583868 674420 583896
rect 673880 583856 673886 583868
rect 673638 583720 673644 583772
rect 673696 583760 673702 583772
rect 673822 583760 673828 583772
rect 673696 583732 673828 583760
rect 673696 583720 673702 583732
rect 673822 583720 673828 583732
rect 673880 583720 673886 583772
rect 674392 583704 674420 583868
rect 674742 583720 674748 583772
rect 674800 583760 674806 583772
rect 675478 583760 675484 583772
rect 674800 583732 675484 583760
rect 674800 583720 674806 583732
rect 675478 583720 675484 583732
rect 675536 583720 675542 583772
rect 42426 583652 42432 583704
rect 42484 583692 42490 583704
rect 43254 583692 43260 583704
rect 42484 583664 43260 583692
rect 42484 583652 42490 583664
rect 43254 583652 43260 583664
rect 43312 583652 43318 583704
rect 674374 583652 674380 583704
rect 674432 583652 674438 583704
rect 674558 583652 674564 583704
rect 674616 583692 674622 583704
rect 675202 583692 675208 583704
rect 674616 583664 675208 583692
rect 674616 583652 674622 583664
rect 675202 583652 675208 583664
rect 675260 583652 675266 583704
rect 48958 582360 48964 582412
rect 49016 582400 49022 582412
rect 58434 582400 58440 582412
rect 49016 582372 58440 582400
rect 49016 582360 49022 582372
rect 58434 582360 58440 582372
rect 58492 582360 58498 582412
rect 42150 582088 42156 582140
rect 42208 582128 42214 582140
rect 42886 582128 42892 582140
rect 42208 582100 42892 582128
rect 42208 582088 42214 582100
rect 42886 582088 42892 582100
rect 42944 582088 42950 582140
rect 703998 582088 704004 582140
rect 704056 582128 704062 582140
rect 708874 582128 708880 582140
rect 704056 582100 708880 582128
rect 704056 582088 704062 582100
rect 708874 582088 708880 582100
rect 708932 582088 708938 582140
rect 708046 582060 708052 582072
rect 704844 582032 708052 582060
rect 704844 581936 704872 582032
rect 708046 582020 708052 582032
rect 708104 582020 708110 582072
rect 704918 581952 704924 582004
rect 704976 581992 704982 582004
rect 707954 581992 707960 582004
rect 704976 581964 707960 581992
rect 704976 581952 704982 581964
rect 707954 581952 707960 581964
rect 708012 581952 708018 582004
rect 704826 581884 704832 581936
rect 704884 581884 704890 581936
rect 707034 581924 707040 581936
rect 705764 581896 707040 581924
rect 705764 581800 705792 581896
rect 707034 581884 707040 581896
rect 707092 581884 707098 581936
rect 706666 581856 706672 581868
rect 706224 581828 706672 581856
rect 706224 581800 706252 581828
rect 706666 581816 706672 581828
rect 706724 581816 706730 581868
rect 705746 581748 705752 581800
rect 705804 581748 705810 581800
rect 706206 581748 706212 581800
rect 706264 581748 706270 581800
rect 706298 581748 706304 581800
rect 706356 581788 706362 581800
rect 706574 581788 706580 581800
rect 706356 581760 706580 581788
rect 706356 581748 706362 581760
rect 706574 581748 706580 581760
rect 706632 581748 706638 581800
rect 705838 581680 705844 581732
rect 705896 581720 705902 581732
rect 707034 581720 707040 581732
rect 705896 581692 707040 581720
rect 705896 581680 705902 581692
rect 707034 581680 707040 581692
rect 707092 581680 707098 581732
rect 707586 581680 707592 581732
rect 707644 581680 707650 581732
rect 705378 581612 705384 581664
rect 705436 581652 705442 581664
rect 707494 581652 707500 581664
rect 705436 581624 707500 581652
rect 705436 581612 705442 581624
rect 707494 581612 707500 581624
rect 707552 581612 707558 581664
rect 705286 581544 705292 581596
rect 705344 581584 705350 581596
rect 707604 581584 707632 581680
rect 705344 581556 707632 581584
rect 705344 581544 705350 581556
rect 708506 581544 708512 581596
rect 708564 581544 708570 581596
rect 704458 581476 704464 581528
rect 704516 581516 704522 581528
rect 708414 581516 708420 581528
rect 704516 581488 708420 581516
rect 704516 581476 704522 581488
rect 708414 581476 708420 581488
rect 708472 581476 708478 581528
rect 704366 581408 704372 581460
rect 704424 581448 704430 581460
rect 708524 581448 708552 581544
rect 704424 581420 708552 581448
rect 704424 581408 704430 581420
rect 42150 581272 42156 581324
rect 42208 581312 42214 581324
rect 44174 581312 44180 581324
rect 42208 581284 44180 581312
rect 42208 581272 42214 581284
rect 44174 581272 44180 581284
rect 44232 581272 44238 581324
rect 42150 580252 42156 580304
rect 42208 580292 42214 580304
rect 42794 580292 42800 580304
rect 42208 580264 42800 580292
rect 42208 580252 42214 580264
rect 42794 580252 42800 580264
rect 42852 580252 42858 580304
rect 670234 580184 670240 580236
rect 670292 580224 670298 580236
rect 676030 580224 676036 580236
rect 670292 580196 676036 580224
rect 670292 580184 670298 580196
rect 676030 580184 676036 580196
rect 676088 580184 676094 580236
rect 669130 580048 669136 580100
rect 669188 580088 669194 580100
rect 676214 580088 676220 580100
rect 669188 580060 676220 580088
rect 669188 580048 669194 580060
rect 676214 580048 676220 580060
rect 676272 580048 676278 580100
rect 663794 579912 663800 579964
rect 663852 579952 663858 579964
rect 676122 579952 676128 579964
rect 663852 579924 676128 579952
rect 663852 579912 663858 579924
rect 676122 579912 676128 579924
rect 676180 579912 676186 579964
rect 660942 579776 660948 579828
rect 661000 579816 661006 579828
rect 676306 579816 676312 579828
rect 661000 579788 676312 579816
rect 661000 579776 661006 579788
rect 676306 579776 676312 579788
rect 676364 579776 676370 579828
rect 672534 579232 672540 579284
rect 672592 579272 672598 579284
rect 673270 579272 673276 579284
rect 672592 579244 673276 579272
rect 672592 579232 672598 579244
rect 673270 579232 673276 579244
rect 673328 579272 673334 579284
rect 676214 579272 676220 579284
rect 673328 579244 676220 579272
rect 673328 579232 673334 579244
rect 676214 579232 676220 579244
rect 676272 579232 676278 579284
rect 42150 578960 42156 579012
rect 42208 579000 42214 579012
rect 42702 579000 42708 579012
rect 42208 578972 42708 579000
rect 42208 578960 42214 578972
rect 42702 578960 42708 578972
rect 42760 578960 42766 579012
rect 42150 578416 42156 578468
rect 42208 578456 42214 578468
rect 43622 578456 43628 578468
rect 42208 578428 43628 578456
rect 42208 578416 42214 578428
rect 43622 578416 43628 578428
rect 43680 578416 43686 578468
rect 673086 578416 673092 578468
rect 673144 578456 673150 578468
rect 676214 578456 676220 578468
rect 673144 578428 676220 578456
rect 673144 578416 673150 578428
rect 676214 578416 676220 578428
rect 676272 578416 676278 578468
rect 42150 577804 42156 577856
rect 42208 577844 42214 577856
rect 43162 577844 43168 577856
rect 42208 577816 43168 577844
rect 42208 577804 42214 577816
rect 43162 577804 43168 577816
rect 43220 577804 43226 577856
rect 672718 577600 672724 577652
rect 672776 577640 672782 577652
rect 673178 577640 673184 577652
rect 672776 577612 673184 577640
rect 672776 577600 672782 577612
rect 673178 577600 673184 577612
rect 673236 577640 673242 577652
rect 676214 577640 676220 577652
rect 673236 577612 676220 577640
rect 673236 577600 673242 577612
rect 676214 577600 676220 577612
rect 676272 577600 676278 577652
rect 670510 577124 670516 577176
rect 670568 577164 670574 577176
rect 676214 577164 676220 577176
rect 670568 577136 676220 577164
rect 670568 577124 670574 577136
rect 676214 577124 676220 577136
rect 676272 577124 676278 577176
rect 42150 576920 42156 576972
rect 42208 576960 42214 576972
rect 43990 576960 43996 576972
rect 42208 576932 43996 576960
rect 42208 576920 42214 576932
rect 43990 576920 43996 576932
rect 44048 576920 44054 576972
rect 673362 576920 673368 576972
rect 673420 576960 673426 576972
rect 676030 576960 676036 576972
rect 673420 576932 676036 576960
rect 673420 576920 673426 576932
rect 676030 576920 676036 576932
rect 676088 576920 676094 576972
rect 654502 576852 654508 576904
rect 654560 576892 654566 576904
rect 663886 576892 663892 576904
rect 654560 576864 663892 576892
rect 654560 576852 654566 576864
rect 663886 576852 663892 576864
rect 663944 576852 663950 576904
rect 674466 576784 674472 576836
rect 674524 576824 674530 576836
rect 676030 576824 676036 576836
rect 674524 576796 676036 576824
rect 674524 576784 674530 576796
rect 676030 576784 676036 576796
rect 676088 576784 676094 576836
rect 674006 576036 674012 576088
rect 674064 576076 674070 576088
rect 676030 576076 676036 576088
rect 674064 576048 676036 576076
rect 674064 576036 674070 576048
rect 676030 576036 676036 576048
rect 676088 576036 676094 576088
rect 42150 574676 42156 574728
rect 42208 574716 42214 574728
rect 43714 574716 43720 574728
rect 42208 574688 43720 574716
rect 42208 574676 42214 574688
rect 43714 574676 43720 574688
rect 43772 574676 43778 574728
rect 42150 574064 42156 574116
rect 42208 574104 42214 574116
rect 42978 574104 42984 574116
rect 42208 574076 42984 574104
rect 42208 574064 42214 574076
rect 42978 574064 42984 574076
rect 43036 574064 43042 574116
rect 674190 573588 674196 573640
rect 674248 573628 674254 573640
rect 676030 573628 676036 573640
rect 674248 573600 676036 573628
rect 674248 573588 674254 573600
rect 676030 573588 676036 573600
rect 676088 573588 676094 573640
rect 42150 573452 42156 573504
rect 42208 573492 42214 573504
rect 44082 573492 44088 573504
rect 42208 573464 44088 573492
rect 42208 573452 42214 573464
rect 44082 573452 44088 573464
rect 44140 573452 44146 573504
rect 42058 572840 42064 572892
rect 42116 572880 42122 572892
rect 43898 572880 43904 572892
rect 42116 572852 43904 572880
rect 42116 572840 42122 572852
rect 43898 572840 43904 572852
rect 43956 572840 43962 572892
rect 673914 572772 673920 572824
rect 673972 572812 673978 572824
rect 676030 572812 676036 572824
rect 673972 572784 676036 572812
rect 673972 572772 673978 572784
rect 676030 572772 676036 572784
rect 676088 572772 676094 572824
rect 673546 572364 673552 572416
rect 673604 572404 673610 572416
rect 676030 572404 676036 572416
rect 673604 572376 676036 572404
rect 673604 572364 673610 572376
rect 676030 572364 676036 572376
rect 676088 572364 676094 572416
rect 42058 570868 42064 570920
rect 42116 570908 42122 570920
rect 43806 570908 43812 570920
rect 42116 570880 43812 570908
rect 42116 570868 42122 570880
rect 43806 570868 43812 570880
rect 43864 570868 43870 570920
rect 42150 570392 42156 570444
rect 42208 570432 42214 570444
rect 43438 570432 43444 570444
rect 42208 570404 43444 570432
rect 42208 570392 42214 570404
rect 43438 570392 43444 570404
rect 43496 570392 43502 570444
rect 42058 569576 42064 569628
rect 42116 569616 42122 569628
rect 43530 569616 43536 569628
rect 42116 569588 43536 569616
rect 42116 569576 42122 569588
rect 43530 569576 43536 569588
rect 43588 569576 43594 569628
rect 672534 568556 672540 568608
rect 672592 568596 672598 568608
rect 678974 568596 678980 568608
rect 672592 568568 678980 568596
rect 672592 568556 672598 568568
rect 678974 568556 678980 568568
rect 679032 568556 679038 568608
rect 673546 559512 673552 559564
rect 673604 559552 673610 559564
rect 675478 559552 675484 559564
rect 673604 559524 675484 559552
rect 673604 559512 673610 559524
rect 675478 559512 675484 559524
rect 675536 559512 675542 559564
rect 41506 558764 41512 558816
rect 41564 558804 41570 558816
rect 48958 558804 48964 558816
rect 41564 558776 48964 558804
rect 41564 558764 41570 558776
rect 48958 558764 48964 558776
rect 49016 558764 49022 558816
rect 41506 558288 41512 558340
rect 41564 558328 41570 558340
rect 53742 558328 53748 558340
rect 41564 558300 53748 558328
rect 41564 558288 41570 558300
rect 53742 558288 53748 558300
rect 53800 558288 53806 558340
rect 41782 558220 41788 558272
rect 41840 558260 41846 558272
rect 58434 558260 58440 558272
rect 41840 558232 58440 558260
rect 41840 558220 41846 558232
rect 58434 558220 58440 558232
rect 58492 558220 58498 558272
rect 49050 557540 49056 557592
rect 49108 557580 49114 557592
rect 57974 557580 57980 557592
rect 49108 557552 57980 557580
rect 49108 557540 49114 557552
rect 57974 557540 57980 557552
rect 58032 557540 58038 557592
rect 654318 556112 654324 556164
rect 654376 556152 654382 556164
rect 675294 556152 675300 556164
rect 654376 556124 675300 556152
rect 654376 556112 654382 556124
rect 675294 556112 675300 556124
rect 675352 556112 675358 556164
rect 674190 555228 674196 555280
rect 674248 555268 674254 555280
rect 675386 555268 675392 555280
rect 674248 555240 675392 555268
rect 674248 555228 674254 555240
rect 675386 555228 675392 555240
rect 675444 555228 675450 555280
rect 673454 554548 673460 554600
rect 673512 554588 673518 554600
rect 675386 554588 675392 554600
rect 673512 554560 675392 554588
rect 673512 554548 673518 554560
rect 675386 554548 675392 554560
rect 675444 554548 675450 554600
rect 673914 553732 673920 553784
rect 673972 553772 673978 553784
rect 675386 553772 675392 553784
rect 673972 553744 675392 553772
rect 673972 553732 673978 553744
rect 675386 553732 675392 553744
rect 675444 553732 675450 553784
rect 673638 553188 673644 553240
rect 673696 553228 673702 553240
rect 675386 553228 675392 553240
rect 673696 553200 675392 553228
rect 673696 553188 673702 553200
rect 675386 553188 675392 553200
rect 675444 553188 675450 553240
rect 674006 551896 674012 551948
rect 674064 551936 674070 551948
rect 675386 551936 675392 551948
rect 674064 551908 675392 551936
rect 674064 551896 674070 551908
rect 675386 551896 675392 551908
rect 675444 551896 675450 551948
rect 655054 550196 655060 550248
rect 655112 550236 655118 550248
rect 669130 550236 669136 550248
rect 655112 550208 669136 550236
rect 655112 550196 655118 550208
rect 669130 550196 669136 550208
rect 669188 550196 669194 550248
rect 674466 548836 674472 548888
rect 674524 548876 674530 548888
rect 675294 548876 675300 548888
rect 674524 548848 675300 548876
rect 674524 548836 674530 548848
rect 675294 548836 675300 548848
rect 675352 548836 675358 548888
rect 674650 548224 674656 548276
rect 674708 548264 674714 548276
rect 675294 548264 675300 548276
rect 674708 548236 675300 548264
rect 674708 548224 674714 548236
rect 675294 548224 675300 548236
rect 675352 548224 675358 548276
rect 41414 547272 41420 547324
rect 41472 547312 41478 547324
rect 48958 547312 48964 547324
rect 41472 547284 48964 547312
rect 41472 547272 41478 547284
rect 48958 547272 48964 547284
rect 49016 547272 49022 547324
rect 673086 546252 673092 546304
rect 673144 546292 673150 546304
rect 679066 546292 679072 546304
rect 673144 546264 679072 546292
rect 673144 546252 673150 546264
rect 679066 546252 679072 546264
rect 679124 546252 679130 546304
rect 53834 543736 53840 543788
rect 53892 543776 53898 543788
rect 59170 543776 59176 543788
rect 53892 543748 59176 543776
rect 53892 543736 53898 543748
rect 59170 543736 59176 543748
rect 59228 543736 59234 543788
rect 41598 543124 41604 543176
rect 41656 543164 41662 543176
rect 43254 543164 43260 543176
rect 41656 543136 43260 543164
rect 41656 543124 41662 543136
rect 43254 543124 43260 543136
rect 43312 543124 43318 543176
rect 41506 542444 41512 542496
rect 41564 542484 41570 542496
rect 42794 542484 42800 542496
rect 41564 542456 42800 542484
rect 41564 542444 41570 542456
rect 42794 542444 42800 542456
rect 42852 542444 42858 542496
rect 41782 541016 41788 541068
rect 41840 541016 41846 541068
rect 43898 541016 43904 541068
rect 43956 541056 43962 541068
rect 50982 541056 50988 541068
rect 43956 541028 50988 541056
rect 43956 541016 43962 541028
rect 50982 541016 50988 541028
rect 51040 541016 51046 541068
rect 41800 540796 41828 541016
rect 41782 540744 41788 540796
rect 41840 540744 41846 540796
rect 42058 538908 42064 538960
rect 42116 538948 42122 538960
rect 42702 538948 42708 538960
rect 42116 538920 42708 538948
rect 42116 538908 42122 538920
rect 42702 538908 42708 538920
rect 42760 538908 42766 538960
rect 42150 538092 42156 538144
rect 42208 538132 42214 538144
rect 43898 538132 43904 538144
rect 42208 538104 43904 538132
rect 42208 538092 42214 538104
rect 43898 538092 43904 538104
rect 43956 538092 43962 538144
rect 703446 537140 703452 537192
rect 703504 537180 703510 537192
rect 703504 537152 709012 537180
rect 703504 537140 703510 537152
rect 708984 537124 709012 537152
rect 42058 537072 42064 537124
rect 42116 537112 42122 537124
rect 42886 537112 42892 537124
rect 42116 537084 42892 537112
rect 42116 537072 42122 537084
rect 42886 537072 42892 537084
rect 42944 537072 42950 537124
rect 703538 537072 703544 537124
rect 703596 537112 703602 537124
rect 708874 537112 708880 537124
rect 703596 537084 708880 537112
rect 703596 537072 703602 537084
rect 708874 537072 708880 537084
rect 708932 537072 708938 537124
rect 708966 537072 708972 537124
rect 709024 537072 709030 537124
rect 708046 537044 708052 537056
rect 704844 537016 708052 537044
rect 704844 536920 704872 537016
rect 708046 537004 708052 537016
rect 708104 537004 708110 537056
rect 704918 536936 704924 536988
rect 704976 536976 704982 536988
rect 707954 536976 707960 536988
rect 704976 536948 707960 536976
rect 704976 536936 704982 536948
rect 707954 536936 707960 536948
rect 708012 536936 708018 536988
rect 42978 536868 42984 536920
rect 43036 536908 43042 536920
rect 43346 536908 43352 536920
rect 43036 536880 43352 536908
rect 43036 536868 43042 536880
rect 43346 536868 43352 536880
rect 43404 536868 43410 536920
rect 704826 536868 704832 536920
rect 704884 536868 704890 536920
rect 707034 536908 707040 536920
rect 705764 536880 707040 536908
rect 705764 536784 705792 536880
rect 707034 536868 707040 536880
rect 707092 536868 707098 536920
rect 706666 536840 706672 536852
rect 706224 536812 706672 536840
rect 706224 536784 706252 536812
rect 706666 536800 706672 536812
rect 706724 536800 706730 536852
rect 43346 536732 43352 536784
rect 43404 536772 43410 536784
rect 43530 536772 43536 536784
rect 43404 536744 43536 536772
rect 43404 536732 43410 536744
rect 43530 536732 43536 536744
rect 43588 536732 43594 536784
rect 705746 536732 705752 536784
rect 705804 536732 705810 536784
rect 706206 536732 706212 536784
rect 706264 536732 706270 536784
rect 706298 536732 706304 536784
rect 706356 536772 706362 536784
rect 706574 536772 706580 536784
rect 706356 536744 706580 536772
rect 706356 536732 706362 536744
rect 706574 536732 706580 536744
rect 706632 536732 706638 536784
rect 705838 536664 705844 536716
rect 705896 536704 705902 536716
rect 707034 536704 707040 536716
rect 705896 536676 707040 536704
rect 705896 536664 705902 536676
rect 707034 536664 707040 536676
rect 707092 536664 707098 536716
rect 707586 536664 707592 536716
rect 707644 536664 707650 536716
rect 705378 536596 705384 536648
rect 705436 536636 705442 536648
rect 707494 536636 707500 536648
rect 705436 536608 707500 536636
rect 705436 536596 705442 536608
rect 707494 536596 707500 536608
rect 707552 536596 707558 536648
rect 705286 536528 705292 536580
rect 705344 536568 705350 536580
rect 707604 536568 707632 536664
rect 705344 536540 707632 536568
rect 705344 536528 705350 536540
rect 708506 536528 708512 536580
rect 708564 536528 708570 536580
rect 704458 536460 704464 536512
rect 704516 536500 704522 536512
rect 708414 536500 708420 536512
rect 704516 536472 708420 536500
rect 704516 536460 704522 536472
rect 708414 536460 708420 536472
rect 708472 536460 708478 536512
rect 654686 536392 654692 536444
rect 654744 536432 654750 536444
rect 667106 536432 667112 536444
rect 654744 536404 667112 536432
rect 654744 536392 654750 536404
rect 667106 536392 667112 536404
rect 667164 536392 667170 536444
rect 704366 536392 704372 536444
rect 704424 536432 704430 536444
rect 708524 536432 708552 536528
rect 704424 536404 708552 536432
rect 704424 536392 704430 536404
rect 42150 535780 42156 535832
rect 42208 535820 42214 535832
rect 42794 535820 42800 535832
rect 42208 535792 42800 535820
rect 42208 535780 42214 535792
rect 42794 535780 42800 535792
rect 42852 535780 42858 535832
rect 666462 535712 666468 535764
rect 666520 535752 666526 535764
rect 676214 535752 676220 535764
rect 666520 535724 676220 535752
rect 666520 535712 666526 535724
rect 676214 535712 676220 535724
rect 676272 535712 676278 535764
rect 663702 535576 663708 535628
rect 663760 535616 663766 535628
rect 676030 535616 676036 535628
rect 663760 535588 676036 535616
rect 663760 535576 663766 535588
rect 676030 535576 676036 535588
rect 676088 535576 676094 535628
rect 42058 535032 42064 535084
rect 42116 535072 42122 535084
rect 43438 535072 43444 535084
rect 42116 535044 43444 535072
rect 42116 535032 42122 535044
rect 43438 535032 43444 535044
rect 43496 535032 43502 535084
rect 673270 534896 673276 534948
rect 673328 534936 673334 534948
rect 676030 534936 676036 534948
rect 673328 534908 676036 534936
rect 673328 534896 673334 534908
rect 676030 534896 676036 534908
rect 676088 534896 676094 534948
rect 42150 534556 42156 534608
rect 42208 534596 42214 534608
rect 43254 534596 43260 534608
rect 42208 534568 43260 534596
rect 42208 534556 42214 534568
rect 43254 534556 43260 534568
rect 43312 534556 43318 534608
rect 42150 533740 42156 533792
rect 42208 533780 42214 533792
rect 43162 533780 43168 533792
rect 42208 533752 43168 533780
rect 42208 533740 42214 533752
rect 43162 533740 43168 533752
rect 43220 533740 43226 533792
rect 673178 533264 673184 533316
rect 673236 533304 673242 533316
rect 676030 533304 676036 533316
rect 673236 533276 676036 533304
rect 673236 533264 673242 533276
rect 676030 533264 676036 533276
rect 676088 533264 676094 533316
rect 667198 532856 667204 532908
rect 667256 532896 667262 532908
rect 678974 532896 678980 532908
rect 667256 532868 678980 532896
rect 667256 532856 667262 532868
rect 678974 532856 678980 532868
rect 679032 532856 679038 532908
rect 670050 532788 670056 532840
rect 670108 532828 670114 532840
rect 675846 532828 675852 532840
rect 670108 532800 675852 532828
rect 670108 532788 670114 532800
rect 675846 532788 675852 532800
rect 675904 532828 675910 532840
rect 676122 532828 676128 532840
rect 675904 532800 676128 532828
rect 675904 532788 675910 532800
rect 676122 532788 676128 532800
rect 676180 532788 676186 532840
rect 674742 532652 674748 532704
rect 674800 532692 674806 532704
rect 676030 532692 676036 532704
rect 674800 532664 676036 532692
rect 674800 532652 674806 532664
rect 676030 532652 676036 532664
rect 676088 532652 676094 532704
rect 672810 532584 672816 532636
rect 672868 532624 672874 532636
rect 673362 532624 673368 532636
rect 672868 532596 673368 532624
rect 672868 532584 672874 532596
rect 673362 532584 673368 532596
rect 673420 532624 673426 532636
rect 676214 532624 676220 532636
rect 673420 532596 676220 532624
rect 673420 532584 673426 532596
rect 676214 532584 676220 532596
rect 676272 532584 676278 532636
rect 42150 531428 42156 531480
rect 42208 531468 42214 531480
rect 43806 531468 43812 531480
rect 42208 531440 43812 531468
rect 42208 531428 42214 531440
rect 43806 531428 43812 531440
rect 43864 531428 43870 531480
rect 674282 531088 674288 531140
rect 674340 531128 674346 531140
rect 676030 531128 676036 531140
rect 674340 531100 676036 531128
rect 674340 531088 674346 531100
rect 676030 531088 676036 531100
rect 676088 531088 676094 531140
rect 42150 530680 42156 530732
rect 42208 530720 42214 530732
rect 43714 530720 43720 530732
rect 42208 530692 43720 530720
rect 42208 530680 42214 530692
rect 43714 530680 43720 530692
rect 43772 530680 43778 530732
rect 42150 530272 42156 530324
rect 42208 530312 42214 530324
rect 43070 530312 43076 530324
rect 42208 530284 43076 530312
rect 42208 530272 42214 530284
rect 43070 530272 43076 530284
rect 43128 530272 43134 530324
rect 674558 529864 674564 529916
rect 674616 529904 674622 529916
rect 676030 529904 676036 529916
rect 674616 529876 676036 529904
rect 674616 529864 674622 529876
rect 676030 529864 676036 529876
rect 676088 529864 676094 529916
rect 42150 529592 42156 529644
rect 42208 529632 42214 529644
rect 42886 529632 42892 529644
rect 42208 529604 42892 529632
rect 42208 529592 42214 529604
rect 42886 529592 42892 529604
rect 42944 529592 42950 529644
rect 674374 529456 674380 529508
rect 674432 529496 674438 529508
rect 676030 529496 676036 529508
rect 674432 529468 676036 529496
rect 674432 529456 674438 529468
rect 676030 529456 676036 529468
rect 676088 529456 676094 529508
rect 673730 527824 673736 527876
rect 673788 527864 673794 527876
rect 676030 527864 676036 527876
rect 673788 527836 676036 527864
rect 673788 527824 673794 527836
rect 676030 527824 676036 527836
rect 676088 527824 676094 527876
rect 42058 527212 42064 527264
rect 42116 527252 42122 527264
rect 43346 527252 43352 527264
rect 42116 527224 43352 527252
rect 42116 527212 42122 527224
rect 43346 527212 43352 527224
rect 43404 527212 43410 527264
rect 42150 527144 42156 527196
rect 42208 527184 42214 527196
rect 43622 527184 43628 527196
rect 42208 527156 43628 527184
rect 42208 527144 42214 527156
rect 43622 527144 43628 527156
rect 43680 527144 43686 527196
rect 673822 527076 673828 527128
rect 673880 527116 673886 527128
rect 676030 527116 676036 527128
rect 673880 527088 676036 527116
rect 673880 527076 673886 527088
rect 676030 527076 676036 527088
rect 676088 527076 676094 527128
rect 42150 526600 42156 526652
rect 42208 526640 42214 526652
rect 42978 526640 42984 526652
rect 42208 526612 42984 526640
rect 42208 526600 42214 526612
rect 42978 526600 42984 526612
rect 43036 526600 43042 526652
rect 672626 524424 672632 524476
rect 672684 524464 672690 524476
rect 678974 524464 678980 524476
rect 672684 524436 678980 524464
rect 672684 524424 672690 524436
rect 678974 524424 678980 524436
rect 679032 524424 679038 524476
rect 677502 524356 677508 524408
rect 677560 524396 677566 524408
rect 679066 524396 679072 524408
rect 677560 524368 679072 524396
rect 677560 524356 677566 524368
rect 679066 524356 679072 524368
rect 679124 524356 679130 524408
rect 654134 522452 654140 522504
rect 654192 522492 654198 522504
rect 661218 522492 661224 522504
rect 654192 522464 661224 522492
rect 654192 522452 654198 522464
rect 661218 522452 661224 522464
rect 661276 522452 661282 522504
rect 51258 518916 51264 518968
rect 51316 518956 51322 518968
rect 58434 518956 58440 518968
rect 51316 518928 58440 518956
rect 51316 518916 51322 518928
rect 58434 518916 58440 518928
rect 58492 518916 58498 518968
rect 654778 510620 654784 510672
rect 654836 510660 654842 510672
rect 667014 510660 667020 510672
rect 654836 510632 667020 510660
rect 654836 510620 654842 510632
rect 667014 510620 667020 510632
rect 667072 510620 667078 510672
rect 50982 505112 50988 505164
rect 51040 505152 51046 505164
rect 58434 505152 58440 505164
rect 51040 505124 58440 505152
rect 51040 505112 51046 505124
rect 58434 505112 58440 505124
rect 58492 505112 58498 505164
rect 656802 497632 656808 497684
rect 656860 497672 656866 497684
rect 663794 497672 663800 497684
rect 656860 497644 663800 497672
rect 656860 497632 656866 497644
rect 663794 497632 663800 497644
rect 663852 497632 663858 497684
rect 704366 493076 704372 493128
rect 704424 493116 704430 493128
rect 704424 493088 708552 493116
rect 704424 493076 704430 493088
rect 704458 493008 704464 493060
rect 704516 493048 704522 493060
rect 708414 493048 708420 493060
rect 704516 493020 708420 493048
rect 704516 493008 704522 493020
rect 708414 493008 708420 493020
rect 708472 493008 708478 493060
rect 708524 492992 708552 493088
rect 705378 492940 705384 492992
rect 705436 492980 705442 492992
rect 705436 492952 707402 492980
rect 705436 492940 705442 492952
rect 707034 492912 707040 492924
rect 705764 492884 707040 492912
rect 705764 492856 705792 492884
rect 707034 492872 707040 492884
rect 707092 492872 707098 492924
rect 705746 492804 705752 492856
rect 705804 492804 705810 492856
rect 706206 492804 706212 492856
rect 706264 492844 706270 492856
rect 706574 492844 706580 492856
rect 706264 492816 706580 492844
rect 706264 492804 706270 492816
rect 706574 492804 706580 492816
rect 706632 492804 706638 492856
rect 707374 492844 707402 492952
rect 708506 492940 708512 492992
rect 708564 492940 708570 492992
rect 707586 492844 707592 492856
rect 707374 492816 707592 492844
rect 707586 492804 707592 492816
rect 707644 492804 707650 492856
rect 705838 492736 705844 492788
rect 705896 492776 705902 492788
rect 707034 492776 707040 492788
rect 705896 492748 707040 492776
rect 705896 492736 705902 492748
rect 707034 492736 707040 492748
rect 707092 492736 707098 492788
rect 706298 492668 706304 492720
rect 706356 492708 706362 492720
rect 706574 492708 706580 492720
rect 706356 492680 706580 492708
rect 706356 492668 706362 492680
rect 706574 492668 706580 492680
rect 706632 492668 706638 492720
rect 705378 492600 705384 492652
rect 705436 492640 705442 492652
rect 707494 492640 707500 492652
rect 705436 492612 707500 492640
rect 705436 492600 705442 492612
rect 707494 492600 707500 492612
rect 707552 492600 707558 492652
rect 704826 492532 704832 492584
rect 704884 492572 704890 492584
rect 707954 492572 707960 492584
rect 704884 492544 707960 492572
rect 704884 492532 704890 492544
rect 707954 492532 707960 492544
rect 708012 492532 708018 492584
rect 703906 492464 703912 492516
rect 703964 492504 703970 492516
rect 708874 492504 708880 492516
rect 703964 492476 708880 492504
rect 703964 492464 703970 492476
rect 708874 492464 708880 492476
rect 708932 492464 708938 492516
rect 704918 492396 704924 492448
rect 704976 492436 704982 492448
rect 707954 492436 707960 492448
rect 704976 492408 707960 492436
rect 704976 492396 704982 492408
rect 707954 492396 707960 492408
rect 708012 492396 708018 492448
rect 703538 492328 703544 492380
rect 703596 492368 703602 492380
rect 708874 492368 708880 492380
rect 703596 492340 708880 492368
rect 703596 492328 703602 492340
rect 708874 492328 708880 492340
rect 708932 492328 708938 492380
rect 669038 491648 669044 491700
rect 669096 491688 669102 491700
rect 676030 491688 676036 491700
rect 669096 491660 676036 491688
rect 669096 491648 669102 491660
rect 676030 491648 676036 491660
rect 676088 491648 676094 491700
rect 663886 491512 663892 491564
rect 663944 491552 663950 491564
rect 676030 491552 676036 491564
rect 663944 491524 676036 491552
rect 663944 491512 663950 491524
rect 676030 491512 676036 491524
rect 676088 491512 676094 491564
rect 661034 491376 661040 491428
rect 661092 491416 661098 491428
rect 675938 491416 675944 491428
rect 661092 491388 675944 491416
rect 661092 491376 661098 491388
rect 675938 491376 675944 491388
rect 675996 491376 676002 491428
rect 49142 491308 49148 491360
rect 49200 491348 49206 491360
rect 57974 491348 57980 491360
rect 49200 491320 57980 491348
rect 49200 491308 49206 491320
rect 57974 491308 57980 491320
rect 58032 491308 58038 491360
rect 676214 491240 676220 491292
rect 676272 491280 676278 491292
rect 677502 491280 677508 491292
rect 676272 491252 677508 491280
rect 676272 491240 676278 491252
rect 677502 491240 677508 491252
rect 677560 491240 677566 491292
rect 676122 490192 676128 490204
rect 676048 490164 676128 490192
rect 676048 490000 676076 490164
rect 676122 490152 676128 490164
rect 676180 490152 676186 490204
rect 676030 489948 676036 490000
rect 676088 489948 676094 490000
rect 669590 488520 669596 488572
rect 669648 488560 669654 488572
rect 675570 488560 675576 488572
rect 669648 488532 675576 488560
rect 669648 488520 669654 488532
rect 675570 488520 675576 488532
rect 675628 488560 675634 488572
rect 675938 488560 675944 488572
rect 675628 488532 675944 488560
rect 675628 488520 675634 488532
rect 675938 488520 675944 488532
rect 675996 488520 676002 488572
rect 669682 488044 669688 488096
rect 669740 488084 669746 488096
rect 675202 488084 675208 488096
rect 669740 488056 675208 488084
rect 669740 488044 669746 488056
rect 675202 488044 675208 488056
rect 675260 488044 675266 488096
rect 674466 487840 674472 487892
rect 674524 487880 674530 487892
rect 676030 487880 676036 487892
rect 674524 487852 676036 487880
rect 674524 487840 674530 487852
rect 676030 487840 676036 487852
rect 676088 487840 676094 487892
rect 673546 487432 673552 487484
rect 673604 487472 673610 487484
rect 675938 487472 675944 487484
rect 673604 487444 675944 487472
rect 673604 487432 673610 487444
rect 675938 487432 675944 487444
rect 675996 487432 676002 487484
rect 674190 487092 674196 487144
rect 674248 487132 674254 487144
rect 676030 487132 676036 487144
rect 674248 487104 676036 487132
rect 674248 487092 674254 487104
rect 676030 487092 676036 487104
rect 676088 487092 676094 487144
rect 674650 485732 674656 485784
rect 674708 485772 674714 485784
rect 676030 485772 676036 485784
rect 674708 485744 676036 485772
rect 674708 485732 674714 485744
rect 676030 485732 676036 485744
rect 676088 485732 676094 485784
rect 674006 485460 674012 485512
rect 674064 485500 674070 485512
rect 676030 485500 676036 485512
rect 674064 485472 676036 485500
rect 674064 485460 674070 485472
rect 676030 485460 676036 485472
rect 676088 485460 676094 485512
rect 673914 483828 673920 483880
rect 673972 483868 673978 483880
rect 676030 483868 676036 483880
rect 673972 483840 676036 483868
rect 673972 483828 673978 483840
rect 676030 483828 676036 483840
rect 676088 483828 676094 483880
rect 655054 483284 655060 483336
rect 655112 483324 655118 483336
rect 670050 483324 670056 483336
rect 655112 483296 670056 483324
rect 655112 483284 655118 483296
rect 670050 483284 670056 483296
rect 670108 483284 670114 483336
rect 673638 482944 673644 482996
rect 673696 482984 673702 482996
rect 676030 482984 676036 482996
rect 673696 482956 676036 482984
rect 673696 482944 673702 482956
rect 676030 482944 676036 482956
rect 676088 482944 676094 482996
rect 673454 482876 673460 482928
rect 673512 482916 673518 482928
rect 675938 482916 675944 482928
rect 673512 482888 675944 482916
rect 673512 482876 673518 482888
rect 675938 482876 675944 482888
rect 675996 482876 676002 482928
rect 676030 481148 676036 481160
rect 673426 481120 676036 481148
rect 672718 481040 672724 481092
rect 672776 481080 672782 481092
rect 673426 481080 673454 481120
rect 676030 481108 676036 481120
rect 676088 481108 676094 481160
rect 672776 481052 673454 481080
rect 672776 481040 672782 481052
rect 51166 480224 51172 480276
rect 51224 480264 51230 480276
rect 58434 480264 58440 480276
rect 51224 480236 58440 480264
rect 51224 480224 51230 480236
rect 58434 480224 58440 480236
rect 58492 480224 58498 480276
rect 675570 478864 675576 478916
rect 675628 478904 675634 478916
rect 676122 478904 676128 478916
rect 675628 478876 676128 478904
rect 675628 478864 675634 478876
rect 676122 478864 676128 478876
rect 676180 478864 676186 478916
rect 654870 470500 654876 470552
rect 654928 470540 654934 470552
rect 663702 470540 663708 470552
rect 654928 470512 663708 470540
rect 654928 470500 654934 470512
rect 663702 470500 663708 470512
rect 663760 470500 663766 470552
rect 54018 466420 54024 466472
rect 54076 466460 54082 466472
rect 58618 466460 58624 466472
rect 54076 466432 58624 466460
rect 54076 466420 54082 466432
rect 58618 466420 58624 466432
rect 58676 466420 58682 466472
rect 654134 457308 654140 457360
rect 654192 457348 654198 457360
rect 661034 457348 661040 457360
rect 654192 457320 661040 457348
rect 654192 457308 654198 457320
rect 661034 457308 661040 457320
rect 661092 457308 661098 457360
rect 53742 452616 53748 452668
rect 53800 452656 53806 452668
rect 59170 452656 59176 452668
rect 53800 452628 59176 452656
rect 53800 452616 53806 452628
rect 59170 452616 59176 452628
rect 59228 452616 59234 452668
rect 656802 444456 656808 444508
rect 656860 444496 656866 444508
rect 663886 444496 663892 444508
rect 656860 444468 663892 444496
rect 656860 444456 656866 444468
rect 663886 444456 663892 444468
rect 663944 444456 663950 444508
rect 51074 438880 51080 438932
rect 51132 438920 51138 438932
rect 58434 438920 58440 438932
rect 51132 438892 58440 438920
rect 51132 438880 51138 438892
rect 58434 438880 58440 438892
rect 58492 438880 58498 438932
rect 43990 430652 43996 430704
rect 44048 430692 44054 430704
rect 62390 430692 62396 430704
rect 44048 430664 62396 430692
rect 44048 430652 44054 430664
rect 62390 430652 62396 430664
rect 62448 430652 62454 430704
rect 41782 430584 41788 430636
rect 41840 430624 41846 430636
rect 59262 430624 59268 430636
rect 41840 430596 59268 430624
rect 41840 430584 41846 430596
rect 59262 430584 59268 430596
rect 59320 430584 59326 430636
rect 654870 430584 654876 430636
rect 654928 430624 654934 430636
rect 666462 430624 666468 430636
rect 654928 430596 666468 430624
rect 654928 430584 654934 430596
rect 666462 430584 666468 430596
rect 666520 430584 666526 430636
rect 53926 427864 53932 427916
rect 53984 427904 53990 427916
rect 57974 427904 57980 427916
rect 53984 427876 57980 427904
rect 53984 427864 53990 427876
rect 57974 427864 57980 427876
rect 58032 427864 58038 427916
rect 41782 427796 41788 427848
rect 41840 427836 41846 427848
rect 44082 427836 44088 427848
rect 41840 427808 44088 427836
rect 41840 427796 41846 427808
rect 44082 427796 44088 427808
rect 44140 427836 44146 427848
rect 62942 427836 62948 427848
rect 44140 427808 62948 427836
rect 44140 427796 44146 427808
rect 62942 427796 62948 427808
rect 63000 427796 63006 427848
rect 655054 417460 655060 417512
rect 655112 417500 655118 417512
rect 660942 417500 660948 417512
rect 655112 417472 660948 417500
rect 655112 417460 655118 417472
rect 660942 417460 660948 417472
rect 661000 417460 661006 417512
rect 41782 416304 41788 416356
rect 41840 416344 41846 416356
rect 43070 416344 43076 416356
rect 41840 416316 43076 416344
rect 41840 416304 41846 416316
rect 43070 416304 43076 416316
rect 43128 416304 43134 416356
rect 49234 413992 49240 414044
rect 49292 414032 49298 414044
rect 58434 414032 58440 414044
rect 49292 414004 58440 414032
rect 49292 413992 49298 414004
rect 58434 413992 58440 414004
rect 58492 413992 58498 414044
rect 41874 413380 41880 413432
rect 41932 413380 41938 413432
rect 41892 413160 41920 413380
rect 41874 413108 41880 413160
rect 41932 413108 41938 413160
rect 42794 411340 42800 411392
rect 42852 411340 42858 411392
rect 42150 411272 42156 411324
rect 42208 411312 42214 411324
rect 42812 411312 42840 411340
rect 42208 411284 42840 411312
rect 42208 411272 42214 411284
rect 42150 410660 42156 410712
rect 42208 410700 42214 410712
rect 49050 410700 49056 410712
rect 42208 410672 49056 410700
rect 42208 410660 42214 410672
rect 49050 410660 49056 410672
rect 49108 410660 49114 410712
rect 42150 409368 42156 409420
rect 42208 409408 42214 409420
rect 42978 409408 42984 409420
rect 42208 409380 42984 409408
rect 42208 409368 42214 409380
rect 42978 409368 42984 409380
rect 43036 409368 43042 409420
rect 42058 408144 42064 408196
rect 42116 408184 42122 408196
rect 42518 408184 42524 408196
rect 42116 408156 42524 408184
rect 42116 408144 42122 408156
rect 42518 408144 42524 408156
rect 42576 408144 42582 408196
rect 42150 407464 42156 407516
rect 42208 407504 42214 407516
rect 43346 407504 43352 407516
rect 42208 407476 43352 407504
rect 42208 407464 42214 407476
rect 43346 407464 43352 407476
rect 43404 407464 43410 407516
rect 42058 406988 42064 407040
rect 42116 407028 42122 407040
rect 43070 407028 43076 407040
rect 42116 407000 43076 407028
rect 42116 406988 42122 407000
rect 43070 406988 43076 407000
rect 43128 406988 43134 407040
rect 42150 406172 42156 406224
rect 42208 406212 42214 406224
rect 43438 406212 43444 406224
rect 42208 406184 43444 406212
rect 42208 406172 42214 406184
rect 43438 406172 43444 406184
rect 43496 406172 43502 406224
rect 703556 404960 709012 404988
rect 703556 404932 703584 404960
rect 708984 404932 709012 404960
rect 703538 404880 703544 404932
rect 703596 404880 703602 404932
rect 703998 404880 704004 404932
rect 704056 404920 704062 404932
rect 708874 404920 708880 404932
rect 704056 404892 708880 404920
rect 704056 404880 704062 404892
rect 708874 404880 708880 404892
rect 708932 404880 708938 404932
rect 708966 404880 708972 404932
rect 709024 404880 709030 404932
rect 708046 404852 708052 404864
rect 704844 404824 708052 404852
rect 704844 404728 704872 404824
rect 708046 404812 708052 404824
rect 708104 404812 708110 404864
rect 704918 404744 704924 404796
rect 704976 404784 704982 404796
rect 707954 404784 707960 404796
rect 704976 404756 707960 404784
rect 704976 404744 704982 404756
rect 707954 404744 707960 404756
rect 708012 404744 708018 404796
rect 704826 404676 704832 404728
rect 704884 404676 704890 404728
rect 707034 404716 707040 404728
rect 705856 404688 707040 404716
rect 705746 404540 705752 404592
rect 705804 404580 705810 404592
rect 705856 404580 705884 404688
rect 707034 404676 707040 404688
rect 707092 404676 707098 404728
rect 706666 404648 706672 404660
rect 706224 404620 706672 404648
rect 706224 404592 706252 404620
rect 706666 404608 706672 404620
rect 706724 404608 706730 404660
rect 705804 404552 705884 404580
rect 705804 404540 705810 404552
rect 706206 404540 706212 404592
rect 706264 404540 706270 404592
rect 706298 404540 706304 404592
rect 706356 404580 706362 404592
rect 706574 404580 706580 404592
rect 706356 404552 706580 404580
rect 706356 404540 706362 404552
rect 706574 404540 706580 404552
rect 706632 404540 706638 404592
rect 705838 404472 705844 404524
rect 705896 404512 705902 404524
rect 707034 404512 707040 404524
rect 705896 404484 707040 404512
rect 705896 404472 705902 404484
rect 707034 404472 707040 404484
rect 707092 404472 707098 404524
rect 707586 404472 707592 404524
rect 707644 404472 707650 404524
rect 705378 404404 705384 404456
rect 705436 404444 705442 404456
rect 707494 404444 707500 404456
rect 705436 404416 707500 404444
rect 705436 404404 705442 404416
rect 707494 404404 707500 404416
rect 707552 404404 707558 404456
rect 705286 404336 705292 404388
rect 705344 404376 705350 404388
rect 707604 404376 707632 404472
rect 705344 404348 707632 404376
rect 705344 404336 705350 404348
rect 708506 404336 708512 404388
rect 708564 404336 708570 404388
rect 704458 404268 704464 404320
rect 704516 404308 704522 404320
rect 708414 404308 708420 404320
rect 704516 404280 708420 404308
rect 704516 404268 704522 404280
rect 708414 404268 708420 404280
rect 708472 404268 708478 404320
rect 704366 404200 704372 404252
rect 704424 404240 704430 404252
rect 708524 404240 708552 404336
rect 704424 404212 708552 404240
rect 704424 404200 704430 404212
rect 654870 403996 654876 404048
rect 654928 404036 654934 404048
rect 661126 404036 661132 404048
rect 654928 404008 661132 404036
rect 654928 403996 654934 404008
rect 661126 403996 661132 404008
rect 661184 403996 661190 404048
rect 42150 403860 42156 403912
rect 42208 403900 42214 403912
rect 43990 403900 43996 403912
rect 42208 403872 43996 403900
rect 42208 403860 42214 403872
rect 43990 403860 43996 403872
rect 44048 403860 44054 403912
rect 669130 403384 669136 403436
rect 669188 403424 669194 403436
rect 675938 403424 675944 403436
rect 669188 403396 675944 403424
rect 669188 403384 669194 403396
rect 675938 403384 675944 403396
rect 675996 403384 676002 403436
rect 42150 403316 42156 403368
rect 42208 403356 42214 403368
rect 43622 403356 43628 403368
rect 42208 403328 43628 403356
rect 42208 403316 42214 403328
rect 43622 403316 43628 403328
rect 43680 403316 43686 403368
rect 667106 403248 667112 403300
rect 667164 403288 667170 403300
rect 676214 403288 676220 403300
rect 667164 403260 676220 403288
rect 667164 403248 667170 403260
rect 676214 403248 676220 403260
rect 676272 403248 676278 403300
rect 661218 403112 661224 403164
rect 661276 403152 661282 403164
rect 675938 403152 675944 403164
rect 661276 403124 675944 403152
rect 661276 403112 661282 403124
rect 675938 403112 675944 403124
rect 675996 403112 676002 403164
rect 42150 402500 42156 402552
rect 42208 402540 42214 402552
rect 43806 402540 43812 402552
rect 42208 402512 43812 402540
rect 42208 402500 42214 402512
rect 43806 402500 43812 402512
rect 43864 402500 43870 402552
rect 42150 402024 42156 402076
rect 42208 402064 42214 402076
rect 43162 402064 43168 402076
rect 42208 402036 43168 402064
rect 42208 402024 42214 402036
rect 43162 402024 43168 402036
rect 43220 402024 43226 402076
rect 674650 401208 674656 401260
rect 674708 401248 674714 401260
rect 676122 401248 676128 401260
rect 674708 401220 676128 401248
rect 674708 401208 674714 401220
rect 676122 401208 676128 401220
rect 676180 401208 676186 401260
rect 49050 400188 49056 400240
rect 49108 400228 49114 400240
rect 58434 400228 58440 400240
rect 49108 400200 58440 400228
rect 49108 400188 49114 400200
rect 58434 400188 58440 400200
rect 58492 400188 58498 400240
rect 42150 399984 42156 400036
rect 42208 400024 42214 400036
rect 43254 400024 43260 400036
rect 42208 399996 43260 400024
rect 42208 399984 42214 399996
rect 43254 399984 43260 399996
rect 43312 399984 43318 400036
rect 42150 399440 42156 399492
rect 42208 399480 42214 399492
rect 43806 399480 43812 399492
rect 42208 399452 43812 399480
rect 42208 399440 42214 399452
rect 43806 399440 43812 399452
rect 43864 399440 43870 399492
rect 674374 399440 674380 399492
rect 674432 399480 674438 399492
rect 676030 399480 676036 399492
rect 674432 399452 676036 399480
rect 674432 399440 674438 399452
rect 676030 399440 676036 399452
rect 676088 399440 676094 399492
rect 42150 398964 42156 399016
rect 42208 399004 42214 399016
rect 42886 399004 42892 399016
rect 42208 398976 42892 399004
rect 42208 398964 42214 398976
rect 42886 398964 42892 398976
rect 42944 398964 42950 399016
rect 674466 398216 674472 398268
rect 674524 398256 674530 398268
rect 676030 398256 676036 398268
rect 674524 398228 676036 398256
rect 674524 398216 674530 398228
rect 676030 398216 676036 398228
rect 676088 398216 676094 398268
rect 673730 397604 673736 397656
rect 673788 397644 673794 397656
rect 675938 397644 675944 397656
rect 673788 397616 675944 397644
rect 673788 397604 673794 397616
rect 675938 397604 675944 397616
rect 675996 397604 676002 397656
rect 674282 397536 674288 397588
rect 674340 397576 674346 397588
rect 676122 397576 676128 397588
rect 674340 397548 676128 397576
rect 674340 397536 674346 397548
rect 676122 397536 676128 397548
rect 676180 397536 676186 397588
rect 674926 397468 674932 397520
rect 674984 397508 674990 397520
rect 676030 397508 676036 397520
rect 674984 397480 676036 397508
rect 674984 397468 674990 397480
rect 676030 397468 676036 397480
rect 676088 397468 676094 397520
rect 673454 396584 673460 396636
rect 673512 396624 673518 396636
rect 676030 396624 676036 396636
rect 673512 396596 676036 396624
rect 673512 396584 673518 396596
rect 676030 396584 676036 396596
rect 676088 396584 676094 396636
rect 673546 395360 673552 395412
rect 673604 395400 673610 395412
rect 675938 395400 675944 395412
rect 673604 395372 675944 395400
rect 673604 395360 673610 395372
rect 675938 395360 675944 395372
rect 675996 395360 676002 395412
rect 675110 394952 675116 395004
rect 675168 394992 675174 395004
rect 676030 394992 676036 395004
rect 675168 394964 676036 394992
rect 675168 394952 675174 394964
rect 676030 394952 676036 394964
rect 676088 394952 676094 395004
rect 673638 394816 673644 394868
rect 673696 394856 673702 394868
rect 675938 394856 675944 394868
rect 673696 394828 675944 394856
rect 673696 394816 673702 394828
rect 675938 394816 675944 394828
rect 675996 394816 676002 394868
rect 675018 394748 675024 394800
rect 675076 394788 675082 394800
rect 676122 394788 676128 394800
rect 675076 394760 676128 394788
rect 675076 394748 675082 394760
rect 676122 394748 676128 394760
rect 676180 394748 676186 394800
rect 675202 394680 675208 394732
rect 675260 394720 675266 394732
rect 676030 394720 676036 394732
rect 675260 394692 676036 394720
rect 675260 394680 675266 394692
rect 676030 394680 676036 394692
rect 676088 394680 676094 394732
rect 673822 394136 673828 394188
rect 673880 394176 673886 394188
rect 676030 394176 676036 394188
rect 673880 394148 676036 394176
rect 673880 394136 673886 394148
rect 676030 394136 676036 394148
rect 676088 394136 676094 394188
rect 672902 392028 672908 392080
rect 672960 392068 672966 392080
rect 678974 392068 678980 392080
rect 672960 392040 678980 392068
rect 672960 392028 672966 392040
rect 678974 392028 678980 392040
rect 679032 392028 679038 392080
rect 674006 391960 674012 392012
rect 674064 392000 674070 392012
rect 676030 392000 676036 392012
rect 674064 391972 676036 392000
rect 674064 391960 674070 391972
rect 676030 391960 676036 391972
rect 676088 391960 676094 392012
rect 674742 390532 674748 390584
rect 674800 390572 674806 390584
rect 675754 390572 675760 390584
rect 674800 390544 675760 390572
rect 674800 390532 674806 390544
rect 675754 390532 675760 390544
rect 675812 390532 675818 390584
rect 674558 390464 674564 390516
rect 674616 390504 674622 390516
rect 675662 390504 675668 390516
rect 674616 390476 675668 390504
rect 674616 390464 674622 390476
rect 675662 390464 675668 390476
rect 675720 390464 675726 390516
rect 654134 389784 654140 389836
rect 654192 389824 654198 389836
rect 669590 389824 669596 389836
rect 654192 389796 669596 389824
rect 654192 389784 654198 389796
rect 669590 389784 669596 389796
rect 669648 389784 669654 389836
rect 53834 389172 53840 389224
rect 53892 389212 53898 389224
rect 57974 389212 57980 389224
rect 53892 389184 57980 389212
rect 53892 389172 53898 389184
rect 57974 389172 57980 389184
rect 58032 389172 58038 389224
rect 41506 387948 41512 388000
rect 41564 387988 41570 388000
rect 51166 387988 51172 388000
rect 41564 387960 51172 387988
rect 41564 387948 41570 387960
rect 51166 387948 51172 387960
rect 51224 387948 51230 388000
rect 41782 387404 41788 387456
rect 41840 387444 41846 387456
rect 54018 387444 54024 387456
rect 41840 387416 54024 387444
rect 41840 387404 41846 387416
rect 54018 387404 54024 387416
rect 54076 387404 54082 387456
rect 41506 387132 41512 387184
rect 41564 387172 41570 387184
rect 49142 387172 49148 387184
rect 41564 387144 49148 387172
rect 41564 387132 41570 387144
rect 49142 387132 49148 387144
rect 49200 387132 49206 387184
rect 42794 386384 42800 386436
rect 42852 386424 42858 386436
rect 63126 386424 63132 386436
rect 42852 386396 63132 386424
rect 42852 386384 42858 386396
rect 63126 386384 63132 386396
rect 63184 386384 63190 386436
rect 675754 386384 675760 386436
rect 675812 386384 675818 386436
rect 675772 386164 675800 386384
rect 675754 386112 675760 386164
rect 675812 386112 675818 386164
rect 674466 384956 674472 385008
rect 674524 384996 674530 385008
rect 675294 384996 675300 385008
rect 674524 384968 675300 384996
rect 674524 384956 674530 384968
rect 675294 384956 675300 384968
rect 675352 384956 675358 385008
rect 675202 384072 675208 384124
rect 675260 384072 675266 384124
rect 675220 383908 675248 384072
rect 675294 383908 675300 383920
rect 675220 383880 675300 383908
rect 675294 383868 675300 383880
rect 675352 383868 675358 383920
rect 674926 383120 674932 383172
rect 674984 383160 674990 383172
rect 675386 383160 675392 383172
rect 674984 383132 675392 383160
rect 674984 383120 674990 383132
rect 675386 383120 675392 383132
rect 675444 383120 675450 383172
rect 675110 382440 675116 382492
rect 675168 382480 675174 382492
rect 675386 382480 675392 382492
rect 675168 382452 675392 382480
rect 675168 382440 675174 382452
rect 675386 382440 675392 382452
rect 675444 382440 675450 382492
rect 674374 382304 674380 382356
rect 674432 382344 674438 382356
rect 675110 382344 675116 382356
rect 674432 382316 675116 382344
rect 674432 382304 674438 382316
rect 675110 382304 675116 382316
rect 675168 382304 675174 382356
rect 675018 381896 675024 381948
rect 675076 381936 675082 381948
rect 675386 381936 675392 381948
rect 675076 381908 675392 381936
rect 675076 381896 675082 381908
rect 675386 381896 675392 381908
rect 675444 381896 675450 381948
rect 673730 379448 673736 379500
rect 673788 379488 673794 379500
rect 675294 379488 675300 379500
rect 673788 379460 675300 379488
rect 673788 379448 673794 379460
rect 675294 379448 675300 379460
rect 675352 379448 675358 379500
rect 656802 378156 656808 378208
rect 656860 378196 656866 378208
rect 669682 378196 669688 378208
rect 656860 378168 669688 378196
rect 656860 378156 656866 378168
rect 669682 378156 669688 378168
rect 669740 378156 669746 378208
rect 673638 378156 673644 378208
rect 673696 378196 673702 378208
rect 675294 378196 675300 378208
rect 673696 378168 675300 378196
rect 673696 378156 673702 378168
rect 675294 378156 675300 378168
rect 675352 378156 675358 378208
rect 673822 377952 673828 378004
rect 673880 377992 673886 378004
rect 675478 377992 675484 378004
rect 673880 377964 675484 377992
rect 673880 377952 673886 377964
rect 675478 377952 675484 377964
rect 675536 377952 675542 378004
rect 674006 376932 674012 376984
rect 674064 376972 674070 376984
rect 675478 376972 675484 376984
rect 674064 376944 675484 376972
rect 674064 376932 674070 376944
rect 675478 376932 675484 376944
rect 675536 376932 675542 376984
rect 673546 376864 673552 376916
rect 673604 376904 673610 376916
rect 675294 376904 675300 376916
rect 673604 376876 675300 376904
rect 673604 376864 673610 376876
rect 675294 376864 675300 376876
rect 675352 376864 675358 376916
rect 41414 376456 41420 376508
rect 41472 376496 41478 376508
rect 46750 376496 46756 376508
rect 41472 376468 46756 376496
rect 41472 376456 41478 376468
rect 46750 376456 46756 376468
rect 46808 376456 46814 376508
rect 49142 375368 49148 375420
rect 49200 375408 49206 375420
rect 58434 375408 58440 375420
rect 49200 375380 58440 375408
rect 49200 375368 49206 375380
rect 58434 375368 58440 375380
rect 58492 375368 58498 375420
rect 675110 374076 675116 374128
rect 675168 374116 675174 374128
rect 675294 374116 675300 374128
rect 675168 374088 675300 374116
rect 675168 374076 675174 374088
rect 675294 374076 675300 374088
rect 675352 374076 675358 374128
rect 674282 373872 674288 373924
rect 674340 373912 674346 373924
rect 675386 373912 675392 373924
rect 674340 373884 675392 373912
rect 674340 373872 674346 373884
rect 675386 373872 675392 373884
rect 675444 373872 675450 373924
rect 675294 372852 675300 372904
rect 675352 372852 675358 372904
rect 675312 372700 675340 372852
rect 675294 372648 675300 372700
rect 675352 372648 675358 372700
rect 673454 372036 673460 372088
rect 673512 372076 673518 372088
rect 675386 372076 675392 372088
rect 673512 372048 675392 372076
rect 673512 372036 673518 372048
rect 675386 372036 675392 372048
rect 675444 372036 675450 372088
rect 42794 371764 42800 371816
rect 42852 371804 42858 371816
rect 43346 371804 43352 371816
rect 42852 371776 43352 371804
rect 42852 371764 42858 371776
rect 43346 371764 43352 371776
rect 43404 371764 43410 371816
rect 41506 371424 41512 371476
rect 41564 371464 41570 371476
rect 42794 371464 42800 371476
rect 41564 371436 42800 371464
rect 41564 371424 41570 371436
rect 42794 371424 42800 371436
rect 42852 371424 42858 371476
rect 674742 370744 674748 370796
rect 674800 370784 674806 370796
rect 675754 370784 675760 370796
rect 674800 370756 675760 370784
rect 674800 370744 674806 370756
rect 675754 370744 675760 370756
rect 675812 370744 675818 370796
rect 674558 370676 674564 370728
rect 674616 370716 674622 370728
rect 675662 370716 675668 370728
rect 674616 370688 675668 370716
rect 674616 370676 674622 370688
rect 675662 370676 675668 370688
rect 675720 370676 675726 370728
rect 42150 369928 42156 369980
rect 42208 369968 42214 369980
rect 42334 369968 42340 369980
rect 42208 369940 42340 369968
rect 42208 369928 42214 369940
rect 42334 369928 42340 369940
rect 42392 369928 42398 369980
rect 42150 368092 42156 368144
rect 42208 368132 42214 368144
rect 42702 368132 42708 368144
rect 42208 368104 42708 368132
rect 42208 368092 42214 368104
rect 42702 368092 42708 368104
rect 42760 368092 42766 368144
rect 42150 366800 42156 366852
rect 42208 366840 42214 366852
rect 50982 366840 50988 366852
rect 42208 366812 50988 366840
rect 42208 366800 42214 366812
rect 50982 366800 50988 366812
rect 51040 366800 51046 366852
rect 42150 366256 42156 366308
rect 42208 366296 42214 366308
rect 43070 366296 43076 366308
rect 42208 366268 43076 366296
rect 42208 366256 42214 366268
rect 43070 366256 43076 366268
rect 43128 366256 43134 366308
rect 42150 364964 42156 365016
rect 42208 365004 42214 365016
rect 42794 365004 42800 365016
rect 42208 364976 42800 365004
rect 42208 364964 42214 364976
rect 42794 364964 42800 364976
rect 42852 364964 42858 365016
rect 42150 364420 42156 364472
rect 42208 364460 42214 364472
rect 43254 364460 43260 364472
rect 42208 364432 43260 364460
rect 42208 364420 42214 364432
rect 43254 364420 43260 364432
rect 43312 364420 43318 364472
rect 656802 364352 656808 364404
rect 656860 364392 656866 364404
rect 667106 364392 667112 364404
rect 656860 364364 667112 364392
rect 656860 364352 656866 364364
rect 667106 364352 667112 364364
rect 667164 364352 667170 364404
rect 42150 363808 42156 363860
rect 42208 363848 42214 363860
rect 43162 363848 43168 363860
rect 42208 363820 43168 363848
rect 42208 363808 42214 363820
rect 43162 363808 43168 363820
rect 43220 363808 43226 363860
rect 42150 363128 42156 363180
rect 42208 363168 42214 363180
rect 43346 363168 43352 363180
rect 42208 363140 43352 363168
rect 42208 363128 42214 363140
rect 43346 363128 43352 363140
rect 43404 363128 43410 363180
rect 43162 362788 43168 362840
rect 43220 362828 43226 362840
rect 43622 362828 43628 362840
rect 43220 362800 43628 362828
rect 43220 362788 43226 362800
rect 43622 362788 43628 362800
rect 43680 362788 43686 362840
rect 703446 361700 703452 361752
rect 703504 361740 703510 361752
rect 709334 361740 709340 361752
rect 703504 361712 709340 361740
rect 703504 361700 703510 361712
rect 709334 361700 709340 361712
rect 709392 361700 709398 361752
rect 51166 361564 51172 361616
rect 51224 361604 51230 361616
rect 58434 361604 58440 361616
rect 51224 361576 58440 361604
rect 51224 361564 51230 361576
rect 58434 361564 58440 361576
rect 58492 361564 58498 361616
rect 42058 360680 42064 360732
rect 42116 360720 42122 360732
rect 43070 360720 43076 360732
rect 42116 360692 43076 360720
rect 42116 360680 42122 360692
rect 43070 360680 43076 360692
rect 43128 360680 43134 360732
rect 42150 359932 42156 359984
rect 42208 359972 42214 359984
rect 43806 359972 43812 359984
rect 42208 359944 43812 359972
rect 42208 359932 42214 359944
rect 43806 359932 43812 359944
rect 43864 359932 43870 359984
rect 708506 359700 708512 359712
rect 704384 359672 708512 359700
rect 704384 359576 704412 359672
rect 708506 359660 708512 359672
rect 708564 359660 708570 359712
rect 704458 359592 704464 359644
rect 704516 359632 704522 359644
rect 708414 359632 708420 359644
rect 704516 359604 708420 359632
rect 704516 359592 704522 359604
rect 708414 359592 708420 359604
rect 708472 359592 708478 359644
rect 704366 359524 704372 359576
rect 704424 359524 704430 359576
rect 707494 359564 707500 359576
rect 705304 359536 707500 359564
rect 42150 359456 42156 359508
rect 42208 359496 42214 359508
rect 43622 359496 43628 359508
rect 42208 359468 43628 359496
rect 42208 359456 42214 359468
rect 43622 359456 43628 359468
rect 43680 359456 43686 359508
rect 705304 359440 705332 359536
rect 707494 359524 707500 359536
rect 707552 359524 707558 359576
rect 707034 359496 707040 359508
rect 705764 359468 707040 359496
rect 705764 359440 705792 359468
rect 707034 359456 707040 359468
rect 707092 359456 707098 359508
rect 705286 359388 705292 359440
rect 705344 359388 705350 359440
rect 705746 359388 705752 359440
rect 705804 359388 705810 359440
rect 706206 359388 706212 359440
rect 706264 359428 706270 359440
rect 706574 359428 706580 359440
rect 706264 359400 706580 359428
rect 706264 359388 706270 359400
rect 706574 359388 706580 359400
rect 706632 359388 706638 359440
rect 705838 359320 705844 359372
rect 705896 359360 705902 359372
rect 707034 359360 707040 359372
rect 705896 359332 707040 359360
rect 705896 359320 705902 359332
rect 707034 359320 707040 359332
rect 707092 359320 707098 359372
rect 706298 359252 706304 359304
rect 706356 359292 706362 359304
rect 706574 359292 706580 359304
rect 706356 359264 706580 359292
rect 706356 359252 706362 359264
rect 706574 359252 706580 359264
rect 706632 359252 706638 359304
rect 705378 359184 705384 359236
rect 705436 359224 705442 359236
rect 707494 359224 707500 359236
rect 705436 359196 707500 359224
rect 705436 359184 705442 359196
rect 707494 359184 707500 359196
rect 707552 359184 707558 359236
rect 708046 359184 708052 359236
rect 708104 359184 708110 359236
rect 704918 359116 704924 359168
rect 704976 359156 704982 359168
rect 707954 359156 707960 359168
rect 704976 359128 707960 359156
rect 704976 359116 704982 359128
rect 707954 359116 707960 359128
rect 708012 359116 708018 359168
rect 704826 359048 704832 359100
rect 704884 359088 704890 359100
rect 708064 359088 708092 359184
rect 704884 359060 708092 359088
rect 704884 359048 704890 359060
rect 703814 358844 703820 358896
rect 703872 358844 703878 358896
rect 708874 358844 708880 358896
rect 708932 358844 708938 358896
rect 42058 358776 42064 358828
rect 42116 358816 42122 358828
rect 42886 358816 42892 358828
rect 42116 358788 42892 358816
rect 42116 358776 42122 358788
rect 42886 358776 42892 358788
rect 42944 358776 42950 358828
rect 703832 358748 703860 358844
rect 708892 358748 708920 358844
rect 703832 358720 708920 358748
rect 673270 357008 673276 357060
rect 673328 357048 673334 357060
rect 675570 357048 675576 357060
rect 673328 357020 675576 357048
rect 673328 357008 673334 357020
rect 675570 357008 675576 357020
rect 675628 357008 675634 357060
rect 42058 356940 42064 356992
rect 42116 356980 42122 356992
rect 42978 356980 42984 356992
rect 42116 356952 42984 356980
rect 42116 356940 42122 356952
rect 42978 356940 42984 356952
rect 43036 356940 43042 356992
rect 670050 356464 670056 356516
rect 670108 356504 670114 356516
rect 676030 356504 676036 356516
rect 670108 356476 676036 356504
rect 670108 356464 670114 356476
rect 676030 356464 676036 356476
rect 676088 356464 676094 356516
rect 667014 356328 667020 356380
rect 667072 356368 667078 356380
rect 675938 356368 675944 356380
rect 667072 356340 675944 356368
rect 667072 356328 667078 356340
rect 675938 356328 675944 356340
rect 675996 356328 676002 356380
rect 42150 356260 42156 356312
rect 42208 356300 42214 356312
rect 43162 356300 43168 356312
rect 42208 356272 43168 356300
rect 42208 356260 42214 356272
rect 43162 356260 43168 356272
rect 43220 356260 43226 356312
rect 663794 356192 663800 356244
rect 663852 356232 663858 356244
rect 675846 356232 675852 356244
rect 663852 356204 675852 356232
rect 663852 356192 663858 356204
rect 675846 356192 675852 356204
rect 675904 356192 675910 356244
rect 673362 356124 673368 356176
rect 673420 356164 673426 356176
rect 676030 356164 676036 356176
rect 673420 356136 676036 356164
rect 673420 356124 673426 356136
rect 676030 356124 676036 356136
rect 676088 356124 676094 356176
rect 669498 356056 669504 356108
rect 669556 356096 669562 356108
rect 672994 356096 673000 356108
rect 669556 356068 673000 356096
rect 669556 356056 669562 356068
rect 672994 356056 673000 356068
rect 673052 356096 673058 356108
rect 673270 356096 673276 356108
rect 673052 356068 673276 356096
rect 673052 356056 673058 356068
rect 673270 356056 673276 356068
rect 673328 356056 673334 356108
rect 673178 355376 673184 355428
rect 673236 355416 673242 355428
rect 676030 355416 676036 355428
rect 673236 355388 676036 355416
rect 673236 355376 673242 355388
rect 676030 355376 676036 355388
rect 676088 355376 676094 355428
rect 673270 354560 673276 354612
rect 673328 354600 673334 354612
rect 676030 354600 676036 354612
rect 673328 354572 676036 354600
rect 673328 354560 673334 354572
rect 676030 354560 676036 354572
rect 676088 354560 676094 354612
rect 669406 353472 669412 353524
rect 669464 353512 669470 353524
rect 673086 353512 673092 353524
rect 669464 353484 673092 353512
rect 669464 353472 669470 353484
rect 673086 353472 673092 353484
rect 673144 353512 673150 353524
rect 673270 353512 673276 353524
rect 673144 353484 673276 353512
rect 673144 353472 673150 353484
rect 673270 353472 673276 353484
rect 673328 353472 673334 353524
rect 673546 353472 673552 353524
rect 673604 353512 673610 353524
rect 676030 353512 676036 353524
rect 673604 353484 676036 353512
rect 673604 353472 673610 353484
rect 676030 353472 676036 353484
rect 676088 353472 676094 353524
rect 669314 353336 669320 353388
rect 669372 353376 669378 353388
rect 673178 353376 673184 353388
rect 669372 353348 673184 353376
rect 669372 353336 669378 353348
rect 673178 353336 673184 353348
rect 673236 353336 673242 353388
rect 674006 353268 674012 353320
rect 674064 353308 674070 353320
rect 676030 353308 676036 353320
rect 674064 353280 676036 353308
rect 674064 353268 674070 353280
rect 676030 353268 676036 353280
rect 676088 353268 676094 353320
rect 674558 351432 674564 351484
rect 674616 351472 674622 351484
rect 676030 351472 676036 351484
rect 674616 351444 676036 351472
rect 674616 351432 674622 351444
rect 676030 351432 676036 351444
rect 676088 351432 676094 351484
rect 673454 351024 673460 351076
rect 673512 351064 673518 351076
rect 675938 351064 675944 351076
rect 673512 351036 675944 351064
rect 673512 351024 673518 351036
rect 675938 351024 675944 351036
rect 675996 351024 676002 351076
rect 674650 350616 674656 350668
rect 674708 350656 674714 350668
rect 675938 350656 675944 350668
rect 674708 350628 675944 350656
rect 674708 350616 674714 350628
rect 675938 350616 675944 350628
rect 675996 350616 676002 350668
rect 654870 350548 654876 350600
rect 654928 350588 654934 350600
rect 669406 350588 669412 350600
rect 654928 350560 669412 350588
rect 654928 350548 654934 350560
rect 669406 350548 669412 350560
rect 669464 350548 669470 350600
rect 674742 350548 674748 350600
rect 674800 350588 674806 350600
rect 676030 350588 676036 350600
rect 674800 350560 676036 350588
rect 674800 350548 674806 350560
rect 676030 350548 676036 350560
rect 676088 350548 676094 350600
rect 673730 349800 673736 349852
rect 673788 349840 673794 349852
rect 676030 349840 676036 349852
rect 673788 349812 676036 349840
rect 673788 349800 673794 349812
rect 676030 349800 676036 349812
rect 676088 349800 676094 349852
rect 673822 347896 673828 347948
rect 673880 347936 673886 347948
rect 675846 347936 675852 347948
rect 673880 347908 675852 347936
rect 673880 347896 673886 347908
rect 675846 347896 675852 347908
rect 675904 347896 675910 347948
rect 673914 347828 673920 347880
rect 673972 347868 673978 347880
rect 675938 347868 675944 347880
rect 673972 347840 675944 347868
rect 673972 347828 673978 347840
rect 675938 347828 675944 347840
rect 675996 347828 676002 347880
rect 50982 347760 50988 347812
rect 51040 347800 51046 347812
rect 58434 347800 58440 347812
rect 51040 347772 58440 347800
rect 51040 347760 51046 347772
rect 58434 347760 58440 347772
rect 58492 347760 58498 347812
rect 674834 347760 674840 347812
rect 674892 347800 674898 347812
rect 676030 347800 676036 347812
rect 674892 347772 676036 347800
rect 674892 347760 674898 347772
rect 676030 347760 676036 347772
rect 676088 347760 676094 347812
rect 44358 344972 44364 345024
rect 44416 345012 44422 345024
rect 48406 345012 48412 345024
rect 44416 344984 48412 345012
rect 44416 344972 44422 344984
rect 48406 344972 48412 344984
rect 48464 344972 48470 345024
rect 41506 344224 41512 344276
rect 41564 344264 41570 344276
rect 53926 344264 53932 344276
rect 41564 344236 53932 344264
rect 41564 344224 41570 344236
rect 53926 344224 53932 344236
rect 53984 344224 53990 344276
rect 41782 344156 41788 344208
rect 41840 344196 41846 344208
rect 49234 344196 49240 344208
rect 41840 344168 49240 344196
rect 41840 344156 41846 344168
rect 49234 344156 49240 344168
rect 49292 344156 49298 344208
rect 41506 344088 41512 344140
rect 41564 344128 41570 344140
rect 43530 344128 43536 344140
rect 41564 344100 43536 344128
rect 41564 344088 41570 344100
rect 43530 344088 43536 344100
rect 43588 344088 43594 344140
rect 41598 343884 41604 343936
rect 41656 343924 41662 343936
rect 51074 343924 51080 343936
rect 41656 343896 51080 343924
rect 41656 343884 41662 343896
rect 51074 343884 51080 343896
rect 51132 343884 51138 343936
rect 41782 343340 41788 343392
rect 41840 343380 41846 343392
rect 44358 343380 44364 343392
rect 41840 343352 44364 343380
rect 41840 343340 41846 343352
rect 44358 343340 44364 343352
rect 44416 343340 44422 343392
rect 672994 342388 673000 342440
rect 673052 342428 673058 342440
rect 675754 342428 675760 342440
rect 673052 342400 675760 342428
rect 673052 342388 673058 342400
rect 675754 342388 675760 342400
rect 675812 342388 675818 342440
rect 674006 340960 674012 341012
rect 674064 341000 674070 341012
rect 675478 341000 675484 341012
rect 674064 340972 675484 341000
rect 674064 340960 674070 340972
rect 675478 340960 675484 340972
rect 675536 340960 675542 341012
rect 673546 339736 673552 339788
rect 673604 339776 673610 339788
rect 675478 339776 675484 339788
rect 673604 339748 675484 339776
rect 673604 339736 673610 339748
rect 675478 339736 675484 339748
rect 675536 339736 675542 339788
rect 674558 337900 674564 337952
rect 674616 337940 674622 337952
rect 675478 337940 675484 337952
rect 674616 337912 675484 337940
rect 674616 337900 674622 337912
rect 675478 337900 675484 337912
rect 675536 337900 675542 337952
rect 674742 337016 674748 337068
rect 674800 337056 674806 337068
rect 675386 337056 675392 337068
rect 674800 337028 675392 337056
rect 674800 337016 674806 337028
rect 675386 337016 675392 337028
rect 675444 337016 675450 337068
rect 654318 336812 654324 336864
rect 654376 336852 654382 336864
rect 667014 336852 667020 336864
rect 654376 336824 667020 336852
rect 654376 336812 654382 336824
rect 667014 336812 667020 336824
rect 667072 336812 667078 336864
rect 48406 336744 48412 336796
rect 48464 336784 48470 336796
rect 58434 336784 58440 336796
rect 48464 336756 58440 336784
rect 48464 336744 48470 336756
rect 58434 336744 58440 336756
rect 58492 336744 58498 336796
rect 674650 336540 674656 336592
rect 674708 336580 674714 336592
rect 675386 336580 675392 336592
rect 674708 336552 675392 336580
rect 674708 336540 674714 336552
rect 675386 336540 675392 336552
rect 675444 336540 675450 336592
rect 674834 336064 674840 336116
rect 674892 336104 674898 336116
rect 675478 336104 675484 336116
rect 674892 336076 675484 336104
rect 674892 336064 674898 336076
rect 675478 336064 675484 336076
rect 675536 336064 675542 336116
rect 673454 333548 673460 333600
rect 673512 333588 673518 333600
rect 675386 333588 675392 333600
rect 673512 333560 675392 333588
rect 673512 333548 673518 333560
rect 675386 333548 675392 333560
rect 675444 333548 675450 333600
rect 41506 333208 41512 333260
rect 41564 333248 41570 333260
rect 46198 333248 46204 333260
rect 41564 333220 46204 333248
rect 41564 333208 41570 333220
rect 46198 333208 46204 333220
rect 46256 333208 46262 333260
rect 673914 332936 673920 332988
rect 673972 332976 673978 332988
rect 675386 332976 675392 332988
rect 673972 332948 675392 332976
rect 673972 332936 673978 332948
rect 675386 332936 675392 332948
rect 675444 332936 675450 332988
rect 673730 332188 673736 332240
rect 673788 332228 673794 332240
rect 675386 332228 675392 332240
rect 673788 332200 675392 332228
rect 673788 332188 673794 332200
rect 675386 332188 675392 332200
rect 675444 332188 675450 332240
rect 673822 331576 673828 331628
rect 673880 331616 673886 331628
rect 675386 331616 675392 331628
rect 673880 331588 675392 331616
rect 673880 331576 673886 331588
rect 675386 331576 675392 331588
rect 675444 331576 675450 331628
rect 33042 330080 33048 330132
rect 33100 330120 33106 330132
rect 41874 330120 41880 330132
rect 33100 330092 41880 330120
rect 33100 330080 33106 330092
rect 41874 330080 41880 330092
rect 41932 330080 41938 330132
rect 32950 329944 32956 329996
rect 33008 329984 33014 329996
rect 42886 329984 42892 329996
rect 33008 329956 42892 329984
rect 33008 329944 33014 329956
rect 42886 329944 42892 329956
rect 42944 329944 42950 329996
rect 32674 329876 32680 329928
rect 32732 329916 32738 329928
rect 42794 329916 42800 329928
rect 32732 329888 42800 329916
rect 32732 329876 32738 329888
rect 42794 329876 42800 329888
rect 42852 329876 42858 329928
rect 32858 329808 32864 329860
rect 32916 329848 32922 329860
rect 43346 329848 43352 329860
rect 32916 329820 43352 329848
rect 32916 329808 32922 329820
rect 43346 329808 43352 329820
rect 43404 329808 43410 329860
rect 41874 326952 41880 327004
rect 41932 326952 41938 327004
rect 41892 326800 41920 326952
rect 41874 326748 41880 326800
rect 41932 326748 41938 326800
rect 42058 324912 42064 324964
rect 42116 324952 42122 324964
rect 42794 324952 42800 324964
rect 42116 324924 42800 324952
rect 42116 324912 42122 324924
rect 42794 324912 42800 324924
rect 42852 324912 42858 324964
rect 42794 324776 42800 324828
rect 42852 324816 42858 324828
rect 43070 324816 43076 324828
rect 42852 324788 43076 324816
rect 42852 324776 42858 324788
rect 43070 324776 43076 324788
rect 43128 324776 43134 324828
rect 654318 323892 654324 323944
rect 654376 323932 654382 323944
rect 669130 323932 669136 323944
rect 654376 323904 669136 323932
rect 654376 323892 654382 323904
rect 669130 323892 669136 323904
rect 669188 323892 669194 323944
rect 53926 323484 53932 323536
rect 53984 323524 53990 323536
rect 58158 323524 58164 323536
rect 53984 323496 58164 323524
rect 53984 323484 53990 323496
rect 58158 323484 58164 323496
rect 58216 323484 58222 323536
rect 42150 323280 42156 323332
rect 42208 323320 42214 323332
rect 42610 323320 42616 323332
rect 42208 323292 42616 323320
rect 42208 323280 42214 323292
rect 42610 323280 42616 323292
rect 42668 323280 42674 323332
rect 42058 323076 42064 323128
rect 42116 323116 42122 323128
rect 42886 323116 42892 323128
rect 42116 323088 42892 323116
rect 42116 323076 42122 323088
rect 42886 323076 42892 323088
rect 42944 323076 42950 323128
rect 42150 321784 42156 321836
rect 42208 321824 42214 321836
rect 43162 321824 43168 321836
rect 42208 321796 43168 321824
rect 42208 321784 42214 321796
rect 43162 321784 43168 321796
rect 43220 321784 43226 321836
rect 42150 321036 42156 321088
rect 42208 321076 42214 321088
rect 43346 321076 43352 321088
rect 42208 321048 43352 321076
rect 42208 321036 42214 321048
rect 43346 321036 43352 321048
rect 43404 321036 43410 321088
rect 42150 320560 42156 320612
rect 42208 320600 42214 320612
rect 42978 320600 42984 320612
rect 42208 320572 42984 320600
rect 42208 320560 42214 320572
rect 42978 320560 42984 320572
rect 43036 320560 43042 320612
rect 42610 320084 42616 320136
rect 42668 320124 42674 320136
rect 53742 320124 53748 320136
rect 42668 320096 53748 320124
rect 42668 320084 42674 320096
rect 53742 320084 53748 320096
rect 53800 320084 53806 320136
rect 42150 317432 42156 317484
rect 42208 317472 42214 317484
rect 42794 317472 42800 317484
rect 42208 317444 42800 317472
rect 42208 317432 42214 317444
rect 42794 317432 42800 317444
rect 42852 317432 42858 317484
rect 703998 314712 704004 314764
rect 704056 314752 704062 314764
rect 708874 314752 708880 314764
rect 704056 314724 708880 314752
rect 704056 314712 704062 314724
rect 708874 314712 708880 314724
rect 708932 314712 708938 314764
rect 708506 314684 708512 314696
rect 704384 314656 708512 314684
rect 658458 314576 658464 314628
rect 658516 314616 658522 314628
rect 671154 314616 671160 314628
rect 658516 314588 671160 314616
rect 658516 314576 658522 314588
rect 671154 314576 671160 314588
rect 671212 314576 671218 314628
rect 704384 314560 704412 314656
rect 708506 314644 708512 314656
rect 708564 314644 708570 314696
rect 704458 314576 704464 314628
rect 704516 314616 704522 314628
rect 708414 314616 708420 314628
rect 704516 314588 708420 314616
rect 704516 314576 704522 314588
rect 708414 314576 708420 314588
rect 708472 314576 708478 314628
rect 704366 314508 704372 314560
rect 704424 314508 704430 314560
rect 707494 314548 707500 314560
rect 705304 314520 707500 314548
rect 705304 314424 705332 314520
rect 707494 314508 707500 314520
rect 707552 314508 707558 314560
rect 707034 314480 707040 314492
rect 705764 314452 707040 314480
rect 705764 314424 705792 314452
rect 707034 314440 707040 314452
rect 707092 314440 707098 314492
rect 705286 314372 705292 314424
rect 705344 314372 705350 314424
rect 705746 314372 705752 314424
rect 705804 314372 705810 314424
rect 706206 314372 706212 314424
rect 706264 314412 706270 314424
rect 706574 314412 706580 314424
rect 706264 314384 706580 314412
rect 706264 314372 706270 314384
rect 706574 314372 706580 314384
rect 706632 314372 706638 314424
rect 705838 314304 705844 314356
rect 705896 314344 705902 314356
rect 707034 314344 707040 314356
rect 705896 314316 707040 314344
rect 705896 314304 705902 314316
rect 707034 314304 707040 314316
rect 707092 314304 707098 314356
rect 706298 314236 706304 314288
rect 706356 314276 706362 314288
rect 706574 314276 706580 314288
rect 706356 314248 706580 314276
rect 706356 314236 706362 314248
rect 706574 314236 706580 314248
rect 706632 314236 706638 314288
rect 705378 314168 705384 314220
rect 705436 314208 705442 314220
rect 707494 314208 707500 314220
rect 705436 314180 707500 314208
rect 705436 314168 705442 314180
rect 707494 314168 707500 314180
rect 707552 314168 707558 314220
rect 708046 314168 708052 314220
rect 708104 314168 708110 314220
rect 704918 314100 704924 314152
rect 704976 314140 704982 314152
rect 707954 314140 707960 314152
rect 704976 314112 707960 314140
rect 704976 314100 704982 314112
rect 707954 314100 707960 314112
rect 708012 314100 708018 314152
rect 704826 314032 704832 314084
rect 704884 314072 704890 314084
rect 708064 314072 708092 314168
rect 704884 314044 708092 314072
rect 704884 314032 704890 314044
rect 703538 313964 703544 314016
rect 703596 314004 703602 314016
rect 708874 314004 708880 314016
rect 703596 313976 708880 314004
rect 703596 313964 703602 313976
rect 708874 313964 708880 313976
rect 708932 313964 708938 314016
rect 663702 313284 663708 313336
rect 663760 313324 663766 313336
rect 676030 313324 676036 313336
rect 663760 313296 676036 313324
rect 663760 313284 663766 313296
rect 676030 313284 676036 313296
rect 676088 313284 676094 313336
rect 663886 312876 663892 312928
rect 663944 312916 663950 312928
rect 676030 312916 676036 312928
rect 663944 312888 676036 312916
rect 663944 312876 663950 312888
rect 676030 312876 676036 312888
rect 676088 312876 676094 312928
rect 673178 312468 673184 312520
rect 673236 312508 673242 312520
rect 676030 312508 676036 312520
rect 673236 312480 676036 312508
rect 673236 312468 673242 312480
rect 676030 312468 676036 312480
rect 676088 312468 676094 312520
rect 671154 312060 671160 312112
rect 671212 312100 671218 312112
rect 672258 312100 672264 312112
rect 671212 312072 672264 312100
rect 671212 312060 671218 312072
rect 672258 312060 672264 312072
rect 672316 312100 672322 312112
rect 676030 312100 676036 312112
rect 672316 312072 676036 312100
rect 672316 312060 672322 312072
rect 676030 312060 676036 312072
rect 676088 312060 676094 312112
rect 661034 311992 661040 312044
rect 661092 312032 661098 312044
rect 676214 312032 676220 312044
rect 661092 312004 676220 312032
rect 661092 311992 661098 312004
rect 676214 311992 676220 312004
rect 676272 311992 676278 312044
rect 658366 311788 658372 311840
rect 658424 311828 658430 311840
rect 671154 311828 671160 311840
rect 658424 311800 671160 311828
rect 658424 311788 658430 311800
rect 671154 311788 671160 311800
rect 671212 311788 671218 311840
rect 654134 311652 654140 311704
rect 654192 311692 654198 311704
rect 669314 311692 669320 311704
rect 654192 311664 669320 311692
rect 654192 311652 654198 311664
rect 669314 311652 669320 311664
rect 669372 311652 669378 311704
rect 673362 311652 673368 311704
rect 673420 311692 673426 311704
rect 676030 311692 676036 311704
rect 673420 311664 676036 311692
rect 673420 311652 673426 311664
rect 676030 311652 676036 311664
rect 676088 311652 676094 311704
rect 674742 310972 674748 311024
rect 674800 311012 674806 311024
rect 676030 311012 676036 311024
rect 674800 310984 676036 311012
rect 674800 310972 674806 310984
rect 676030 310972 676036 310984
rect 676088 310972 676094 311024
rect 673270 310836 673276 310888
rect 673328 310876 673334 310888
rect 676030 310876 676036 310888
rect 673328 310848 676036 310876
rect 673328 310836 673334 310848
rect 676030 310836 676036 310848
rect 676088 310836 676094 310888
rect 655422 310428 655428 310480
rect 655480 310468 655486 310480
rect 671890 310468 671896 310480
rect 655480 310440 671896 310468
rect 655480 310428 655486 310440
rect 671890 310428 671896 310440
rect 671948 310468 671954 310480
rect 676030 310468 676036 310480
rect 671948 310440 676036 310468
rect 671948 310428 671954 310440
rect 676030 310428 676036 310440
rect 676088 310428 676094 310480
rect 673086 310020 673092 310072
rect 673144 310060 673150 310072
rect 676030 310060 676036 310072
rect 673144 310032 676036 310060
rect 673144 310020 673150 310032
rect 676030 310020 676036 310032
rect 676088 310020 676094 310072
rect 671154 309612 671160 309664
rect 671212 309652 671218 309664
rect 673178 309652 673184 309664
rect 671212 309624 673184 309652
rect 671212 309612 671218 309624
rect 673178 309612 673184 309624
rect 673236 309652 673242 309664
rect 676030 309652 676036 309664
rect 673236 309624 676036 309652
rect 673236 309612 673242 309624
rect 676030 309612 676036 309624
rect 676088 309612 676094 309664
rect 674190 309136 674196 309188
rect 674248 309176 674254 309188
rect 676030 309176 676036 309188
rect 674248 309148 676036 309176
rect 674248 309136 674254 309148
rect 676030 309136 676036 309148
rect 676088 309136 676094 309188
rect 673546 308048 673552 308100
rect 673604 308088 673610 308100
rect 676030 308088 676036 308100
rect 673604 308060 676036 308088
rect 673604 308048 673610 308060
rect 676030 308048 676036 308060
rect 676088 308048 676094 308100
rect 674466 306824 674472 306876
rect 674524 306864 674530 306876
rect 676030 306864 676036 306876
rect 674524 306836 676036 306864
rect 674524 306824 674530 306836
rect 676030 306824 676036 306836
rect 676088 306824 676094 306876
rect 673454 306484 673460 306536
rect 673512 306524 673518 306536
rect 675938 306524 675944 306536
rect 673512 306496 675944 306524
rect 673512 306484 673518 306496
rect 675938 306484 675944 306496
rect 675996 306484 676002 306536
rect 673914 306416 673920 306468
rect 673972 306456 673978 306468
rect 676122 306456 676128 306468
rect 673972 306428 676128 306456
rect 673972 306416 673978 306428
rect 676122 306416 676128 306428
rect 676180 306416 676186 306468
rect 676030 306388 676036 306400
rect 675128 306360 676036 306388
rect 675128 306264 675156 306360
rect 676030 306348 676036 306360
rect 676088 306348 676094 306400
rect 675110 306212 675116 306264
rect 675168 306212 675174 306264
rect 673730 305056 673736 305108
rect 673788 305096 673794 305108
rect 676122 305096 676128 305108
rect 673788 305068 676128 305096
rect 673788 305056 673794 305068
rect 676122 305056 676128 305068
rect 676180 305056 676186 305108
rect 674650 304784 674656 304836
rect 674708 304824 674714 304836
rect 676030 304824 676036 304836
rect 674708 304796 676036 304824
rect 674708 304784 674714 304796
rect 676030 304784 676036 304796
rect 676088 304784 676094 304836
rect 673822 304240 673828 304292
rect 673880 304280 673886 304292
rect 676122 304280 676128 304292
rect 673880 304252 676128 304280
rect 673880 304240 673886 304252
rect 676122 304240 676128 304252
rect 676180 304240 676186 304292
rect 673638 303764 673644 303816
rect 673696 303804 673702 303816
rect 675938 303804 675944 303816
rect 673696 303776 675944 303804
rect 673696 303764 673702 303776
rect 675938 303764 675944 303776
rect 675996 303764 676002 303816
rect 674006 303696 674012 303748
rect 674064 303736 674070 303748
rect 676122 303736 676128 303748
rect 674064 303708 676128 303736
rect 674064 303696 674070 303708
rect 676122 303696 676128 303708
rect 676180 303696 676186 303748
rect 674558 303628 674564 303680
rect 674616 303668 674622 303680
rect 676030 303668 676036 303680
rect 674616 303640 676036 303668
rect 674616 303628 674622 303640
rect 676030 303628 676036 303640
rect 676088 303628 676094 303680
rect 41506 301588 41512 301640
rect 41564 301628 41570 301640
rect 49142 301628 49148 301640
rect 41564 301600 49148 301628
rect 41564 301588 41570 301600
rect 49142 301588 49148 301600
rect 49200 301588 49206 301640
rect 41782 300908 41788 300960
rect 41840 300948 41846 300960
rect 51166 300948 51172 300960
rect 41840 300920 51172 300948
rect 41840 300908 41846 300920
rect 51166 300908 51172 300920
rect 51224 300908 51230 300960
rect 673086 300840 673092 300892
rect 673144 300880 673150 300892
rect 679066 300880 679072 300892
rect 673144 300852 679072 300880
rect 673144 300840 673150 300852
rect 679066 300840 679072 300852
rect 679124 300840 679130 300892
rect 656802 298392 656808 298444
rect 656860 298432 656866 298444
rect 669498 298432 669504 298444
rect 656860 298404 669504 298432
rect 656860 298392 656866 298404
rect 669498 298392 669504 298404
rect 669556 298392 669562 298444
rect 675754 296148 675760 296200
rect 675812 296148 675818 296200
rect 675772 295996 675800 296148
rect 675754 295944 675760 295996
rect 675812 295944 675818 295996
rect 675202 295060 675208 295112
rect 675260 295100 675266 295112
rect 675386 295100 675392 295112
rect 675260 295072 675392 295100
rect 675260 295060 675266 295072
rect 675386 295060 675392 295072
rect 675444 295060 675450 295112
rect 674190 294516 674196 294568
rect 674248 294556 674254 294568
rect 675386 294556 675392 294568
rect 674248 294528 675392 294556
rect 674248 294516 674254 294528
rect 675386 294516 675392 294528
rect 675444 294516 675450 294568
rect 674466 292884 674472 292936
rect 674524 292924 674530 292936
rect 675386 292924 675392 292936
rect 674524 292896 675392 292924
rect 674524 292884 674530 292896
rect 675386 292884 675392 292896
rect 675444 292884 675450 292936
rect 674650 291524 674656 291576
rect 674708 291564 674714 291576
rect 675386 291564 675392 291576
rect 674708 291536 675392 291564
rect 674708 291524 674714 291536
rect 675386 291524 675392 291536
rect 675444 291524 675450 291576
rect 674558 291048 674564 291100
rect 674616 291088 674622 291100
rect 675386 291088 675392 291100
rect 674616 291060 675392 291088
rect 674616 291048 674622 291060
rect 675386 291048 675392 291060
rect 675444 291048 675450 291100
rect 673914 288532 673920 288584
rect 673972 288572 673978 288584
rect 675386 288572 675392 288584
rect 673972 288544 675392 288572
rect 673972 288532 673978 288544
rect 675386 288532 675392 288544
rect 675444 288532 675450 288584
rect 674006 287920 674012 287972
rect 674064 287960 674070 287972
rect 675386 287960 675392 287972
rect 674064 287932 675392 287960
rect 674064 287920 674070 287932
rect 675386 287920 675392 287932
rect 675444 287920 675450 287972
rect 673822 287172 673828 287224
rect 673880 287212 673886 287224
rect 675478 287212 675484 287224
rect 673880 287184 675484 287212
rect 673880 287172 673886 287184
rect 675478 287172 675484 287184
rect 675536 287172 675542 287224
rect 35802 286968 35808 287020
rect 35860 287008 35866 287020
rect 42702 287008 42708 287020
rect 35860 286980 42708 287008
rect 35860 286968 35866 286980
rect 42702 286968 42708 286980
rect 42760 286968 42766 287020
rect 673638 286560 673644 286612
rect 673696 286600 673702 286612
rect 675386 286600 675392 286612
rect 673696 286572 675392 286600
rect 673696 286560 673702 286572
rect 675386 286560 675392 286572
rect 675444 286560 675450 286612
rect 32858 285744 32864 285796
rect 32916 285784 32922 285796
rect 42794 285784 42800 285796
rect 32916 285756 42800 285784
rect 32916 285744 32922 285756
rect 42794 285744 42800 285756
rect 42852 285744 42858 285796
rect 32950 285676 32956 285728
rect 33008 285716 33014 285728
rect 43254 285716 43260 285728
rect 33008 285688 43260 285716
rect 33008 285676 33014 285688
rect 43254 285676 43260 285688
rect 43312 285676 43318 285728
rect 32674 285608 32680 285660
rect 32732 285648 32738 285660
rect 41874 285648 41880 285660
rect 32732 285620 41880 285648
rect 32732 285608 32738 285620
rect 41874 285608 41880 285620
rect 41932 285608 41938 285660
rect 673730 285540 673736 285592
rect 673788 285580 673794 285592
rect 675478 285580 675484 285592
rect 673788 285552 675484 285580
rect 673788 285540 673794 285552
rect 675478 285540 675484 285552
rect 675536 285540 675542 285592
rect 655698 284724 655704 284776
rect 655756 284764 655762 284776
rect 670050 284764 670056 284776
rect 655756 284736 670056 284764
rect 655756 284724 655762 284736
rect 670050 284724 670056 284736
rect 670108 284724 670114 284776
rect 41874 283772 41880 283824
rect 41932 283772 41938 283824
rect 41892 283620 41920 283772
rect 673546 283704 673552 283756
rect 673604 283744 673610 283756
rect 675478 283744 675484 283756
rect 673604 283716 675484 283744
rect 673604 283704 673610 283716
rect 675478 283704 675484 283716
rect 675536 283704 675542 283756
rect 41874 283568 41880 283620
rect 41932 283568 41938 283620
rect 673454 281868 673460 281920
rect 673512 281908 673518 281920
rect 675386 281908 675392 281920
rect 673512 281880 675392 281908
rect 673512 281868 673518 281880
rect 675386 281868 675392 281880
rect 675444 281868 675450 281920
rect 42150 281732 42156 281784
rect 42208 281772 42214 281784
rect 42702 281772 42708 281784
rect 42208 281744 42708 281772
rect 42208 281732 42214 281744
rect 42702 281732 42708 281744
rect 42760 281732 42766 281784
rect 42150 281052 42156 281104
rect 42208 281092 42214 281104
rect 49050 281092 49056 281104
rect 42208 281064 49056 281092
rect 42208 281052 42214 281064
rect 49050 281052 49056 281064
rect 49108 281052 49114 281104
rect 42150 279828 42156 279880
rect 42208 279868 42214 279880
rect 42978 279868 42984 279880
rect 42208 279840 42984 279868
rect 42208 279828 42214 279840
rect 42978 279828 42984 279840
rect 43036 279828 43042 279880
rect 42058 278604 42064 278656
rect 42116 278644 42122 278656
rect 43346 278644 43352 278656
rect 42116 278616 43352 278644
rect 42116 278604 42122 278616
rect 43346 278604 43352 278616
rect 43404 278604 43410 278656
rect 46474 278536 46480 278588
rect 46532 278576 46538 278588
rect 670602 278576 670608 278588
rect 46532 278548 670608 278576
rect 46532 278536 46538 278548
rect 670602 278536 670608 278548
rect 670660 278536 670666 278588
rect 46566 278468 46572 278520
rect 46624 278508 46630 278520
rect 670418 278508 670424 278520
rect 46624 278480 670424 278508
rect 46624 278468 46630 278480
rect 670418 278468 670424 278480
rect 670476 278468 670482 278520
rect 62574 278400 62580 278452
rect 62632 278440 62638 278452
rect 670510 278440 670516 278452
rect 62632 278412 670516 278440
rect 62632 278400 62638 278412
rect 670510 278400 670516 278412
rect 670568 278400 670574 278452
rect 62022 278332 62028 278384
rect 62080 278372 62086 278384
rect 669866 278372 669872 278384
rect 62080 278344 669872 278372
rect 62080 278332 62086 278344
rect 669866 278332 669872 278344
rect 669924 278332 669930 278384
rect 62390 278264 62396 278316
rect 62448 278304 62454 278316
rect 670142 278304 670148 278316
rect 62448 278276 670148 278304
rect 62448 278264 62454 278276
rect 670142 278264 670148 278276
rect 670200 278264 670206 278316
rect 62758 278196 62764 278248
rect 62816 278236 62822 278248
rect 670326 278236 670332 278248
rect 62816 278208 670332 278236
rect 62816 278196 62822 278208
rect 670326 278196 670332 278208
rect 670384 278196 670390 278248
rect 62942 278128 62948 278180
rect 63000 278168 63006 278180
rect 668578 278168 668584 278180
rect 63000 278140 668584 278168
rect 63000 278128 63006 278140
rect 668578 278128 668584 278140
rect 668636 278128 668642 278180
rect 63310 278060 63316 278112
rect 63368 278100 63374 278112
rect 669958 278100 669964 278112
rect 63368 278072 669964 278100
rect 63368 278060 63374 278072
rect 669958 278060 669964 278072
rect 670016 278060 670022 278112
rect 42150 277992 42156 278044
rect 42208 278032 42214 278044
rect 43162 278032 43168 278044
rect 42208 278004 43168 278032
rect 42208 277992 42214 278004
rect 43162 277992 43168 278004
rect 43220 277992 43226 278044
rect 63126 277992 63132 278044
rect 63184 278032 63190 278044
rect 669774 278032 669780 278044
rect 63184 278004 669780 278032
rect 63184 277992 63190 278004
rect 669774 277992 669780 278004
rect 669832 277992 669838 278044
rect 42150 277380 42156 277432
rect 42208 277420 42214 277432
rect 43622 277420 43628 277432
rect 42208 277392 43628 277420
rect 42208 277380 42214 277392
rect 43622 277380 43628 277392
rect 43680 277380 43686 277432
rect 42058 276700 42064 276752
rect 42116 276740 42122 276752
rect 42794 276740 42800 276752
rect 42116 276712 42800 276740
rect 42116 276700 42122 276712
rect 42794 276700 42800 276712
rect 42852 276700 42858 276752
rect 345106 275952 345112 276004
rect 345164 275992 345170 276004
rect 471330 275992 471336 276004
rect 345164 275964 471336 275992
rect 345164 275952 345170 275964
rect 471330 275952 471336 275964
rect 471388 275952 471394 276004
rect 343726 275884 343732 275936
rect 343784 275924 343790 275936
rect 467834 275924 467840 275936
rect 343784 275896 467840 275924
rect 343784 275884 343790 275896
rect 467834 275884 467840 275896
rect 467892 275884 467898 275936
rect 349062 275816 349068 275868
rect 349120 275856 349126 275868
rect 482002 275856 482008 275868
rect 349120 275828 482008 275856
rect 349120 275816 349126 275828
rect 482002 275816 482008 275828
rect 482060 275816 482066 275868
rect 350166 275748 350172 275800
rect 350224 275788 350230 275800
rect 485498 275788 485504 275800
rect 350224 275760 485504 275788
rect 350224 275748 350230 275760
rect 485498 275748 485504 275760
rect 485556 275748 485562 275800
rect 354398 275680 354404 275732
rect 354456 275720 354462 275732
rect 496170 275720 496176 275732
rect 354456 275692 496176 275720
rect 354456 275680 354462 275692
rect 496170 275680 496176 275692
rect 496228 275680 496234 275732
rect 355778 275612 355784 275664
rect 355836 275652 355842 275664
rect 499758 275652 499764 275664
rect 355836 275624 499764 275652
rect 355836 275612 355842 275624
rect 499758 275612 499764 275624
rect 499816 275612 499822 275664
rect 358446 275544 358452 275596
rect 358504 275584 358510 275596
rect 506842 275584 506848 275596
rect 358504 275556 506848 275584
rect 358504 275544 358510 275556
rect 506842 275544 506848 275556
rect 506900 275544 506906 275596
rect 361114 275476 361120 275528
rect 361172 275516 361178 275528
rect 513926 275516 513932 275528
rect 361172 275488 513932 275516
rect 361172 275476 361178 275488
rect 513926 275476 513932 275488
rect 513984 275476 513990 275528
rect 364058 275408 364064 275460
rect 364116 275448 364122 275460
rect 521010 275448 521016 275460
rect 364116 275420 521016 275448
rect 364116 275408 364122 275420
rect 521010 275408 521016 275420
rect 521068 275408 521074 275460
rect 366450 275340 366456 275392
rect 366508 275380 366514 275392
rect 528094 275380 528100 275392
rect 366508 275352 528100 275380
rect 366508 275340 366514 275352
rect 528094 275340 528100 275352
rect 528152 275340 528158 275392
rect 369118 275272 369124 275324
rect 369176 275312 369182 275324
rect 535178 275312 535184 275324
rect 369176 275284 535184 275312
rect 369176 275272 369182 275284
rect 535178 275272 535184 275284
rect 535236 275272 535242 275324
rect 371786 275204 371792 275256
rect 371844 275244 371850 275256
rect 542262 275244 542268 275256
rect 371844 275216 542268 275244
rect 371844 275204 371850 275216
rect 542262 275204 542268 275216
rect 542320 275204 542326 275256
rect 374914 275136 374920 275188
rect 374972 275176 374978 275188
rect 550542 275176 550548 275188
rect 374972 275148 550548 275176
rect 374972 275136 374978 275148
rect 550542 275136 550548 275148
rect 550600 275136 550606 275188
rect 377582 275068 377588 275120
rect 377640 275108 377646 275120
rect 557626 275108 557632 275120
rect 377640 275080 557632 275108
rect 377640 275068 377646 275080
rect 557626 275068 557632 275080
rect 557684 275068 557690 275120
rect 380250 275000 380256 275052
rect 380308 275040 380314 275052
rect 564710 275040 564716 275052
rect 380308 275012 564716 275040
rect 380308 275000 380314 275012
rect 564710 275000 564716 275012
rect 564768 275000 564774 275052
rect 382918 274932 382924 274984
rect 382976 274972 382982 274984
rect 571794 274972 571800 274984
rect 382976 274944 571800 274972
rect 382976 274932 382982 274944
rect 571794 274932 571800 274944
rect 571852 274932 571858 274984
rect 385586 274864 385592 274916
rect 385644 274904 385650 274916
rect 578878 274904 578884 274916
rect 385644 274876 578884 274904
rect 385644 274864 385650 274876
rect 578878 274864 578884 274876
rect 578936 274864 578942 274916
rect 318886 274796 318892 274848
rect 318944 274836 318950 274848
rect 401594 274836 401600 274848
rect 318944 274808 401600 274836
rect 318944 274796 318950 274808
rect 401594 274796 401600 274808
rect 401652 274796 401658 274848
rect 403894 274796 403900 274848
rect 403952 274836 403958 274848
rect 403952 274808 420868 274836
rect 403952 274796 403958 274808
rect 320174 274728 320180 274780
rect 320232 274768 320238 274780
rect 405182 274768 405188 274780
rect 320232 274740 405188 274768
rect 320232 274728 320238 274740
rect 405182 274728 405188 274740
rect 405240 274728 405246 274780
rect 406562 274728 406568 274780
rect 406620 274768 406626 274780
rect 420840 274768 420868 274808
rect 420914 274796 420920 274848
rect 420972 274836 420978 274848
rect 620278 274836 620284 274848
rect 420972 274808 620284 274836
rect 420972 274796 420978 274808
rect 620278 274796 620284 274808
rect 620336 274796 620342 274848
rect 627362 274768 627368 274780
rect 406620 274740 414980 274768
rect 420840 274740 627368 274768
rect 406620 274728 406626 274740
rect 321002 274660 321008 274712
rect 321060 274700 321066 274712
rect 407482 274700 407488 274712
rect 321060 274672 407488 274700
rect 321060 274660 321066 274672
rect 407482 274660 407488 274672
rect 407540 274660 407546 274712
rect 409230 274660 409236 274712
rect 409288 274700 409294 274712
rect 414952 274700 414980 274740
rect 627362 274728 627368 274740
rect 627420 274728 627426 274780
rect 634446 274700 634452 274712
rect 409288 274672 411208 274700
rect 414952 274672 634452 274700
rect 409288 274660 409294 274672
rect 322750 274592 322756 274644
rect 322808 274632 322814 274644
rect 411070 274632 411076 274644
rect 322808 274604 411076 274632
rect 322808 274592 322814 274604
rect 411070 274592 411076 274604
rect 411128 274592 411134 274644
rect 411180 274632 411208 274672
rect 634446 274660 634452 274672
rect 634504 274660 634510 274712
rect 641622 274632 641628 274644
rect 411180 274604 641628 274632
rect 641622 274592 641628 274604
rect 641680 274592 641686 274644
rect 342530 274524 342536 274576
rect 342588 274564 342594 274576
rect 464246 274564 464252 274576
rect 342588 274536 464252 274564
rect 342588 274524 342594 274536
rect 464246 274524 464252 274536
rect 464304 274524 464310 274576
rect 341058 274456 341064 274508
rect 341116 274496 341122 274508
rect 460658 274496 460664 274508
rect 341116 274468 460664 274496
rect 341116 274456 341122 274468
rect 460658 274456 460664 274468
rect 460716 274456 460722 274508
rect 337102 274388 337108 274440
rect 337160 274428 337166 274440
rect 450078 274428 450084 274440
rect 337160 274400 450084 274428
rect 337160 274388 337166 274400
rect 450078 274388 450084 274400
rect 450136 274388 450142 274440
rect 336090 274320 336096 274372
rect 336148 274360 336154 274372
rect 446490 274360 446496 274372
rect 336148 274332 446496 274360
rect 336148 274320 336154 274332
rect 446490 274320 446496 274332
rect 446548 274320 446554 274372
rect 42150 274252 42156 274304
rect 42208 274292 42214 274304
rect 43070 274292 43076 274304
rect 42208 274264 43076 274292
rect 42208 274252 42214 274264
rect 43070 274252 43076 274264
rect 43128 274252 43134 274304
rect 333146 274252 333152 274304
rect 333204 274292 333210 274304
rect 439406 274292 439412 274304
rect 333204 274264 439412 274292
rect 333204 274252 333210 274264
rect 439406 274252 439412 274264
rect 439464 274252 439470 274304
rect 334342 274184 334348 274236
rect 334400 274224 334406 274236
rect 442994 274224 443000 274236
rect 334400 274196 443000 274224
rect 334400 274184 334406 274196
rect 442994 274184 443000 274196
rect 443052 274184 443058 274236
rect 332134 274116 332140 274168
rect 332192 274156 332198 274168
rect 437014 274156 437020 274168
rect 332192 274128 437020 274156
rect 332192 274116 332198 274128
rect 437014 274116 437020 274128
rect 437072 274116 437078 274168
rect 351822 274048 351828 274100
rect 351880 274088 351886 274100
rect 432322 274088 432328 274100
rect 351880 274060 432328 274088
rect 351880 274048 351886 274060
rect 432322 274048 432328 274060
rect 432380 274048 432386 274100
rect 331674 273980 331680 274032
rect 331732 274020 331738 274032
rect 435910 274020 435916 274032
rect 331732 273992 435916 274020
rect 331732 273980 331738 273992
rect 435910 273980 435916 273992
rect 435968 273980 435974 274032
rect 327718 273912 327724 273964
rect 327776 273952 327782 273964
rect 425238 273952 425244 273964
rect 327776 273924 425244 273952
rect 327776 273912 327782 273924
rect 425238 273912 425244 273924
rect 425296 273912 425302 273964
rect 329006 273844 329012 273896
rect 329064 273884 329070 273896
rect 428826 273884 428832 273896
rect 329064 273856 428832 273884
rect 329064 273844 329070 273856
rect 428826 273844 428832 273856
rect 428884 273844 428890 273896
rect 326798 273776 326804 273828
rect 326856 273816 326862 273828
rect 422846 273816 422852 273828
rect 326856 273788 422852 273816
rect 326856 273776 326862 273788
rect 422846 273776 422852 273788
rect 422904 273776 422910 273828
rect 42058 273708 42064 273760
rect 42116 273748 42122 273760
rect 42886 273748 42892 273760
rect 42116 273720 42892 273748
rect 42116 273708 42122 273720
rect 42886 273708 42892 273720
rect 42944 273708 42950 273760
rect 325418 273708 325424 273760
rect 325476 273748 325482 273760
rect 418154 273748 418160 273760
rect 325476 273720 418160 273748
rect 325476 273708 325482 273720
rect 418154 273708 418160 273720
rect 418212 273708 418218 273760
rect 326338 273640 326344 273692
rect 326396 273680 326402 273692
rect 326396 273652 409828 273680
rect 326396 273640 326402 273652
rect 323670 273572 323676 273624
rect 323728 273612 323734 273624
rect 409800 273612 409828 273652
rect 421650 273612 421656 273624
rect 323728 273584 400214 273612
rect 409800 273584 421656 273612
rect 323728 273572 323734 273584
rect 330386 273504 330392 273556
rect 330444 273544 330450 273556
rect 351822 273544 351828 273556
rect 330444 273516 351828 273544
rect 330444 273504 330450 273516
rect 351822 273504 351828 273516
rect 351880 273504 351886 273556
rect 400186 273544 400214 273584
rect 421650 273572 421656 273584
rect 421708 273572 421714 273624
rect 414566 273544 414572 273556
rect 400186 273516 414572 273544
rect 414566 273504 414572 273516
rect 414624 273504 414630 273556
rect 401134 273436 401140 273488
rect 401192 273476 401198 273488
rect 420914 273476 420920 273488
rect 401192 273448 420920 273476
rect 401192 273436 401198 273448
rect 420914 273436 420920 273448
rect 420972 273436 420978 273488
rect 226150 273204 226156 273216
rect 168346 273176 226156 273204
rect 155678 273096 155684 273148
rect 155736 273136 155742 273148
rect 168346 273136 168374 273176
rect 226150 273164 226156 273176
rect 226208 273164 226214 273216
rect 263226 273164 263232 273216
rect 263284 273204 263290 273216
rect 266722 273204 266728 273216
rect 263284 273176 266728 273204
rect 263284 273164 263290 273176
rect 266722 273164 266728 273176
rect 266780 273164 266786 273216
rect 292022 273164 292028 273216
rect 292080 273204 292086 273216
rect 329466 273204 329472 273216
rect 292080 273176 329472 273204
rect 292080 273164 292086 273176
rect 329466 273164 329472 273176
rect 329524 273164 329530 273216
rect 339494 273164 339500 273216
rect 339552 273204 339558 273216
rect 344830 273204 344836 273216
rect 339552 273176 344836 273204
rect 339552 273164 339558 273176
rect 344830 273164 344836 273176
rect 344888 273164 344894 273216
rect 354858 273164 354864 273216
rect 354916 273204 354922 273216
rect 354916 273176 362908 273204
rect 354916 273164 354922 273176
rect 155736 273108 168374 273136
rect 155736 273096 155742 273108
rect 177850 273096 177856 273148
rect 177908 273136 177914 273148
rect 227070 273136 227076 273148
rect 177908 273108 227076 273136
rect 177908 273096 177914 273108
rect 227070 273096 227076 273108
rect 227128 273096 227134 273148
rect 264422 273096 264428 273148
rect 264480 273136 264486 273148
rect 267182 273136 267188 273148
rect 264480 273108 267188 273136
rect 264480 273096 264486 273108
rect 267182 273096 267188 273108
rect 267240 273096 267246 273148
rect 292574 273096 292580 273148
rect 292632 273136 292638 273148
rect 331858 273136 331864 273148
rect 292632 273108 331864 273136
rect 292632 273096 292638 273108
rect 331858 273096 331864 273108
rect 331916 273096 331922 273148
rect 355318 273096 355324 273148
rect 355376 273136 355382 273148
rect 362880 273136 362908 273176
rect 362954 273164 362960 273216
rect 363012 273204 363018 273216
rect 491478 273204 491484 273216
rect 363012 273176 491484 273204
rect 363012 273164 363018 273176
rect 491478 273164 491484 273176
rect 491536 273164 491542 273216
rect 497366 273136 497372 273148
rect 355376 273108 362816 273136
rect 362880 273108 497372 273136
rect 355376 273096 355382 273108
rect 148594 273028 148600 273080
rect 148652 273068 148658 273080
rect 223482 273068 223488 273080
rect 148652 273040 223488 273068
rect 148652 273028 148658 273040
rect 223482 273028 223488 273040
rect 223540 273028 223546 273080
rect 243170 273028 243176 273080
rect 243228 273068 243234 273080
rect 259178 273068 259184 273080
rect 243228 273040 259184 273068
rect 243228 273028 243234 273040
rect 259178 273028 259184 273040
rect 259236 273028 259242 273080
rect 260926 273028 260932 273080
rect 260984 273068 260990 273080
rect 265802 273068 265808 273080
rect 260984 273040 265808 273068
rect 260984 273028 260990 273040
rect 265802 273028 265808 273040
rect 265860 273028 265866 273080
rect 293862 273028 293868 273080
rect 293920 273068 293926 273080
rect 335354 273068 335360 273080
rect 293920 273040 335360 273068
rect 293920 273028 293926 273040
rect 335354 273028 335360 273040
rect 335412 273028 335418 273080
rect 358814 273028 358820 273080
rect 358872 273068 358878 273080
rect 362788 273068 362816 273108
rect 497366 273096 497372 273108
rect 497424 273096 497430 273148
rect 498562 273068 498568 273080
rect 358872 273040 362724 273068
rect 362788 273040 498568 273068
rect 358872 273028 358878 273040
rect 149790 272960 149796 273012
rect 149848 273000 149854 273012
rect 224402 273000 224408 273012
rect 149848 272972 224408 273000
rect 149848 272960 149854 272972
rect 224402 272960 224408 272972
rect 224460 272960 224466 273012
rect 241974 272960 241980 273012
rect 242032 273000 242038 273012
rect 258718 273000 258724 273012
rect 242032 272972 258724 273000
rect 242032 272960 242038 272972
rect 258718 272960 258724 272972
rect 258776 272960 258782 273012
rect 293402 272960 293408 273012
rect 293460 273000 293466 273012
rect 334158 273000 334164 273012
rect 293460 272972 334164 273000
rect 293460 272960 293466 272972
rect 334158 272960 334164 272972
rect 334216 272960 334222 273012
rect 344002 272960 344008 273012
rect 344060 273000 344066 273012
rect 362586 273000 362592 273012
rect 344060 272972 362592 273000
rect 344060 272960 344066 272972
rect 362586 272960 362592 272972
rect 362644 272960 362650 273012
rect 362696 273000 362724 273040
rect 498562 273028 498568 273040
rect 498620 273028 498626 273080
rect 498838 273028 498844 273080
rect 498896 273068 498902 273080
rect 617978 273068 617984 273080
rect 498896 273040 617984 273068
rect 498896 273028 498902 273040
rect 617978 273028 617984 273040
rect 618036 273028 618042 273080
rect 504450 273000 504456 273012
rect 362696 272972 504456 273000
rect 504450 272960 504456 272972
rect 504508 272960 504514 273012
rect 42150 272892 42156 272944
rect 42208 272932 42214 272944
rect 43254 272932 43260 272944
rect 42208 272904 43260 272932
rect 42208 272892 42214 272904
rect 43254 272892 43260 272904
rect 43312 272892 43318 272944
rect 150986 272892 150992 272944
rect 151044 272932 151050 272944
rect 223942 272932 223948 272944
rect 151044 272904 223948 272932
rect 151044 272892 151050 272904
rect 223942 272892 223948 272904
rect 224000 272892 224006 272944
rect 239582 272892 239588 272944
rect 239640 272932 239646 272944
rect 257798 272932 257804 272944
rect 239640 272904 257804 272932
rect 239640 272892 239646 272904
rect 257798 272892 257804 272904
rect 257856 272892 257862 272944
rect 304902 272892 304908 272944
rect 304960 272932 304966 272944
rect 346026 272932 346032 272944
rect 304960 272904 346032 272932
rect 304960 272892 304966 272904
rect 346026 272892 346032 272904
rect 346084 272892 346090 272944
rect 357986 272892 357992 272944
rect 358044 272932 358050 272944
rect 505646 272932 505652 272944
rect 358044 272904 505652 272932
rect 358044 272892 358050 272904
rect 505646 272892 505652 272904
rect 505704 272892 505710 272944
rect 143902 272824 143908 272876
rect 143960 272864 143966 272876
rect 221274 272864 221280 272876
rect 143960 272836 221280 272864
rect 143960 272824 143966 272836
rect 221274 272824 221280 272836
rect 221332 272824 221338 272876
rect 236086 272824 236092 272876
rect 236144 272864 236150 272876
rect 256418 272864 256424 272876
rect 236144 272836 256424 272864
rect 236144 272824 236150 272836
rect 256418 272824 256424 272836
rect 256476 272824 256482 272876
rect 307846 272824 307852 272876
rect 307904 272864 307910 272876
rect 348418 272864 348424 272876
rect 307904 272836 348424 272864
rect 307904 272824 307910 272836
rect 348418 272824 348424 272836
rect 348476 272824 348482 272876
rect 360654 272824 360660 272876
rect 360712 272864 360718 272876
rect 512730 272864 512736 272876
rect 360712 272836 512736 272864
rect 360712 272824 360718 272836
rect 512730 272824 512736 272836
rect 512788 272824 512794 272876
rect 145006 272756 145012 272808
rect 145064 272796 145070 272808
rect 222194 272796 222200 272808
rect 145064 272768 222200 272796
rect 145064 272756 145070 272768
rect 222194 272756 222200 272768
rect 222252 272756 222258 272808
rect 234890 272756 234896 272808
rect 234948 272796 234954 272808
rect 256050 272796 256056 272808
rect 234948 272768 256056 272796
rect 234948 272756 234954 272768
rect 256050 272756 256056 272768
rect 256108 272756 256114 272808
rect 300762 272756 300768 272808
rect 300820 272796 300826 272808
rect 353110 272796 353116 272808
rect 300820 272768 353116 272796
rect 300820 272756 300826 272768
rect 353110 272756 353116 272768
rect 353168 272756 353174 272808
rect 360562 272756 360568 272808
rect 360620 272796 360626 272808
rect 511534 272796 511540 272808
rect 360620 272768 511540 272796
rect 360620 272756 360626 272768
rect 511534 272756 511540 272768
rect 511592 272756 511598 272808
rect 511626 272756 511632 272808
rect 511684 272796 511690 272808
rect 610802 272796 610808 272808
rect 511684 272768 610808 272796
rect 511684 272756 511690 272768
rect 610802 272756 610808 272768
rect 610860 272756 610866 272808
rect 146202 272688 146208 272740
rect 146260 272728 146266 272740
rect 223022 272728 223028 272740
rect 146260 272700 223028 272728
rect 146260 272688 146266 272700
rect 223022 272688 223028 272700
rect 223080 272688 223086 272740
rect 232498 272688 232504 272740
rect 232556 272728 232562 272740
rect 255130 272728 255136 272740
rect 232556 272700 255136 272728
rect 232556 272688 232562 272700
rect 255130 272688 255136 272700
rect 255188 272688 255194 272740
rect 294874 272688 294880 272740
rect 294932 272728 294938 272740
rect 338942 272728 338948 272740
rect 294932 272700 338948 272728
rect 294932 272688 294938 272700
rect 338942 272688 338948 272700
rect 339000 272688 339006 272740
rect 344738 272688 344744 272740
rect 344796 272728 344802 272740
rect 470134 272728 470140 272740
rect 344796 272700 470140 272728
rect 344796 272688 344802 272700
rect 470134 272688 470140 272700
rect 470192 272688 470198 272740
rect 471974 272688 471980 272740
rect 472032 272728 472038 272740
rect 625062 272728 625068 272740
rect 472032 272700 625068 272728
rect 472032 272688 472038 272700
rect 625062 272688 625068 272700
rect 625120 272688 625126 272740
rect 139118 272620 139124 272672
rect 139176 272660 139182 272672
rect 220354 272660 220360 272672
rect 139176 272632 220360 272660
rect 139176 272620 139182 272632
rect 220354 272620 220360 272632
rect 220412 272620 220418 272672
rect 237282 272620 237288 272672
rect 237340 272660 237346 272672
rect 257154 272660 257160 272672
rect 237340 272632 257160 272660
rect 237340 272620 237346 272632
rect 257154 272620 257160 272632
rect 257212 272620 257218 272672
rect 301406 272620 301412 272672
rect 301464 272660 301470 272672
rect 355502 272660 355508 272672
rect 301464 272632 355508 272660
rect 301464 272620 301470 272632
rect 355502 272620 355508 272632
rect 355560 272620 355566 272672
rect 363138 272620 363144 272672
rect 363196 272660 363202 272672
rect 518618 272660 518624 272672
rect 363196 272632 518624 272660
rect 363196 272620 363202 272632
rect 518618 272620 518624 272632
rect 518676 272620 518682 272672
rect 137922 272552 137928 272604
rect 137980 272592 137986 272604
rect 219158 272592 219164 272604
rect 137980 272564 219164 272592
rect 137980 272552 137986 272564
rect 219158 272552 219164 272564
rect 219216 272552 219222 272604
rect 233694 272552 233700 272604
rect 233752 272592 233758 272604
rect 255590 272592 255596 272604
rect 233752 272564 255596 272592
rect 233752 272552 233758 272564
rect 255590 272552 255596 272564
rect 255648 272552 255654 272604
rect 300670 272552 300676 272604
rect 300728 272592 300734 272604
rect 351914 272592 351920 272604
rect 300728 272564 351920 272592
rect 300728 272552 300734 272564
rect 351914 272552 351920 272564
rect 351972 272552 351978 272604
rect 353110 272552 353116 272604
rect 353168 272592 353174 272604
rect 362954 272592 362960 272604
rect 353168 272564 362960 272592
rect 353168 272552 353174 272564
rect 362954 272552 362960 272564
rect 363012 272552 363018 272604
rect 368198 272552 368204 272604
rect 368256 272592 368262 272604
rect 532786 272592 532792 272604
rect 368256 272564 532792 272592
rect 368256 272552 368262 272564
rect 532786 272552 532792 272564
rect 532844 272552 532850 272604
rect 136818 272484 136824 272536
rect 136876 272524 136882 272536
rect 218606 272524 218612 272536
rect 136876 272496 218612 272524
rect 136876 272484 136882 272496
rect 218606 272484 218612 272496
rect 218664 272484 218670 272536
rect 230198 272484 230204 272536
rect 230256 272524 230262 272536
rect 254210 272524 254216 272536
rect 230256 272496 254216 272524
rect 230256 272484 230262 272496
rect 254210 272484 254216 272496
rect 254268 272484 254274 272536
rect 296070 272484 296076 272536
rect 296128 272524 296134 272536
rect 341334 272524 341340 272536
rect 296128 272496 341340 272524
rect 296128 272484 296134 272496
rect 341334 272484 341340 272496
rect 341392 272484 341398 272536
rect 342070 272484 342076 272536
rect 342128 272524 342134 272536
rect 463050 272524 463056 272536
rect 342128 272496 463056 272524
rect 342128 272484 342134 272496
rect 463050 272484 463056 272496
rect 463108 272484 463114 272536
rect 465902 272484 465908 272536
rect 465960 272524 465966 272536
rect 632146 272524 632152 272536
rect 465960 272496 632152 272524
rect 465960 272484 465966 272496
rect 632146 272484 632152 272496
rect 632204 272484 632210 272536
rect 132034 272416 132040 272468
rect 132092 272456 132098 272468
rect 217686 272456 217692 272468
rect 132092 272428 217692 272456
rect 132092 272416 132098 272428
rect 217686 272416 217692 272428
rect 217744 272416 217750 272468
rect 301866 272416 301872 272468
rect 301924 272456 301930 272468
rect 356698 272456 356704 272468
rect 301924 272428 356704 272456
rect 301924 272416 301930 272428
rect 356698 272416 356704 272428
rect 356756 272416 356762 272468
rect 373166 272416 373172 272468
rect 373224 272456 373230 272468
rect 545850 272456 545856 272468
rect 373224 272428 545856 272456
rect 373224 272416 373230 272428
rect 545850 272416 545856 272428
rect 545908 272416 545914 272468
rect 124950 272348 124956 272400
rect 125008 272388 125014 272400
rect 215018 272388 215024 272400
rect 125008 272360 215024 272388
rect 125008 272348 125014 272360
rect 215018 272348 215024 272360
rect 215076 272348 215082 272400
rect 303338 272348 303344 272400
rect 303396 272388 303402 272400
rect 360194 272388 360200 272400
rect 303396 272360 360200 272388
rect 303396 272348 303402 272360
rect 360194 272348 360200 272360
rect 360252 272348 360258 272400
rect 376662 272348 376668 272400
rect 376720 272388 376726 272400
rect 555234 272388 555240 272400
rect 376720 272360 555240 272388
rect 376720 272348 376726 272360
rect 555234 272348 555240 272360
rect 555292 272348 555298 272400
rect 129642 272280 129648 272332
rect 129700 272320 129706 272332
rect 215662 272320 215668 272332
rect 129700 272292 215668 272320
rect 129700 272280 129706 272292
rect 215662 272280 215668 272292
rect 215720 272280 215726 272332
rect 294782 272280 294788 272332
rect 294840 272320 294846 272332
rect 337746 272320 337752 272332
rect 294840 272292 337752 272320
rect 294840 272280 294846 272292
rect 337746 272280 337752 272292
rect 337804 272280 337810 272332
rect 339310 272280 339316 272332
rect 339368 272320 339374 272332
rect 455966 272320 455972 272332
rect 339368 272292 455972 272320
rect 339368 272280 339374 272292
rect 455966 272280 455972 272292
rect 456024 272280 456030 272332
rect 459462 272280 459468 272332
rect 459520 272320 459526 272332
rect 639230 272320 639236 272332
rect 459520 272292 639236 272320
rect 459520 272280 459526 272292
rect 639230 272280 639236 272292
rect 639288 272280 639294 272332
rect 117866 272212 117872 272264
rect 117924 272252 117930 272264
rect 206646 272252 206652 272264
rect 117924 272224 206652 272252
rect 117924 272212 117930 272224
rect 206646 272212 206652 272224
rect 206704 272212 206710 272264
rect 302786 272212 302792 272264
rect 302844 272252 302850 272264
rect 358998 272252 359004 272264
rect 302844 272224 359004 272252
rect 302844 272212 302850 272224
rect 358998 272212 359004 272224
rect 359056 272212 359062 272264
rect 381998 272212 382004 272264
rect 382056 272252 382062 272264
rect 569494 272252 569500 272264
rect 382056 272224 569500 272252
rect 382056 272212 382062 272224
rect 569494 272212 569500 272224
rect 569552 272212 569558 272264
rect 93026 272144 93032 272196
rect 93084 272184 93090 272196
rect 184934 272184 184940 272196
rect 93084 272156 184940 272184
rect 93084 272144 93090 272156
rect 184934 272144 184940 272156
rect 184992 272144 184998 272196
rect 188798 272144 188804 272196
rect 188856 272184 188862 272196
rect 234614 272184 234620 272196
rect 188856 272156 234620 272184
rect 188856 272144 188862 272156
rect 234614 272144 234620 272156
rect 234672 272144 234678 272196
rect 238478 272144 238484 272196
rect 238536 272184 238542 272196
rect 257246 272184 257252 272196
rect 238536 272156 257252 272184
rect 238536 272144 238542 272156
rect 257246 272144 257252 272156
rect 257304 272144 257310 272196
rect 306282 272144 306288 272196
rect 306340 272184 306346 272196
rect 367278 272184 367284 272196
rect 306340 272156 367284 272184
rect 306340 272144 306346 272156
rect 367278 272144 367284 272156
rect 367336 272144 367342 272196
rect 384666 272144 384672 272196
rect 384724 272184 384730 272196
rect 576578 272184 576584 272196
rect 384724 272156 576584 272184
rect 384724 272144 384730 272156
rect 576578 272144 576584 272156
rect 576636 272144 576642 272196
rect 104894 272076 104900 272128
rect 104952 272116 104958 272128
rect 202782 272116 202788 272128
rect 104952 272088 202788 272116
rect 104952 272076 104958 272088
rect 202782 272076 202788 272088
rect 202840 272076 202846 272128
rect 205358 272076 205364 272128
rect 205416 272116 205422 272128
rect 240134 272116 240140 272128
rect 205416 272088 240140 272116
rect 205416 272076 205422 272088
rect 240134 272076 240140 272088
rect 240192 272076 240198 272128
rect 308950 272076 308956 272128
rect 309008 272116 309014 272128
rect 374362 272116 374368 272128
rect 309008 272088 374368 272116
rect 309008 272076 309014 272088
rect 374362 272076 374368 272088
rect 374420 272076 374426 272128
rect 387334 272076 387340 272128
rect 387392 272116 387398 272128
rect 583662 272116 583668 272128
rect 387392 272088 583668 272116
rect 387392 272076 387398 272088
rect 583662 272076 583668 272088
rect 583720 272076 583726 272128
rect 89530 272008 89536 272060
rect 89588 272048 89594 272060
rect 178034 272048 178040 272060
rect 89588 272020 178040 272048
rect 89588 272008 89594 272020
rect 178034 272008 178040 272020
rect 178092 272008 178098 272060
rect 178126 272008 178132 272060
rect 178184 272048 178190 272060
rect 197262 272048 197268 272060
rect 178184 272020 197268 272048
rect 178184 272008 178190 272020
rect 197262 272008 197268 272020
rect 197320 272008 197326 272060
rect 199470 272008 199476 272060
rect 199528 272048 199534 272060
rect 242618 272048 242624 272060
rect 199528 272020 242624 272048
rect 199528 272008 199534 272020
rect 242618 272008 242624 272020
rect 242676 272008 242682 272060
rect 284202 272008 284208 272060
rect 284260 272048 284266 272060
rect 309410 272048 309416 272060
rect 284260 272020 309416 272048
rect 284260 272008 284266 272020
rect 309410 272008 309416 272020
rect 309468 272008 309474 272060
rect 311618 272008 311624 272060
rect 311676 272048 311682 272060
rect 381538 272048 381544 272060
rect 311676 272020 381544 272048
rect 311676 272008 311682 272020
rect 381538 272008 381544 272020
rect 381596 272008 381602 272060
rect 394602 272008 394608 272060
rect 394660 272048 394666 272060
rect 590746 272048 590752 272060
rect 394660 272020 590752 272048
rect 394660 272008 394666 272020
rect 590746 272008 590752 272020
rect 590804 272008 590810 272060
rect 75270 271940 75276 271992
rect 75328 271980 75334 271992
rect 195422 271980 195428 271992
rect 75328 271952 195428 271980
rect 75328 271940 75334 271952
rect 195422 271940 195428 271952
rect 195480 271940 195486 271992
rect 201770 271940 201776 271992
rect 201828 271980 201834 271992
rect 243538 271980 243544 271992
rect 201828 271952 243544 271980
rect 201828 271940 201834 271952
rect 243538 271940 243544 271952
rect 243596 271940 243602 271992
rect 285398 271940 285404 271992
rect 285456 271980 285462 271992
rect 312906 271980 312912 271992
rect 285456 271952 312912 271980
rect 285456 271940 285462 271952
rect 312906 271940 312912 271952
rect 312964 271940 312970 271992
rect 314286 271940 314292 271992
rect 314344 271980 314350 271992
rect 388622 271980 388628 271992
rect 314344 271952 388628 271980
rect 314344 271940 314350 271952
rect 388622 271940 388628 271952
rect 388680 271940 388686 271992
rect 395430 271940 395436 271992
rect 395488 271980 395494 271992
rect 604914 271980 604920 271992
rect 395488 271952 604920 271980
rect 395488 271940 395494 271952
rect 604914 271940 604920 271952
rect 604972 271940 604978 271992
rect 66990 271872 66996 271924
rect 67048 271912 67054 271924
rect 192478 271912 192484 271924
rect 67048 271884 192484 271912
rect 67048 271872 67054 271884
rect 192478 271872 192484 271884
rect 192536 271872 192542 271924
rect 242250 271912 242256 271924
rect 198706 271884 242256 271912
rect 65886 271804 65892 271856
rect 65944 271844 65950 271856
rect 192110 271844 192116 271856
rect 65944 271816 192116 271844
rect 65944 271804 65950 271816
rect 192110 271804 192116 271816
rect 192168 271804 192174 271856
rect 197170 271844 197176 271856
rect 194612 271816 197176 271844
rect 120258 271736 120264 271788
rect 120316 271776 120322 271788
rect 156782 271776 156788 271788
rect 120316 271748 156788 271776
rect 120316 271736 120322 271748
rect 156782 271736 156788 271748
rect 156840 271736 156846 271788
rect 156874 271736 156880 271788
rect 156932 271776 156938 271788
rect 177850 271776 177856 271788
rect 156932 271748 177856 271776
rect 156932 271736 156938 271748
rect 177850 271736 177856 271748
rect 177908 271736 177914 271788
rect 177942 271736 177948 271788
rect 178000 271776 178006 271788
rect 194502 271776 194508 271788
rect 178000 271748 194508 271776
rect 178000 271736 178006 271748
rect 194502 271736 194508 271748
rect 194560 271736 194566 271788
rect 130838 271668 130844 271720
rect 130896 271708 130902 271720
rect 194612 271708 194640 271816
rect 197170 271804 197176 271816
rect 197228 271804 197234 271856
rect 198274 271804 198280 271856
rect 198332 271844 198338 271856
rect 198706 271844 198734 271884
rect 242250 271872 242256 271884
rect 242308 271872 242314 271924
rect 244366 271872 244372 271924
rect 244424 271912 244430 271924
rect 259546 271912 259552 271924
rect 244424 271884 259552 271912
rect 244424 271872 244430 271884
rect 259546 271872 259552 271884
rect 259604 271872 259610 271924
rect 290274 271872 290280 271924
rect 290332 271912 290338 271924
rect 325970 271912 325976 271924
rect 290332 271884 325976 271912
rect 290332 271872 290338 271884
rect 325970 271872 325976 271884
rect 326028 271872 326034 271924
rect 326706 271872 326712 271924
rect 326764 271912 326770 271924
rect 402790 271912 402796 271924
rect 326764 271884 402796 271912
rect 326764 271872 326770 271884
rect 402790 271872 402796 271884
rect 402848 271872 402854 271924
rect 402882 271872 402888 271924
rect 402940 271912 402946 271924
rect 619082 271912 619088 271924
rect 402940 271884 619088 271912
rect 402940 271872 402946 271884
rect 619082 271872 619088 271884
rect 619140 271872 619146 271924
rect 240870 271844 240876 271856
rect 198332 271816 198734 271844
rect 208412 271816 240876 271844
rect 198332 271804 198338 271816
rect 130896 271680 194640 271708
rect 130896 271668 130902 271680
rect 194686 271668 194692 271720
rect 194744 271708 194750 271720
rect 208412 271708 208440 271816
rect 240870 271804 240876 271816
rect 240928 271804 240934 271856
rect 245562 271804 245568 271856
rect 245620 271844 245626 271856
rect 260006 271844 260012 271856
rect 245620 271816 260012 271844
rect 245620 271804 245626 271816
rect 260006 271804 260012 271816
rect 260064 271804 260070 271856
rect 289354 271804 289360 271856
rect 289412 271844 289418 271856
rect 323578 271844 323584 271856
rect 289412 271816 323584 271844
rect 289412 271804 289418 271816
rect 323578 271804 323584 271816
rect 323636 271804 323642 271856
rect 325602 271804 325608 271856
rect 325660 271844 325666 271856
rect 409874 271844 409880 271856
rect 325660 271816 409880 271844
rect 325660 271804 325666 271816
rect 409874 271804 409880 271816
rect 409932 271804 409938 271856
rect 411990 271804 411996 271856
rect 412048 271844 412054 271856
rect 633342 271844 633348 271856
rect 412048 271816 633348 271844
rect 412048 271804 412054 271816
rect 633342 271804 633348 271816
rect 633400 271804 633406 271856
rect 240778 271736 240784 271788
rect 240836 271776 240842 271788
rect 258258 271776 258264 271788
rect 240836 271748 258264 271776
rect 240836 271736 240842 271748
rect 258258 271736 258264 271748
rect 258316 271736 258322 271788
rect 262122 271736 262128 271788
rect 262180 271776 262186 271788
rect 266262 271776 266268 271788
rect 262180 271748 266268 271776
rect 262180 271736 262186 271748
rect 266262 271736 266268 271748
rect 266320 271736 266326 271788
rect 292482 271736 292488 271788
rect 292540 271776 292546 271788
rect 330662 271776 330668 271788
rect 292540 271748 330668 271776
rect 292540 271736 292546 271748
rect 330662 271736 330668 271748
rect 330720 271736 330726 271788
rect 349982 271736 349988 271788
rect 350040 271776 350046 271788
rect 484302 271776 484308 271788
rect 350040 271748 484308 271776
rect 350040 271736 350046 271748
rect 484302 271736 484308 271748
rect 484360 271736 484366 271788
rect 194744 271680 208440 271708
rect 194744 271668 194750 271680
rect 208486 271668 208492 271720
rect 208544 271708 208550 271720
rect 226334 271708 226340 271720
rect 208544 271680 226340 271708
rect 208544 271668 208550 271680
rect 226334 271668 226340 271680
rect 226392 271668 226398 271720
rect 229002 271668 229008 271720
rect 229060 271708 229066 271720
rect 253750 271708 253756 271720
rect 229060 271680 253756 271708
rect 229060 271668 229066 271680
rect 253750 271668 253756 271680
rect 253808 271668 253814 271720
rect 290734 271668 290740 271720
rect 290792 271708 290798 271720
rect 327074 271708 327080 271720
rect 290792 271680 327080 271708
rect 290792 271668 290798 271680
rect 327074 271668 327080 271680
rect 327132 271668 327138 271720
rect 336734 271668 336740 271720
rect 336792 271708 336798 271720
rect 343634 271708 343640 271720
rect 336792 271680 343640 271708
rect 336792 271668 336798 271680
rect 343634 271668 343640 271680
rect 343692 271668 343698 271720
rect 350902 271668 350908 271720
rect 350960 271708 350966 271720
rect 486694 271708 486700 271720
rect 350960 271680 486700 271708
rect 350960 271668 350966 271680
rect 486694 271668 486700 271680
rect 486752 271668 486758 271720
rect 165154 271600 165160 271652
rect 165212 271640 165218 271652
rect 229278 271640 229284 271652
rect 165212 271612 229284 271640
rect 165212 271600 165218 271612
rect 229278 271600 229284 271612
rect 229336 271600 229342 271652
rect 231394 271600 231400 271652
rect 231452 271640 231458 271652
rect 254670 271640 254676 271652
rect 231452 271612 254676 271640
rect 231452 271600 231458 271612
rect 254670 271600 254676 271612
rect 254728 271600 254734 271652
rect 289814 271600 289820 271652
rect 289872 271640 289878 271652
rect 324774 271640 324780 271652
rect 289872 271612 324780 271640
rect 289872 271600 289878 271612
rect 324774 271600 324780 271612
rect 324832 271600 324838 271652
rect 348234 271600 348240 271652
rect 348292 271640 348298 271652
rect 479610 271640 479616 271652
rect 348292 271612 479616 271640
rect 348292 271600 348298 271612
rect 479610 271600 479616 271612
rect 479668 271600 479674 271652
rect 163958 271532 163964 271584
rect 164016 271572 164022 271584
rect 229738 271572 229744 271584
rect 164016 271544 229744 271572
rect 164016 271532 164022 271544
rect 229738 271532 229744 271544
rect 229796 271532 229802 271584
rect 249058 271532 249064 271584
rect 249116 271572 249122 271584
rect 261386 271572 261392 271584
rect 249116 271544 261392 271572
rect 249116 271532 249122 271544
rect 261386 271532 261392 271544
rect 261444 271532 261450 271584
rect 291194 271532 291200 271584
rect 291252 271572 291258 271584
rect 328270 271572 328276 271584
rect 291252 271544 328276 271572
rect 291252 271532 291258 271544
rect 328270 271532 328276 271544
rect 328328 271532 328334 271584
rect 347590 271532 347596 271584
rect 347648 271572 347654 271584
rect 477218 271572 477224 271584
rect 347648 271544 477224 271572
rect 347648 271532 347654 271544
rect 477218 271532 477224 271544
rect 477276 271532 477282 271584
rect 158070 271464 158076 271516
rect 158128 271504 158134 271516
rect 177942 271504 177948 271516
rect 158128 271476 177948 271504
rect 158128 271464 158134 271476
rect 177942 271464 177948 271476
rect 178000 271464 178006 271516
rect 178126 271464 178132 271516
rect 178184 271504 178190 271516
rect 228818 271504 228824 271516
rect 178184 271476 228824 271504
rect 178184 271464 178190 271476
rect 228818 271464 228824 271476
rect 228876 271464 228882 271516
rect 252646 271464 252652 271516
rect 252704 271504 252710 271516
rect 262858 271504 262864 271516
rect 252704 271476 262864 271504
rect 252704 271464 252710 271476
rect 262858 271464 262864 271476
rect 262916 271464 262922 271516
rect 288986 271464 288992 271516
rect 289044 271504 289050 271516
rect 322382 271504 322388 271516
rect 289044 271476 322388 271504
rect 289044 271464 289050 271476
rect 322382 271464 322388 271476
rect 322440 271464 322446 271516
rect 342806 271464 342812 271516
rect 342864 271504 342870 271516
rect 465442 271504 465448 271516
rect 342864 271476 465448 271504
rect 342864 271464 342870 271476
rect 465442 271464 465448 271476
rect 465500 271464 465506 271516
rect 171042 271396 171048 271448
rect 171100 271436 171106 271448
rect 232406 271436 232412 271448
rect 171100 271408 232412 271436
rect 171100 271396 171106 271408
rect 232406 271396 232412 271408
rect 232464 271396 232470 271448
rect 258534 271396 258540 271448
rect 258592 271436 258598 271448
rect 264882 271436 264888 271448
rect 258592 271408 264888 271436
rect 258592 271396 258598 271408
rect 264882 271396 264888 271408
rect 264940 271396 264946 271448
rect 288526 271396 288532 271448
rect 288584 271436 288590 271448
rect 321186 271436 321192 271448
rect 288584 271408 321192 271436
rect 288584 271396 288590 271408
rect 321186 271396 321192 271408
rect 321244 271396 321250 271448
rect 354766 271396 354772 271448
rect 354824 271436 354830 271448
rect 472526 271436 472532 271448
rect 354824 271408 472532 271436
rect 354824 271396 354830 271408
rect 472526 271396 472532 271408
rect 472584 271396 472590 271448
rect 172238 271328 172244 271380
rect 172296 271368 172302 271380
rect 172296 271340 180012 271368
rect 172296 271328 172302 271340
rect 162762 271260 162768 271312
rect 162820 271300 162826 271312
rect 178126 271300 178132 271312
rect 162820 271272 178132 271300
rect 162820 271260 162826 271272
rect 178126 271260 178132 271272
rect 178184 271260 178190 271312
rect 179984 271300 180012 271340
rect 180058 271328 180064 271380
rect 180116 271368 180122 271380
rect 231486 271368 231492 271380
rect 180116 271340 231492 271368
rect 180116 271328 180122 271340
rect 231486 271328 231492 271340
rect 231544 271328 231550 271380
rect 256142 271328 256148 271380
rect 256200 271368 256206 271380
rect 264054 271368 264060 271380
rect 256200 271340 264060 271368
rect 256200 271328 256206 271340
rect 264054 271328 264060 271340
rect 264112 271328 264118 271380
rect 286594 271328 286600 271380
rect 286652 271368 286658 271380
rect 315298 271368 315304 271380
rect 286652 271340 315304 271368
rect 286652 271328 286658 271340
rect 315298 271328 315304 271340
rect 315356 271328 315362 271380
rect 340230 271328 340236 271380
rect 340288 271368 340294 271380
rect 458358 271368 458364 271380
rect 340288 271340 458364 271368
rect 340288 271328 340294 271340
rect 458358 271328 458364 271340
rect 458416 271328 458422 271380
rect 231762 271300 231768 271312
rect 179984 271272 231768 271300
rect 231762 271260 231768 271272
rect 231820 271260 231826 271312
rect 255038 271260 255044 271312
rect 255096 271300 255102 271312
rect 263594 271300 263600 271312
rect 255096 271272 263600 271300
rect 255096 271260 255102 271272
rect 263594 271260 263600 271272
rect 263652 271260 263658 271312
rect 287606 271260 287612 271312
rect 287664 271300 287670 271312
rect 318794 271300 318800 271312
rect 287664 271272 318800 271300
rect 287664 271260 287670 271272
rect 318794 271260 318800 271272
rect 318852 271260 318858 271312
rect 337470 271260 337476 271312
rect 337528 271300 337534 271312
rect 451274 271300 451280 271312
rect 337528 271272 451280 271300
rect 337528 271260 337534 271272
rect 451274 271260 451280 271272
rect 451332 271260 451338 271312
rect 178034 271192 178040 271244
rect 178092 271232 178098 271244
rect 189258 271232 189264 271244
rect 178092 271204 189264 271232
rect 178092 271192 178098 271204
rect 189258 271192 189264 271204
rect 189316 271192 189322 271244
rect 197262 271192 197268 271244
rect 197320 271232 197326 271244
rect 232682 271232 232688 271244
rect 197320 271204 232688 271232
rect 197320 271192 197326 271204
rect 232682 271192 232688 271204
rect 232740 271192 232746 271244
rect 251450 271192 251456 271244
rect 251508 271232 251514 271244
rect 262214 271232 262220 271244
rect 251508 271204 262220 271232
rect 251508 271192 251514 271204
rect 262214 271192 262220 271204
rect 262272 271192 262278 271244
rect 266814 271192 266820 271244
rect 266872 271232 266878 271244
rect 268010 271232 268016 271244
rect 266872 271204 268016 271232
rect 266872 271192 266878 271204
rect 268010 271192 268016 271204
rect 268068 271192 268074 271244
rect 287146 271192 287152 271244
rect 287204 271232 287210 271244
rect 317690 271232 317696 271244
rect 287204 271204 317696 271232
rect 287204 271192 287210 271204
rect 317690 271192 317696 271204
rect 317748 271192 317754 271244
rect 329742 271192 329748 271244
rect 329800 271232 329806 271244
rect 340138 271232 340144 271244
rect 329800 271204 340144 271232
rect 329800 271192 329806 271204
rect 340138 271192 340144 271204
rect 340196 271192 340202 271244
rect 448882 271232 448888 271244
rect 340248 271204 448888 271232
rect 179322 271124 179328 271176
rect 179380 271164 179386 271176
rect 234522 271164 234528 271176
rect 179380 271136 234528 271164
rect 179380 271124 179386 271136
rect 234522 271124 234528 271136
rect 234580 271124 234586 271176
rect 247862 271124 247868 271176
rect 247920 271164 247926 271176
rect 260926 271164 260932 271176
rect 247920 271136 260932 271164
rect 247920 271124 247926 271136
rect 260926 271124 260932 271136
rect 260984 271124 260990 271176
rect 286686 271124 286692 271176
rect 286744 271164 286750 271176
rect 316494 271164 316500 271176
rect 286744 271136 316500 271164
rect 286744 271124 286750 271136
rect 316494 271124 316500 271136
rect 316552 271124 316558 271176
rect 336642 271124 336648 271176
rect 336700 271164 336706 271176
rect 340248 271164 340276 271204
rect 448882 271192 448888 271204
rect 448940 271192 448946 271244
rect 415302 271164 415308 271176
rect 336700 271136 340276 271164
rect 340340 271136 415308 271164
rect 336700 271124 336706 271136
rect 169846 271056 169852 271108
rect 169904 271096 169910 271108
rect 180058 271096 180064 271108
rect 169904 271068 180064 271096
rect 169904 271056 169910 271068
rect 180058 271056 180064 271068
rect 180116 271056 180122 271108
rect 182910 271056 182916 271108
rect 182968 271096 182974 271108
rect 232958 271096 232964 271108
rect 182968 271068 232964 271096
rect 182968 271056 182974 271068
rect 232958 271056 232964 271068
rect 233016 271056 233022 271108
rect 253842 271056 253848 271108
rect 253900 271096 253906 271108
rect 263134 271096 263140 271108
rect 253900 271068 263140 271096
rect 253900 271056 253906 271068
rect 263134 271056 263140 271068
rect 263192 271056 263198 271108
rect 288158 271056 288164 271108
rect 288216 271096 288222 271108
rect 319990 271096 319996 271108
rect 288216 271068 319996 271096
rect 288216 271056 288222 271068
rect 319990 271056 319996 271068
rect 320048 271056 320054 271108
rect 334802 271056 334808 271108
rect 334860 271096 334866 271108
rect 340340 271096 340368 271136
rect 415302 271124 415308 271136
rect 415360 271124 415366 271176
rect 420914 271124 420920 271176
rect 420972 271164 420978 271176
rect 441798 271164 441804 271176
rect 420972 271136 441804 271164
rect 420972 271124 420978 271136
rect 441798 271124 441804 271136
rect 441856 271124 441862 271176
rect 420730 271096 420736 271108
rect 334860 271068 340368 271096
rect 340432 271068 420736 271096
rect 334860 271056 334866 271068
rect 176930 270988 176936 271040
rect 176988 271028 176994 271040
rect 227622 271028 227628 271040
rect 176988 271000 227628 271028
rect 176988 270988 176994 271000
rect 227622 270988 227628 271000
rect 227680 270988 227686 271040
rect 246758 270988 246764 271040
rect 246816 271028 246822 271040
rect 260466 271028 260472 271040
rect 246816 271000 260472 271028
rect 246816 270988 246822 271000
rect 260466 270988 260472 271000
rect 260524 270988 260530 271040
rect 285858 270988 285864 271040
rect 285916 271028 285922 271040
rect 314102 271028 314108 271040
rect 285916 271000 314108 271028
rect 285916 270988 285922 271000
rect 314102 270988 314108 271000
rect 314160 270988 314166 271040
rect 333974 270988 333980 271040
rect 334032 271028 334038 271040
rect 340432 271028 340460 271068
rect 420730 271056 420736 271068
rect 420788 271056 420794 271108
rect 444190 271096 444196 271108
rect 430546 271068 444196 271096
rect 334032 271000 340460 271028
rect 340524 271000 414152 271028
rect 334032 270988 334038 271000
rect 185210 270920 185216 270972
rect 185268 270960 185274 270972
rect 234706 270960 234712 270972
rect 185268 270932 234712 270960
rect 185268 270920 185274 270932
rect 234706 270920 234712 270932
rect 234764 270920 234770 270972
rect 250254 270920 250260 270972
rect 250312 270960 250318 270972
rect 261846 270960 261852 270972
rect 250312 270932 261852 270960
rect 250312 270920 250318 270932
rect 261846 270920 261852 270932
rect 261904 270920 261910 270972
rect 331306 270920 331312 270972
rect 331364 270960 331370 270972
rect 340524 270960 340552 271000
rect 331364 270932 340552 270960
rect 340616 270932 414060 270960
rect 331364 270920 331370 270932
rect 186406 270852 186412 270904
rect 186464 270892 186470 270904
rect 233418 270892 233424 270904
rect 186464 270864 233424 270892
rect 186464 270852 186470 270864
rect 233418 270852 233424 270864
rect 233476 270852 233482 270904
rect 329926 270852 329932 270904
rect 329984 270892 329990 270904
rect 340616 270892 340644 270932
rect 329984 270864 340644 270892
rect 340708 270864 413876 270892
rect 329984 270852 329990 270864
rect 175826 270784 175832 270836
rect 175884 270824 175890 270836
rect 179322 270824 179328 270836
rect 175884 270796 179328 270824
rect 175884 270784 175890 270796
rect 179322 270784 179328 270796
rect 179380 270784 179386 270836
rect 189994 270784 190000 270836
rect 190052 270824 190058 270836
rect 231854 270824 231860 270836
rect 190052 270796 231860 270824
rect 190052 270784 190058 270796
rect 231854 270784 231860 270796
rect 231912 270784 231918 270836
rect 259730 270784 259736 270836
rect 259788 270824 259794 270836
rect 265434 270824 265440 270836
rect 259788 270796 265440 270824
rect 259788 270784 259794 270796
rect 265434 270784 265440 270796
rect 265492 270784 265498 270836
rect 327258 270784 327264 270836
rect 327316 270824 327322 270836
rect 340708 270824 340736 270864
rect 327316 270796 340736 270824
rect 327316 270784 327322 270796
rect 340782 270784 340788 270836
rect 340840 270824 340846 270836
rect 340840 270796 411254 270824
rect 340840 270784 340846 270796
rect 187602 270716 187608 270768
rect 187660 270756 187666 270768
rect 230750 270756 230756 270768
rect 187660 270728 230756 270756
rect 187660 270716 187666 270728
rect 230750 270716 230756 270728
rect 230808 270716 230814 270768
rect 326430 270716 326436 270768
rect 326488 270756 326494 270768
rect 395706 270756 395712 270768
rect 326488 270728 395712 270756
rect 326488 270716 326494 270728
rect 395706 270716 395712 270728
rect 395764 270716 395770 270768
rect 191190 270648 191196 270700
rect 191248 270688 191254 270700
rect 229094 270688 229100 270700
rect 191248 270660 218054 270688
rect 191248 270648 191254 270660
rect 192294 270512 192300 270564
rect 192352 270552 192358 270564
rect 198642 270552 198648 270564
rect 192352 270524 198648 270552
rect 192352 270512 192358 270524
rect 198642 270512 198648 270524
rect 198700 270512 198706 270564
rect 218026 270552 218054 270660
rect 226536 270660 229100 270688
rect 226536 270552 226564 270660
rect 229094 270648 229100 270660
rect 229152 270648 229158 270700
rect 257338 270648 257344 270700
rect 257396 270688 257402 270700
rect 264514 270688 264520 270700
rect 257396 270660 264520 270688
rect 257396 270648 257402 270660
rect 264514 270648 264520 270660
rect 264572 270648 264578 270700
rect 331122 270648 331128 270700
rect 331180 270688 331186 270700
rect 377950 270688 377956 270700
rect 331180 270660 377956 270688
rect 331180 270648 331186 270660
rect 377950 270648 377956 270660
rect 378008 270648 378014 270700
rect 227806 270580 227812 270632
rect 227864 270620 227870 270632
rect 253382 270620 253388 270632
rect 227864 270592 253388 270620
rect 227864 270580 227870 270592
rect 253382 270580 253388 270592
rect 253440 270580 253446 270632
rect 324590 270580 324596 270632
rect 324648 270620 324654 270632
rect 340782 270620 340788 270632
rect 324648 270592 340788 270620
rect 324648 270580 324654 270592
rect 340782 270580 340788 270592
rect 340840 270580 340846 270632
rect 351730 270580 351736 270632
rect 351788 270620 351794 270632
rect 394510 270620 394516 270632
rect 351788 270592 394516 270620
rect 351788 270580 351794 270592
rect 394510 270580 394516 270592
rect 394568 270580 394574 270632
rect 411226 270620 411254 270796
rect 413848 270688 413876 270864
rect 414032 270824 414060 270932
rect 414124 270892 414152 271000
rect 415302 270988 415308 271040
rect 415360 271028 415366 271040
rect 430546 271028 430574 271068
rect 444190 271056 444196 271068
rect 444248 271056 444254 271108
rect 415360 271000 430574 271028
rect 415360 270988 415366 271000
rect 434714 270892 434720 270904
rect 414124 270864 434720 270892
rect 434714 270852 434720 270864
rect 434772 270852 434778 270904
rect 431126 270824 431132 270836
rect 414032 270796 431132 270824
rect 431126 270784 431132 270796
rect 431184 270784 431190 270836
rect 424042 270688 424048 270700
rect 413848 270660 424048 270688
rect 424042 270648 424048 270660
rect 424100 270648 424106 270700
rect 416958 270620 416964 270632
rect 411226 270592 416964 270620
rect 416958 270580 416964 270592
rect 417016 270580 417022 270632
rect 218026 270524 226564 270552
rect 226610 270512 226616 270564
rect 226668 270552 226674 270564
rect 252922 270552 252928 270564
rect 226668 270524 252928 270552
rect 226668 270512 226674 270524
rect 252922 270512 252928 270524
rect 252980 270512 252986 270564
rect 357434 270512 357440 270564
rect 357492 270552 357498 270564
rect 385034 270552 385040 270564
rect 357492 270524 385040 270552
rect 357492 270512 357498 270524
rect 385034 270512 385040 270524
rect 385092 270512 385098 270564
rect 411806 270512 411812 270564
rect 411864 270552 411870 270564
rect 413094 270552 413100 270564
rect 411864 270524 413100 270552
rect 411864 270512 411870 270524
rect 413094 270512 413100 270524
rect 413152 270512 413158 270564
rect 152182 270444 152188 270496
rect 152240 270484 152246 270496
rect 208026 270484 208032 270496
rect 152240 270456 208032 270484
rect 152240 270444 152246 270456
rect 208026 270444 208032 270456
rect 208084 270444 208090 270496
rect 220814 270484 220820 270496
rect 208228 270456 220820 270484
rect 147398 270376 147404 270428
rect 147456 270416 147462 270428
rect 208118 270416 208124 270428
rect 147456 270388 208124 270416
rect 147456 270376 147462 270388
rect 208118 270376 208124 270388
rect 208176 270376 208182 270428
rect 141510 270308 141516 270360
rect 141568 270348 141574 270360
rect 208228 270348 208256 270456
rect 220814 270444 220820 270456
rect 220872 270444 220878 270496
rect 225414 270444 225420 270496
rect 225472 270484 225478 270496
rect 252462 270484 252468 270496
rect 225472 270456 252468 270484
rect 225472 270444 225478 270456
rect 252462 270444 252468 270456
rect 252520 270444 252526 270496
rect 265618 270444 265624 270496
rect 265676 270484 265682 270496
rect 267550 270484 267556 270496
rect 265676 270456 267556 270484
rect 265676 270444 265682 270456
rect 267550 270444 267556 270456
rect 267608 270444 267614 270496
rect 269850 270444 269856 270496
rect 269908 270484 269914 270496
rect 271506 270484 271512 270496
rect 269908 270456 271512 270484
rect 269908 270444 269914 270456
rect 271506 270444 271512 270456
rect 271564 270444 271570 270496
rect 272058 270444 272064 270496
rect 272116 270484 272122 270496
rect 277486 270484 277492 270496
rect 272116 270456 277492 270484
rect 272116 270444 272122 270456
rect 277486 270444 277492 270456
rect 277544 270444 277550 270496
rect 304074 270444 304080 270496
rect 304132 270484 304138 270496
rect 344002 270484 344008 270496
rect 304132 270456 344008 270484
rect 304132 270444 304138 270456
rect 344002 270444 344008 270456
rect 344060 270444 344066 270496
rect 346854 270444 346860 270496
rect 346912 270484 346918 270496
rect 476114 270484 476120 270496
rect 346912 270456 476120 270484
rect 346912 270444 346918 270456
rect 476114 270444 476120 270456
rect 476172 270444 476178 270496
rect 219986 270416 219992 270428
rect 141568 270320 208256 270348
rect 208320 270388 219992 270416
rect 141568 270308 141574 270320
rect 140314 270240 140320 270292
rect 140372 270280 140378 270292
rect 208320 270280 208348 270388
rect 219986 270376 219992 270388
rect 220044 270376 220050 270428
rect 221918 270376 221924 270428
rect 221976 270416 221982 270428
rect 251082 270416 251088 270428
rect 221976 270388 251088 270416
rect 221976 270376 221982 270388
rect 251082 270376 251088 270388
rect 251140 270376 251146 270428
rect 270310 270376 270316 270428
rect 270368 270416 270374 270428
rect 272702 270416 272708 270428
rect 270368 270388 272708 270416
rect 270368 270376 270374 270388
rect 272702 270376 272708 270388
rect 272760 270376 272766 270428
rect 273714 270376 273720 270428
rect 273772 270416 273778 270428
rect 280982 270416 280988 270428
rect 273772 270388 280988 270416
rect 273772 270376 273778 270388
rect 280982 270376 280988 270388
rect 281040 270376 281046 270428
rect 294322 270376 294328 270428
rect 294380 270416 294386 270428
rect 336550 270416 336556 270428
rect 294380 270388 336556 270416
rect 294380 270376 294386 270388
rect 336550 270376 336556 270388
rect 336608 270376 336614 270428
rect 348602 270376 348608 270428
rect 348660 270416 348666 270428
rect 480806 270416 480812 270428
rect 348660 270388 480812 270416
rect 348660 270376 348666 270388
rect 480806 270376 480812 270388
rect 480864 270376 480870 270428
rect 219066 270348 219072 270360
rect 218026 270320 219072 270348
rect 218026 270280 218054 270320
rect 219066 270308 219072 270320
rect 219124 270308 219130 270360
rect 224218 270308 224224 270360
rect 224276 270348 224282 270360
rect 252002 270348 252008 270360
rect 224276 270320 252008 270348
rect 224276 270308 224282 270320
rect 252002 270308 252008 270320
rect 252060 270308 252066 270360
rect 271138 270308 271144 270360
rect 271196 270348 271202 270360
rect 275094 270348 275100 270360
rect 271196 270320 275100 270348
rect 271196 270308 271202 270320
rect 275094 270308 275100 270320
rect 275152 270308 275158 270360
rect 277394 270308 277400 270360
rect 277452 270348 277458 270360
rect 291654 270348 291660 270360
rect 277452 270320 291660 270348
rect 277452 270308 277458 270320
rect 291654 270308 291660 270320
rect 291712 270308 291718 270360
rect 296990 270308 296996 270360
rect 297048 270348 297054 270360
rect 336734 270348 336740 270360
rect 297048 270320 336740 270348
rect 297048 270308 297054 270320
rect 336734 270308 336740 270320
rect 336792 270308 336798 270360
rect 349522 270308 349528 270360
rect 349580 270348 349586 270360
rect 483198 270348 483204 270360
rect 349580 270320 483204 270348
rect 349580 270308 349586 270320
rect 483198 270308 483204 270320
rect 483256 270308 483262 270360
rect 140372 270252 208348 270280
rect 214760 270252 218054 270280
rect 140372 270240 140378 270252
rect 133230 270172 133236 270224
rect 133288 270212 133294 270224
rect 202506 270212 202512 270224
rect 133288 270184 202512 270212
rect 133288 270172 133294 270184
rect 202506 270172 202512 270184
rect 202564 270172 202570 270224
rect 202598 270172 202604 270224
rect 202656 270212 202662 270224
rect 214650 270212 214656 270224
rect 202656 270184 214656 270212
rect 202656 270172 202662 270184
rect 214650 270172 214656 270184
rect 214708 270172 214714 270224
rect 135622 270104 135628 270156
rect 135680 270144 135686 270156
rect 214760 270144 214788 270252
rect 219526 270240 219532 270292
rect 219584 270280 219590 270292
rect 250254 270280 250260 270292
rect 219584 270252 250260 270280
rect 219584 270240 219590 270252
rect 250254 270240 250260 270252
rect 250312 270240 250318 270292
rect 274266 270240 274272 270292
rect 274324 270280 274330 270292
rect 283374 270280 283380 270292
rect 274324 270252 283380 270280
rect 274324 270240 274330 270252
rect 283374 270240 283380 270252
rect 283432 270240 283438 270292
rect 283466 270240 283472 270292
rect 283524 270280 283530 270292
rect 290458 270280 290464 270292
rect 283524 270252 290464 270280
rect 283524 270240 283530 270252
rect 290458 270240 290464 270252
rect 290516 270240 290522 270292
rect 297450 270240 297456 270292
rect 297508 270280 297514 270292
rect 339494 270280 339500 270292
rect 297508 270252 339500 270280
rect 297508 270240 297514 270252
rect 339494 270240 339500 270252
rect 339552 270240 339558 270292
rect 351270 270240 351276 270292
rect 351328 270280 351334 270292
rect 487890 270280 487896 270292
rect 351328 270252 487896 270280
rect 351328 270240 351334 270252
rect 487890 270240 487896 270252
rect 487948 270240 487954 270292
rect 217134 270172 217140 270224
rect 217192 270212 217198 270224
rect 249334 270212 249340 270224
rect 217192 270184 249340 270212
rect 217192 270172 217198 270184
rect 249334 270172 249340 270184
rect 249392 270172 249398 270224
rect 277854 270172 277860 270224
rect 277912 270212 277918 270224
rect 292850 270212 292856 270224
rect 277912 270184 292856 270212
rect 277912 270172 277918 270184
rect 292850 270172 292856 270184
rect 292908 270172 292914 270224
rect 296530 270172 296536 270224
rect 296588 270212 296594 270224
rect 342438 270212 342444 270224
rect 296588 270184 342444 270212
rect 296588 270172 296594 270184
rect 342438 270172 342444 270184
rect 342496 270172 342502 270224
rect 352190 270172 352196 270224
rect 352248 270212 352254 270224
rect 490282 270212 490288 270224
rect 352248 270184 490288 270212
rect 352248 270172 352254 270184
rect 490282 270172 490288 270184
rect 490340 270172 490346 270224
rect 218146 270144 218152 270156
rect 135680 270116 214788 270144
rect 218026 270116 218152 270144
rect 135680 270104 135686 270116
rect 134426 270036 134432 270088
rect 134484 270076 134490 270088
rect 218026 270076 218054 270116
rect 218146 270104 218152 270116
rect 218204 270104 218210 270156
rect 223114 270104 223120 270156
rect 223172 270144 223178 270156
rect 251542 270144 251548 270156
rect 223172 270116 251548 270144
rect 223172 270104 223178 270116
rect 251542 270104 251548 270116
rect 251600 270104 251606 270156
rect 278590 270104 278596 270156
rect 278648 270144 278654 270156
rect 295150 270144 295156 270156
rect 278648 270116 295156 270144
rect 278648 270104 278654 270116
rect 295150 270104 295156 270116
rect 295208 270104 295214 270156
rect 298278 270104 298284 270156
rect 298336 270144 298342 270156
rect 347222 270144 347228 270156
rect 298336 270116 347228 270144
rect 298336 270104 298342 270116
rect 347222 270104 347228 270116
rect 347280 270104 347286 270156
rect 353570 270104 353576 270156
rect 353628 270144 353634 270156
rect 493778 270144 493784 270156
rect 353628 270116 493784 270144
rect 353628 270104 353634 270116
rect 493778 270104 493784 270116
rect 493836 270104 493842 270156
rect 134484 270048 218054 270076
rect 134484 270036 134490 270048
rect 220722 270036 220728 270088
rect 220780 270076 220786 270088
rect 250714 270076 250720 270088
rect 220780 270048 250720 270076
rect 220780 270036 220786 270048
rect 250714 270036 250720 270048
rect 250772 270036 250778 270088
rect 278314 270036 278320 270088
rect 278372 270076 278378 270088
rect 294046 270076 294052 270088
rect 278372 270048 294052 270076
rect 278372 270036 278378 270048
rect 294046 270036 294052 270048
rect 294104 270036 294110 270088
rect 299198 270036 299204 270088
rect 299256 270076 299262 270088
rect 349614 270076 349620 270088
rect 299256 270048 349620 270076
rect 299256 270036 299262 270048
rect 349614 270036 349620 270048
rect 349672 270036 349678 270088
rect 356238 270036 356244 270088
rect 356296 270076 356302 270088
rect 500862 270076 500868 270088
rect 356296 270048 500868 270076
rect 356296 270036 356302 270048
rect 500862 270036 500868 270048
rect 500920 270036 500926 270088
rect 126146 269968 126152 270020
rect 126204 270008 126210 270020
rect 202598 270008 202604 270020
rect 126204 269980 202604 270008
rect 126204 269968 126210 269980
rect 202598 269968 202604 269980
rect 202656 269968 202662 270020
rect 211890 270008 211896 270020
rect 202708 269980 211896 270008
rect 119062 269900 119068 269952
rect 119120 269940 119126 269952
rect 202708 269940 202736 269980
rect 211890 269968 211896 269980
rect 211948 269968 211954 270020
rect 215938 269968 215944 270020
rect 215996 270008 216002 270020
rect 248874 270008 248880 270020
rect 215996 269980 248880 270008
rect 215996 269968 216002 269980
rect 248874 269968 248880 269980
rect 248932 269968 248938 270020
rect 279142 269968 279148 270020
rect 279200 270008 279206 270020
rect 296346 270008 296352 270020
rect 279200 269980 296352 270008
rect 279200 269968 279206 269980
rect 296346 269968 296352 269980
rect 296404 269968 296410 270020
rect 345474 269968 345480 270020
rect 345532 270008 345538 270020
rect 354766 270008 354772 270020
rect 345532 269980 354772 270008
rect 345532 269968 345538 269980
rect 354766 269968 354772 269980
rect 354824 269968 354830 270020
rect 364702 269968 364708 270020
rect 364760 270008 364766 270020
rect 364760 269980 382412 270008
rect 364760 269968 364766 269980
rect 211062 269940 211068 269952
rect 119120 269912 202736 269940
rect 202800 269912 211068 269940
rect 119120 269900 119126 269912
rect 114278 269832 114284 269884
rect 114336 269872 114342 269884
rect 202800 269872 202828 269912
rect 211062 269900 211068 269912
rect 211120 269900 211126 269952
rect 214834 269900 214840 269952
rect 214892 269940 214898 269952
rect 248414 269940 248420 269952
rect 214892 269912 248420 269940
rect 214892 269900 214898 269912
rect 248414 269900 248420 269912
rect 248472 269900 248478 269952
rect 279602 269900 279608 269952
rect 279660 269940 279666 269952
rect 297542 269940 297548 269952
rect 279660 269912 297548 269940
rect 279660 269900 279666 269912
rect 297542 269900 297548 269912
rect 297600 269900 297606 269952
rect 305454 269900 305460 269952
rect 305512 269940 305518 269952
rect 366082 269940 366088 269952
rect 305512 269912 366088 269940
rect 305512 269900 305518 269912
rect 366082 269900 366088 269912
rect 366140 269900 366146 269952
rect 367370 269900 367376 269952
rect 367428 269940 367434 269952
rect 382384 269940 382412 269980
rect 382458 269968 382464 270020
rect 382516 270008 382522 270020
rect 515122 270008 515128 270020
rect 382516 269980 515128 270008
rect 382516 269968 382522 269980
rect 515122 269968 515128 269980
rect 515180 269968 515186 270020
rect 523402 269940 523408 269952
rect 367428 269912 382136 269940
rect 382384 269912 523408 269940
rect 367428 269900 367434 269912
rect 209682 269872 209688 269884
rect 114336 269844 202828 269872
rect 202892 269844 209688 269872
rect 114336 269832 114342 269844
rect 110782 269764 110788 269816
rect 110840 269804 110846 269816
rect 202892 269804 202920 269844
rect 209682 269832 209688 269844
rect 209740 269832 209746 269884
rect 210050 269832 210056 269884
rect 210108 269872 210114 269884
rect 246666 269872 246672 269884
rect 210108 269844 246672 269872
rect 210108 269832 210114 269844
rect 246666 269832 246672 269844
rect 246724 269832 246730 269884
rect 274726 269832 274732 269884
rect 274784 269872 274790 269884
rect 284570 269872 284576 269884
rect 274784 269844 284576 269872
rect 274784 269832 274790 269844
rect 284570 269832 284576 269844
rect 284628 269832 284634 269884
rect 306742 269832 306748 269884
rect 306800 269872 306806 269884
rect 369670 269872 369676 269884
rect 306800 269844 369676 269872
rect 306800 269832 306806 269844
rect 369670 269832 369676 269844
rect 369728 269832 369734 269884
rect 370038 269832 370044 269884
rect 370096 269872 370102 269884
rect 382108 269872 382136 269912
rect 523402 269900 523408 269912
rect 523460 269900 523466 269952
rect 530486 269872 530492 269884
rect 370096 269844 382044 269872
rect 382108 269844 530492 269872
rect 370096 269832 370102 269844
rect 110840 269776 202920 269804
rect 110840 269764 110846 269776
rect 202966 269764 202972 269816
rect 203024 269804 203030 269816
rect 208394 269804 208400 269816
rect 203024 269776 208400 269804
rect 203024 269764 203030 269776
rect 208394 269764 208400 269776
rect 208452 269764 208458 269816
rect 212442 269764 212448 269816
rect 212500 269804 212506 269816
rect 247586 269804 247592 269816
rect 212500 269776 247592 269804
rect 212500 269764 212506 269776
rect 247586 269764 247592 269776
rect 247644 269764 247650 269816
rect 280522 269764 280528 269816
rect 280580 269804 280586 269816
rect 299934 269804 299940 269816
rect 280580 269776 299940 269804
rect 280580 269764 280586 269776
rect 299934 269764 299940 269776
rect 299992 269764 299998 269816
rect 307202 269764 307208 269816
rect 307260 269804 307266 269816
rect 370866 269804 370872 269816
rect 307260 269776 370872 269804
rect 307260 269764 307266 269776
rect 370866 269764 370872 269776
rect 370924 269764 370930 269816
rect 373258 269804 373264 269816
rect 372586 269776 373264 269804
rect 109586 269696 109592 269748
rect 109644 269736 109650 269748
rect 109644 269708 206508 269736
rect 109644 269696 109650 269708
rect 95418 269628 95424 269680
rect 95476 269668 95482 269680
rect 203518 269668 203524 269680
rect 95476 269640 203524 269668
rect 95476 269628 95482 269640
rect 203518 269628 203524 269640
rect 203576 269628 203582 269680
rect 102502 269560 102508 269612
rect 102560 269600 102566 269612
rect 206186 269600 206192 269612
rect 102560 269572 206192 269600
rect 102560 269560 102566 269572
rect 206186 269560 206192 269572
rect 206244 269560 206250 269612
rect 206480 269600 206508 269708
rect 207750 269696 207756 269748
rect 207808 269736 207814 269748
rect 245746 269736 245752 269748
rect 207808 269708 245752 269736
rect 207808 269696 207814 269708
rect 245746 269696 245752 269708
rect 245804 269696 245810 269748
rect 280062 269696 280068 269748
rect 280120 269736 280126 269748
rect 298738 269736 298744 269748
rect 280120 269708 298744 269736
rect 280120 269696 280126 269708
rect 298738 269696 298744 269708
rect 298796 269696 298802 269748
rect 308122 269696 308128 269748
rect 308180 269736 308186 269748
rect 372586 269736 372614 269776
rect 373258 269764 373264 269776
rect 373316 269764 373322 269816
rect 382016 269804 382044 269844
rect 530486 269832 530492 269844
rect 530544 269832 530550 269884
rect 537570 269804 537576 269816
rect 382016 269776 537576 269804
rect 537570 269764 537576 269776
rect 537628 269764 537634 269816
rect 703556 269776 709012 269804
rect 703556 269748 703584 269776
rect 708984 269748 709012 269776
rect 308180 269708 372614 269736
rect 308180 269696 308186 269708
rect 375374 269696 375380 269748
rect 375432 269736 375438 269748
rect 375432 269708 382412 269736
rect 375432 269696 375438 269708
rect 206554 269628 206560 269680
rect 206612 269668 206618 269680
rect 224126 269668 224132 269680
rect 206612 269640 224132 269668
rect 206612 269628 206618 269640
rect 224126 269628 224132 269640
rect 224184 269628 224190 269680
rect 234614 269628 234620 269680
rect 234672 269668 234678 269680
rect 239122 269668 239128 269680
rect 234672 269640 239128 269668
rect 234672 269628 234678 269640
rect 239122 269628 239128 269640
rect 239180 269628 239186 269680
rect 281810 269628 281816 269680
rect 281868 269668 281874 269680
rect 303430 269668 303436 269680
rect 281868 269640 303436 269668
rect 281868 269628 281874 269640
rect 303430 269628 303436 269640
rect 303488 269628 303494 269680
rect 328638 269628 328644 269680
rect 328696 269668 328702 269680
rect 351914 269668 351920 269680
rect 328696 269640 351920 269668
rect 328696 269628 328702 269640
rect 351914 269628 351920 269640
rect 351972 269628 351978 269680
rect 361574 269628 361580 269680
rect 361632 269668 361638 269680
rect 382274 269668 382280 269680
rect 361632 269640 382280 269668
rect 361632 269628 361638 269640
rect 382274 269628 382280 269640
rect 382332 269628 382338 269680
rect 382384 269668 382412 269708
rect 382458 269696 382464 269748
rect 382516 269736 382522 269748
rect 544654 269736 544660 269748
rect 382516 269708 544660 269736
rect 382516 269696 382522 269708
rect 544654 269696 544660 269708
rect 544712 269696 544718 269748
rect 703538 269696 703544 269748
rect 703596 269696 703602 269748
rect 703998 269696 704004 269748
rect 704056 269736 704062 269748
rect 708874 269736 708880 269748
rect 704056 269708 708880 269736
rect 704056 269696 704062 269708
rect 708874 269696 708880 269708
rect 708932 269696 708938 269748
rect 708966 269696 708972 269748
rect 709024 269696 709030 269748
rect 551738 269668 551744 269680
rect 382384 269640 551744 269668
rect 551738 269628 551744 269640
rect 551796 269628 551802 269680
rect 708046 269668 708052 269680
rect 704844 269640 708052 269668
rect 208854 269600 208860 269612
rect 206480 269572 208860 269600
rect 208854 269560 208860 269572
rect 208912 269560 208918 269612
rect 209130 269560 209136 269612
rect 209188 269600 209194 269612
rect 246206 269600 246212 269612
rect 209188 269572 246212 269600
rect 209188 269560 209194 269572
rect 246206 269560 246212 269572
rect 246264 269560 246270 269612
rect 281442 269560 281448 269612
rect 281500 269600 281506 269612
rect 302326 269600 302332 269612
rect 281500 269572 302332 269600
rect 281500 269560 281506 269572
rect 302326 269560 302332 269572
rect 302384 269560 302390 269612
rect 310790 269560 310796 269612
rect 310848 269600 310854 269612
rect 380342 269600 380348 269612
rect 310848 269572 380348 269600
rect 310848 269560 310854 269572
rect 380342 269560 380348 269572
rect 380400 269560 380406 269612
rect 380710 269560 380716 269612
rect 380768 269600 380774 269612
rect 565906 269600 565912 269612
rect 380768 269572 565912 269600
rect 380768 269560 380774 269572
rect 565906 269560 565912 269572
rect 565964 269560 565970 269612
rect 704844 269544 704872 269640
rect 708046 269628 708052 269640
rect 708104 269628 708110 269680
rect 704918 269560 704924 269612
rect 704976 269600 704982 269612
rect 707954 269600 707960 269612
rect 704976 269572 707960 269600
rect 704976 269560 704982 269572
rect 707954 269560 707960 269572
rect 708012 269560 708018 269612
rect 94222 269492 94228 269544
rect 94280 269532 94286 269544
rect 202598 269532 202604 269544
rect 94280 269504 202604 269532
rect 94280 269492 94286 269504
rect 202598 269492 202604 269504
rect 202656 269492 202662 269544
rect 204162 269492 204168 269544
rect 204220 269532 204226 269544
rect 244458 269532 244464 269544
rect 204220 269504 244464 269532
rect 204220 269492 204226 269504
rect 244458 269492 244464 269504
rect 244516 269492 244522 269544
rect 280982 269492 280988 269544
rect 281040 269532 281046 269544
rect 301130 269532 301136 269544
rect 281040 269504 301136 269532
rect 281040 269492 281046 269504
rect 301130 269492 301136 269504
rect 301188 269492 301194 269544
rect 312078 269492 312084 269544
rect 312136 269532 312142 269544
rect 383838 269532 383844 269544
rect 312136 269504 383844 269532
rect 312136 269492 312142 269504
rect 383838 269492 383844 269504
rect 383896 269492 383902 269544
rect 386046 269492 386052 269544
rect 386104 269532 386110 269544
rect 580074 269532 580080 269544
rect 386104 269504 580080 269532
rect 386104 269492 386110 269504
rect 580074 269492 580080 269504
rect 580132 269492 580138 269544
rect 704826 269492 704832 269544
rect 704884 269492 704890 269544
rect 707034 269532 707040 269544
rect 705764 269504 707040 269532
rect 74074 269424 74080 269476
rect 74132 269464 74138 269476
rect 195882 269464 195888 269476
rect 74132 269436 195888 269464
rect 74132 269424 74138 269436
rect 195882 269424 195888 269436
rect 195940 269424 195946 269476
rect 198642 269424 198648 269476
rect 198700 269464 198706 269476
rect 198700 269436 208348 269464
rect 198700 269424 198706 269436
rect 80054 269356 80060 269408
rect 80112 269396 80118 269408
rect 197262 269396 197268 269408
rect 80112 269368 197268 269396
rect 80112 269356 80118 269368
rect 197262 269356 197268 269368
rect 197320 269356 197326 269408
rect 197354 269356 197360 269408
rect 197412 269396 197418 269408
rect 208320 269396 208348 269436
rect 208394 269424 208400 269476
rect 208452 269464 208458 269476
rect 243998 269464 244004 269476
rect 208452 269436 244004 269464
rect 208452 269424 208458 269436
rect 243998 269424 244004 269436
rect 244056 269424 244062 269476
rect 282730 269424 282736 269476
rect 282788 269464 282794 269476
rect 305822 269464 305828 269476
rect 282788 269436 305828 269464
rect 282788 269424 282794 269436
rect 305822 269424 305828 269436
rect 305880 269424 305886 269476
rect 313458 269424 313464 269476
rect 313516 269464 313522 269476
rect 387426 269464 387432 269476
rect 313516 269436 387432 269464
rect 313516 269424 313522 269436
rect 387426 269424 387432 269436
rect 387484 269424 387490 269476
rect 388714 269424 388720 269476
rect 388772 269464 388778 269476
rect 587158 269464 587164 269476
rect 388772 269436 587164 269464
rect 388772 269424 388778 269436
rect 587158 269424 587164 269436
rect 587216 269424 587222 269476
rect 705764 269408 705792 269504
rect 707034 269492 707040 269504
rect 707092 269492 707098 269544
rect 706666 269464 706672 269476
rect 706224 269436 706672 269464
rect 706224 269408 706252 269436
rect 706666 269424 706672 269436
rect 706724 269424 706730 269476
rect 239950 269396 239956 269408
rect 197412 269368 198734 269396
rect 208320 269368 239956 269396
rect 197412 269356 197418 269368
rect 82354 269288 82360 269340
rect 82412 269328 82418 269340
rect 198550 269328 198556 269340
rect 82412 269300 198556 269328
rect 82412 269288 82418 269300
rect 198550 269288 198556 269300
rect 198608 269288 198614 269340
rect 198706 269328 198734 269368
rect 239950 269356 239956 269368
rect 240008 269356 240014 269408
rect 282270 269356 282276 269408
rect 282328 269396 282334 269408
rect 304626 269396 304632 269408
rect 282328 269368 304632 269396
rect 282328 269356 282334 269368
rect 304626 269356 304632 269368
rect 304684 269356 304690 269408
rect 314838 269356 314844 269408
rect 314896 269396 314902 269408
rect 390922 269396 390928 269408
rect 314896 269368 390928 269396
rect 314896 269356 314902 269368
rect 390922 269356 390928 269368
rect 390980 269356 390986 269408
rect 394050 269356 394056 269408
rect 394108 269396 394114 269408
rect 601418 269396 601424 269408
rect 394108 269368 601424 269396
rect 394108 269356 394114 269368
rect 601418 269356 601424 269368
rect 601476 269356 601482 269408
rect 705746 269356 705752 269408
rect 705804 269356 705810 269408
rect 706206 269356 706212 269408
rect 706264 269356 706270 269408
rect 706298 269356 706304 269408
rect 706356 269396 706362 269408
rect 706574 269396 706580 269408
rect 706356 269368 706580 269396
rect 706356 269356 706362 269368
rect 706574 269356 706580 269368
rect 706632 269356 706638 269408
rect 241790 269328 241796 269340
rect 198706 269300 241796 269328
rect 241790 269288 241796 269300
rect 241848 269288 241854 269340
rect 276934 269288 276940 269340
rect 276992 269328 276998 269340
rect 283466 269328 283472 269340
rect 276992 269300 283472 269328
rect 276992 269288 276998 269300
rect 283466 269288 283472 269300
rect 283524 269288 283530 269340
rect 283650 269288 283656 269340
rect 283708 269328 283714 269340
rect 308214 269328 308220 269340
rect 283708 269300 308220 269328
rect 283708 269288 283714 269300
rect 308214 269288 308220 269300
rect 308272 269288 308278 269340
rect 315206 269288 315212 269340
rect 315264 269328 315270 269340
rect 392118 269328 392124 269340
rect 315264 269300 392124 269328
rect 315264 269288 315270 269300
rect 392118 269288 392124 269300
rect 392176 269288 392182 269340
rect 396718 269288 396724 269340
rect 396776 269328 396782 269340
rect 608502 269328 608508 269340
rect 396776 269300 608508 269328
rect 396776 269288 396782 269300
rect 608502 269288 608508 269300
rect 608560 269288 608566 269340
rect 705838 269288 705844 269340
rect 705896 269328 705902 269340
rect 707034 269328 707040 269340
rect 705896 269300 707040 269328
rect 705896 269288 705902 269300
rect 707034 269288 707040 269300
rect 707092 269288 707098 269340
rect 707586 269288 707592 269340
rect 707644 269288 707650 269340
rect 81250 269220 81256 269272
rect 81308 269260 81314 269272
rect 198090 269260 198096 269272
rect 81308 269232 198096 269260
rect 81308 269220 81314 269232
rect 198090 269220 198096 269232
rect 198148 269220 198154 269272
rect 200574 269220 200580 269272
rect 200632 269260 200638 269272
rect 243078 269260 243084 269272
rect 200632 269232 243084 269260
rect 200632 269220 200638 269232
rect 243078 269220 243084 269232
rect 243136 269220 243142 269272
rect 283190 269220 283196 269272
rect 283248 269260 283254 269272
rect 307018 269260 307024 269272
rect 283248 269232 307024 269260
rect 283248 269220 283254 269232
rect 307018 269220 307024 269232
rect 307076 269220 307082 269272
rect 317874 269220 317880 269272
rect 317932 269260 317938 269272
rect 399202 269260 399208 269272
rect 317932 269232 399208 269260
rect 317932 269220 317938 269232
rect 399202 269220 399208 269232
rect 399260 269220 399266 269272
rect 399386 269220 399392 269272
rect 399444 269260 399450 269272
rect 615586 269260 615592 269272
rect 399444 269232 615592 269260
rect 399444 269220 399450 269232
rect 615586 269220 615592 269232
rect 615644 269220 615650 269272
rect 705378 269220 705384 269272
rect 705436 269260 705442 269272
rect 707494 269260 707500 269272
rect 705436 269232 707500 269260
rect 705436 269220 705442 269232
rect 707494 269220 707500 269232
rect 707552 269220 707558 269272
rect 71774 269152 71780 269204
rect 71832 269192 71838 269204
rect 194594 269192 194600 269204
rect 71832 269164 194600 269192
rect 71832 269152 71838 269164
rect 194594 269152 194600 269164
rect 194652 269152 194658 269204
rect 195790 269152 195796 269204
rect 195848 269192 195854 269204
rect 241330 269192 241336 269204
rect 195848 269164 241336 269192
rect 195848 269152 195854 269164
rect 241330 269152 241336 269164
rect 241388 269152 241394 269204
rect 284938 269152 284944 269204
rect 284996 269192 285002 269204
rect 311710 269192 311716 269204
rect 284996 269164 311716 269192
rect 284996 269152 285002 269164
rect 311710 269152 311716 269164
rect 311768 269152 311774 269204
rect 320542 269152 320548 269204
rect 320600 269192 320606 269204
rect 406286 269192 406292 269204
rect 320600 269164 406292 269192
rect 320600 269152 320606 269164
rect 406286 269152 406292 269164
rect 406344 269152 406350 269204
rect 411438 269152 411444 269204
rect 411496 269192 411502 269204
rect 647510 269192 647516 269204
rect 411496 269164 647516 269192
rect 411496 269152 411502 269164
rect 647510 269152 647516 269164
rect 647568 269152 647574 269204
rect 705286 269152 705292 269204
rect 705344 269192 705350 269204
rect 707604 269192 707632 269288
rect 705344 269164 707632 269192
rect 705344 269152 705350 269164
rect 708506 269152 708512 269204
rect 708564 269152 708570 269204
rect 193490 269084 193496 269136
rect 193548 269124 193554 269136
rect 240410 269124 240416 269136
rect 193548 269096 240416 269124
rect 193548 269084 193554 269096
rect 240410 269084 240416 269096
rect 240468 269084 240474 269136
rect 269390 269084 269396 269136
rect 269448 269124 269454 269136
rect 270402 269124 270408 269136
rect 269448 269096 270408 269124
rect 269448 269084 269454 269096
rect 270402 269084 270408 269096
rect 270460 269084 270466 269136
rect 284478 269084 284484 269136
rect 284536 269124 284542 269136
rect 310514 269124 310520 269136
rect 284536 269096 310520 269124
rect 284536 269084 284542 269096
rect 310514 269084 310520 269096
rect 310572 269084 310578 269136
rect 323210 269084 323216 269136
rect 323268 269124 323274 269136
rect 411806 269124 411812 269136
rect 323268 269096 411812 269124
rect 323268 269084 323274 269096
rect 411806 269084 411812 269096
rect 411864 269084 411870 269136
rect 411898 269084 411904 269136
rect 411956 269124 411962 269136
rect 648706 269124 648712 269136
rect 411956 269096 648712 269124
rect 411956 269084 411962 269096
rect 648706 269084 648712 269096
rect 648764 269084 648770 269136
rect 704458 269084 704464 269136
rect 704516 269124 704522 269136
rect 708414 269124 708420 269136
rect 704516 269096 708420 269124
rect 704516 269084 704522 269096
rect 708414 269084 708420 269096
rect 708472 269084 708478 269136
rect 154482 269016 154488 269068
rect 154540 269056 154546 269068
rect 225322 269056 225328 269068
rect 154540 269028 225328 269056
rect 154540 269016 154546 269028
rect 225322 269016 225328 269028
rect 225380 269016 225386 269068
rect 292942 269016 292948 269068
rect 293000 269056 293006 269068
rect 333054 269056 333060 269068
rect 293000 269028 333060 269056
rect 293000 269016 293006 269028
rect 333054 269016 333060 269028
rect 333112 269016 333118 269068
rect 351822 269056 351828 269068
rect 342226 269028 351828 269056
rect 159266 268948 159272 269000
rect 159324 268988 159330 269000
rect 224034 268988 224040 269000
rect 159324 268960 224040 268988
rect 159324 268948 159330 268960
rect 224034 268948 224040 268960
rect 224092 268948 224098 269000
rect 224126 268948 224132 269000
rect 224184 268988 224190 269000
rect 245286 268988 245292 269000
rect 224184 268960 245292 268988
rect 224184 268948 224190 268960
rect 245286 268948 245292 268960
rect 245344 268948 245350 269000
rect 295610 268948 295616 269000
rect 295668 268988 295674 269000
rect 329742 268988 329748 269000
rect 295668 268960 329748 268988
rect 295668 268948 295674 268960
rect 329742 268948 329748 268960
rect 329800 268948 329806 269000
rect 330846 268948 330852 269000
rect 330904 268988 330910 269000
rect 342226 268988 342254 269028
rect 351822 269016 351828 269028
rect 351880 269016 351886 269068
rect 473722 269056 473728 269068
rect 351932 269028 473728 269056
rect 330904 268960 342254 268988
rect 330904 268948 330910 268960
rect 345934 268948 345940 269000
rect 345992 268988 345998 269000
rect 351932 268988 351960 269028
rect 473722 269016 473728 269028
rect 473780 269016 473786 269068
rect 704366 269016 704372 269068
rect 704424 269056 704430 269068
rect 708524 269056 708552 269152
rect 704424 269028 708552 269056
rect 704424 269016 704430 269028
rect 345992 268960 351960 268988
rect 345992 268948 345998 268960
rect 352006 268948 352012 269000
rect 352064 268988 352070 269000
rect 466638 268988 466644 269000
rect 352064 268960 466644 268988
rect 352064 268948 352070 268960
rect 466638 268948 466644 268960
rect 466696 268948 466702 269000
rect 160462 268880 160468 268932
rect 160520 268920 160526 268932
rect 160520 268892 224080 268920
rect 160520 268880 160526 268892
rect 161566 268812 161572 268864
rect 161624 268852 161630 268864
rect 223758 268852 223764 268864
rect 161624 268824 223764 268852
rect 161624 268812 161630 268824
rect 223758 268812 223764 268824
rect 223816 268812 223822 268864
rect 224052 268852 224080 268892
rect 231854 268880 231860 268932
rect 231912 268920 231918 268932
rect 238662 268920 238668 268932
rect 231912 268892 238668 268920
rect 231912 268880 231918 268892
rect 238662 268880 238668 268892
rect 238720 268880 238726 268932
rect 309870 268880 309876 268932
rect 309928 268920 309934 268932
rect 331122 268920 331128 268932
rect 309928 268892 331128 268920
rect 309928 268880 309934 268892
rect 331122 268880 331128 268892
rect 331180 268880 331186 268932
rect 344186 268880 344192 268932
rect 344244 268920 344250 268932
rect 468938 268920 468944 268932
rect 344244 268892 468944 268920
rect 344244 268880 344250 268892
rect 468938 268880 468944 268892
rect 468996 268880 469002 268932
rect 228450 268852 228456 268864
rect 224052 268824 228456 268852
rect 228450 268812 228456 268824
rect 228508 268812 228514 268864
rect 229094 268812 229100 268864
rect 229152 268852 229158 268864
rect 239582 268852 239588 268864
rect 229152 268824 239588 268852
rect 229152 268812 229158 268824
rect 239582 268812 239588 268824
rect 239640 268812 239646 268864
rect 272978 268812 272984 268864
rect 273036 268852 273042 268864
rect 279786 268852 279792 268864
rect 273036 268824 279792 268852
rect 273036 268812 273042 268824
rect 279786 268812 279792 268824
rect 279844 268812 279850 268864
rect 341518 268812 341524 268864
rect 341576 268852 341582 268864
rect 461854 268852 461860 268864
rect 341576 268824 461860 268852
rect 341576 268812 341582 268824
rect 461854 268812 461860 268824
rect 461912 268812 461918 268864
rect 166350 268744 166356 268796
rect 166408 268784 166414 268796
rect 166408 268756 223804 268784
rect 166408 268744 166414 268756
rect 167546 268676 167552 268728
rect 167604 268716 167610 268728
rect 223776 268716 223804 268756
rect 224034 268744 224040 268796
rect 224092 268784 224098 268796
rect 227530 268784 227536 268796
rect 224092 268756 227536 268784
rect 224092 268744 224098 268756
rect 227530 268744 227536 268756
rect 227588 268744 227594 268796
rect 340598 268744 340604 268796
rect 340656 268784 340662 268796
rect 459554 268784 459560 268796
rect 340656 268756 459560 268784
rect 340656 268744 340662 268756
rect 459554 268744 459560 268756
rect 459612 268744 459618 268796
rect 230198 268716 230204 268728
rect 167604 268688 223712 268716
rect 223776 268688 230204 268716
rect 167604 268676 167610 268688
rect 173434 268608 173440 268660
rect 173492 268648 173498 268660
rect 223574 268648 223580 268660
rect 173492 268620 223580 268648
rect 173492 268608 173498 268620
rect 223574 268608 223580 268620
rect 223632 268608 223638 268660
rect 223684 268648 223712 268688
rect 230198 268676 230204 268688
rect 230256 268676 230262 268728
rect 273806 268676 273812 268728
rect 273864 268716 273870 268728
rect 282178 268716 282184 268728
rect 273864 268688 282184 268716
rect 273864 268676 273870 268688
rect 282178 268676 282184 268688
rect 282236 268676 282242 268728
rect 338850 268676 338856 268728
rect 338908 268716 338914 268728
rect 454770 268716 454776 268728
rect 338908 268688 454776 268716
rect 338908 268676 338914 268688
rect 454770 268676 454776 268688
rect 454828 268676 454834 268728
rect 231118 268648 231124 268660
rect 223684 268620 231124 268648
rect 231118 268608 231124 268620
rect 231176 268608 231182 268660
rect 337930 268608 337936 268660
rect 337988 268648 337994 268660
rect 452470 268648 452476 268660
rect 337988 268620 452476 268648
rect 337988 268608 337994 268620
rect 452470 268608 452476 268620
rect 452528 268608 452534 268660
rect 168650 268540 168656 268592
rect 168708 268580 168714 268592
rect 230658 268580 230664 268592
rect 168708 268552 230664 268580
rect 168708 268540 168714 268552
rect 230658 268540 230664 268552
rect 230716 268540 230722 268592
rect 230750 268540 230756 268592
rect 230808 268580 230814 268592
rect 236638 268580 236644 268592
rect 230808 268552 236644 268580
rect 230808 268540 230814 268552
rect 236638 268540 236644 268552
rect 236696 268540 236702 268592
rect 240134 268540 240140 268592
rect 240192 268580 240198 268592
rect 244918 268580 244924 268592
rect 240192 268552 244924 268580
rect 240192 268540 240198 268552
rect 244918 268540 244924 268552
rect 244976 268540 244982 268592
rect 336182 268540 336188 268592
rect 336240 268580 336246 268592
rect 447686 268580 447692 268592
rect 336240 268552 447692 268580
rect 336240 268540 336246 268552
rect 447686 268540 447692 268552
rect 447744 268540 447750 268592
rect 156782 268472 156788 268524
rect 156840 268512 156846 268524
rect 212810 268512 212816 268524
rect 156840 268484 212816 268512
rect 156840 268472 156846 268484
rect 212810 268472 212816 268484
rect 212868 268472 212874 268524
rect 213638 268472 213644 268524
rect 213696 268512 213702 268524
rect 248046 268512 248052 268524
rect 213696 268484 248052 268512
rect 213696 268472 213702 268484
rect 248046 268472 248052 268484
rect 248104 268472 248110 268524
rect 335262 268472 335268 268524
rect 335320 268512 335326 268524
rect 445294 268512 445300 268524
rect 335320 268484 445300 268512
rect 335320 268472 335326 268484
rect 445294 268472 445300 268484
rect 445352 268472 445358 268524
rect 174630 268404 174636 268456
rect 174688 268444 174694 268456
rect 233786 268444 233792 268456
rect 174688 268416 233792 268444
rect 174688 268404 174694 268416
rect 233786 268404 233792 268416
rect 233844 268404 233850 268456
rect 272518 268404 272524 268456
rect 272576 268444 272582 268456
rect 278682 268444 278688 268456
rect 272576 268416 278688 268444
rect 272576 268404 272582 268416
rect 278682 268404 278688 268416
rect 278740 268404 278746 268456
rect 325970 268404 325976 268456
rect 326028 268444 326034 268456
rect 332778 268444 332784 268456
rect 326028 268416 332784 268444
rect 326028 268404 326034 268416
rect 332778 268404 332784 268416
rect 332836 268404 332842 268456
rect 333514 268404 333520 268456
rect 333572 268444 333578 268456
rect 440602 268444 440608 268456
rect 333572 268416 440608 268444
rect 333572 268404 333578 268416
rect 440602 268404 440608 268416
rect 440660 268404 440666 268456
rect 179322 268336 179328 268388
rect 179380 268376 179386 268388
rect 233326 268376 233332 268388
rect 179380 268348 233332 268376
rect 179380 268336 179386 268348
rect 233326 268336 233332 268348
rect 233384 268336 233390 268388
rect 233418 268336 233424 268388
rect 233476 268376 233482 268388
rect 237282 268376 237288 268388
rect 233476 268348 237288 268376
rect 233476 268336 233482 268348
rect 237282 268336 237288 268348
rect 237340 268336 237346 268388
rect 309410 268336 309416 268388
rect 309468 268376 309474 268388
rect 332502 268376 332508 268388
rect 309468 268348 332508 268376
rect 309468 268336 309474 268348
rect 332502 268336 332508 268348
rect 332560 268336 332566 268388
rect 332594 268336 332600 268388
rect 332652 268376 332658 268388
rect 438210 268376 438216 268388
rect 332652 268348 438216 268376
rect 332652 268336 332658 268348
rect 438210 268336 438216 268348
rect 438268 268336 438274 268388
rect 181714 268268 181720 268320
rect 181772 268308 181778 268320
rect 223574 268308 223580 268320
rect 181772 268280 223580 268308
rect 181772 268268 181778 268280
rect 223574 268268 223580 268280
rect 223632 268268 223638 268320
rect 223666 268268 223672 268320
rect 223724 268308 223730 268320
rect 232866 268308 232872 268320
rect 223724 268280 232872 268308
rect 223724 268268 223730 268280
rect 232866 268268 232872 268280
rect 232924 268268 232930 268320
rect 232958 268268 232964 268320
rect 233016 268308 233022 268320
rect 235994 268308 236000 268320
rect 233016 268280 236000 268308
rect 233016 268268 233022 268280
rect 235994 268268 236000 268280
rect 236052 268268 236058 268320
rect 275186 268268 275192 268320
rect 275244 268308 275250 268320
rect 285766 268308 285772 268320
rect 275244 268280 285772 268308
rect 275244 268268 275250 268280
rect 285766 268268 285772 268280
rect 285824 268268 285830 268320
rect 312538 268268 312544 268320
rect 312596 268308 312602 268320
rect 312596 268280 332640 268308
rect 312596 268268 312602 268280
rect 180518 268200 180524 268252
rect 180576 268240 180582 268252
rect 235534 268240 235540 268252
rect 180576 268212 235540 268240
rect 180576 268200 180582 268212
rect 235534 268200 235540 268212
rect 235592 268200 235598 268252
rect 270678 268200 270684 268252
rect 270736 268240 270742 268252
rect 273898 268240 273904 268252
rect 270736 268212 273904 268240
rect 270736 268200 270742 268212
rect 273898 268200 273904 268212
rect 273956 268200 273962 268252
rect 275646 268200 275652 268252
rect 275704 268240 275710 268252
rect 286870 268240 286876 268252
rect 275704 268212 286876 268240
rect 275704 268200 275710 268212
rect 286870 268200 286876 268212
rect 286928 268200 286934 268252
rect 316126 268200 316132 268252
rect 316184 268240 316190 268252
rect 316184 268212 332364 268240
rect 316184 268200 316190 268212
rect 184106 268132 184112 268184
rect 184164 268172 184170 268184
rect 236914 268172 236920 268184
rect 184164 268144 236920 268172
rect 184164 268132 184170 268144
rect 236914 268132 236920 268144
rect 236972 268132 236978 268184
rect 316586 268132 316592 268184
rect 316644 268172 316650 268184
rect 326430 268172 326436 268184
rect 316644 268144 326436 268172
rect 316644 268132 316650 268144
rect 326430 268132 326436 268144
rect 326488 268132 326494 268184
rect 197170 268064 197176 268116
rect 197228 268104 197234 268116
rect 216858 268104 216864 268116
rect 197228 268076 216864 268104
rect 197228 268064 197234 268076
rect 216858 268064 216864 268076
rect 216916 268064 216922 268116
rect 218330 268064 218336 268116
rect 218388 268104 218394 268116
rect 218388 268076 222792 268104
rect 218388 268064 218394 268076
rect 189258 267996 189264 268048
rect 189316 268036 189322 268048
rect 200758 268036 200764 268048
rect 189316 268008 200764 268036
rect 189316 267996 189322 268008
rect 200758 267996 200764 268008
rect 200816 267996 200822 268048
rect 201310 267996 201316 268048
rect 201368 268036 201374 268048
rect 203886 268036 203892 268048
rect 201368 268008 203892 268036
rect 201368 267996 201374 268008
rect 203886 267996 203892 268008
rect 203944 267996 203950 268048
rect 208118 267996 208124 268048
rect 208176 268036 208182 268048
rect 222654 268036 222660 268048
rect 208176 268008 222660 268036
rect 208176 267996 208182 268008
rect 222654 267996 222660 268008
rect 222712 267996 222718 268048
rect 222764 268036 222792 268076
rect 223574 268064 223580 268116
rect 223632 268104 223638 268116
rect 236454 268104 236460 268116
rect 223632 268076 236460 268104
rect 223632 268064 223638 268076
rect 236454 268064 236460 268076
rect 236512 268064 236518 268116
rect 249794 268104 249800 268116
rect 236564 268076 249800 268104
rect 236564 268036 236592 268076
rect 249794 268064 249800 268076
rect 249852 268064 249858 268116
rect 222764 268008 236592 268036
rect 236638 267996 236644 268048
rect 236696 268036 236702 268048
rect 238202 268036 238208 268048
rect 236696 268008 238208 268036
rect 236696 267996 236702 268008
rect 238202 267996 238208 268008
rect 238260 267996 238266 268048
rect 271598 267996 271604 268048
rect 271656 268036 271662 268048
rect 276290 268036 276296 268048
rect 271656 268008 276296 268036
rect 271656 267996 271662 268008
rect 276290 267996 276296 268008
rect 276348 267996 276354 268048
rect 276382 267996 276388 268048
rect 276440 268036 276446 268048
rect 288066 268036 288072 268048
rect 276440 268008 288072 268036
rect 276440 267996 276446 268008
rect 288066 267996 288072 268008
rect 288124 267996 288130 268048
rect 298738 267996 298744 268048
rect 298796 268036 298802 268048
rect 307846 268036 307852 268048
rect 298796 268008 307852 268036
rect 298796 267996 298802 268008
rect 307846 267996 307852 268008
rect 307904 267996 307910 268048
rect 319254 267996 319260 268048
rect 319312 268036 319318 268048
rect 326706 268036 326712 268048
rect 319312 268008 326712 268036
rect 319312 267996 319318 268008
rect 326706 267996 326712 268008
rect 326764 267996 326770 268048
rect 88334 267928 88340 267980
rect 88392 267968 88398 267980
rect 201218 267968 201224 267980
rect 88392 267940 201224 267968
rect 88392 267928 88398 267940
rect 201218 267928 201224 267940
rect 201276 267928 201282 267980
rect 211246 267928 211252 267980
rect 211304 267968 211310 267980
rect 247126 267968 247132 267980
rect 211304 267940 235212 267968
rect 211304 267928 211310 267940
rect 208026 267860 208032 267912
rect 208084 267900 208090 267912
rect 224862 267900 224868 267912
rect 208084 267872 224868 267900
rect 208084 267860 208090 267872
rect 224862 267860 224868 267872
rect 224920 267860 224926 267912
rect 202506 267792 202512 267844
rect 202564 267832 202570 267844
rect 217318 267832 217324 267844
rect 202564 267804 217324 267832
rect 202564 267792 202570 267804
rect 217318 267792 217324 267804
rect 217376 267792 217382 267844
rect 223758 267792 223764 267844
rect 223816 267832 223822 267844
rect 227990 267832 227996 267844
rect 223816 267804 227996 267832
rect 223816 267792 223822 267804
rect 227990 267792 227996 267804
rect 228048 267792 228054 267844
rect 232682 267792 232688 267844
rect 232740 267832 232746 267844
rect 235074 267832 235080 267844
rect 232740 267804 235080 267832
rect 232740 267792 232746 267804
rect 235074 267792 235080 267804
rect 235132 267792 235138 267844
rect 235184 267832 235212 267940
rect 237346 267940 247132 267968
rect 237346 267832 237374 267940
rect 247126 267928 247132 267940
rect 247184 267928 247190 267980
rect 297910 267928 297916 267980
rect 297968 267968 297974 267980
rect 304902 267968 304908 267980
rect 297968 267940 304908 267968
rect 297968 267928 297974 267940
rect 304902 267928 304908 267940
rect 304960 267928 304966 267980
rect 321922 267928 321928 267980
rect 321980 267968 321986 267980
rect 325602 267968 325608 267980
rect 321980 267940 325608 267968
rect 321980 267928 321986 267940
rect 325602 267928 325608 267940
rect 325660 267928 325666 267980
rect 332336 267968 332364 268212
rect 332612 268036 332640 268280
rect 351822 268268 351828 268320
rect 351880 268308 351886 268320
rect 433518 268308 433524 268320
rect 351880 268280 433524 268308
rect 351880 268268 351886 268280
rect 433518 268268 433524 268280
rect 433576 268268 433582 268320
rect 332686 268200 332692 268252
rect 332744 268240 332750 268252
rect 426434 268240 426440 268252
rect 332744 268212 426440 268240
rect 332744 268200 332750 268212
rect 426434 268200 426440 268212
rect 426492 268200 426498 268252
rect 351914 268132 351920 268184
rect 351972 268172 351978 268184
rect 427630 268172 427636 268184
rect 351972 268144 427636 268172
rect 351972 268132 351978 268144
rect 427630 268132 427636 268144
rect 427688 268132 427694 268184
rect 332778 268064 332784 268116
rect 332836 268104 332842 268116
rect 420546 268104 420552 268116
rect 332836 268076 420552 268104
rect 332836 268064 332842 268076
rect 420546 268064 420552 268076
rect 420604 268064 420610 268116
rect 666462 268064 666468 268116
rect 666520 268104 666526 268116
rect 676214 268104 676220 268116
rect 666520 268076 676220 268104
rect 666520 268064 666526 268076
rect 676214 268064 676220 268076
rect 676272 268064 676278 268116
rect 357434 268036 357440 268048
rect 332612 268008 357440 268036
rect 357434 267996 357440 268008
rect 357492 267996 357498 268048
rect 357526 267996 357532 268048
rect 357584 268036 357590 268048
rect 358722 268036 358728 268048
rect 357584 268008 358728 268036
rect 357584 267996 357590 268008
rect 358722 267996 358728 268008
rect 358780 267996 358786 268048
rect 372706 267996 372712 268048
rect 372764 268036 372770 268048
rect 382458 268036 382464 268048
rect 372764 268008 382464 268036
rect 372764 267996 372770 268008
rect 382458 267996 382464 268008
rect 382516 267996 382522 268048
rect 390002 267996 390008 268048
rect 390060 268036 390066 268048
rect 394602 268036 394608 268048
rect 390060 268008 394608 268036
rect 390060 267996 390066 268008
rect 394602 267996 394608 268008
rect 394660 267996 394666 268048
rect 400766 267996 400772 268048
rect 400824 268036 400830 268048
rect 402882 268036 402888 268048
rect 400824 268008 402888 268036
rect 400824 267996 400830 268008
rect 402882 267996 402888 268008
rect 402940 267996 402946 268048
rect 406102 267996 406108 268048
rect 406160 268036 406166 268048
rect 411990 268036 411996 268048
rect 406160 268008 411996 268036
rect 406160 267996 406166 268008
rect 411990 267996 411996 268008
rect 412048 267996 412054 268048
rect 351730 267968 351736 267980
rect 332336 267940 351736 267968
rect 351730 267928 351736 267940
rect 351788 267928 351794 267980
rect 661126 267928 661132 267980
rect 661184 267968 661190 267980
rect 676030 267968 676036 267980
rect 661184 267940 676036 267968
rect 661184 267928 661190 267940
rect 676030 267928 676036 267940
rect 676088 267928 676094 267980
rect 276474 267860 276480 267912
rect 276532 267900 276538 267912
rect 289262 267900 289268 267912
rect 276532 267872 289268 267900
rect 276532 267860 276538 267872
rect 289262 267860 289268 267872
rect 289320 267860 289326 267912
rect 327994 267860 328000 267912
rect 328052 267900 328058 267912
rect 332686 267900 332692 267912
rect 328052 267872 332692 267900
rect 328052 267860 328058 267872
rect 332686 267860 332692 267872
rect 332744 267860 332750 267912
rect 343266 267860 343272 267912
rect 343324 267900 343330 267912
rect 352006 267900 352012 267912
rect 343324 267872 352012 267900
rect 343324 267860 343330 267872
rect 352006 267860 352012 267872
rect 352064 267860 352070 267912
rect 235184 267804 237374 267832
rect 304534 267792 304540 267844
rect 304592 267832 304598 267844
rect 363782 267832 363788 267844
rect 304592 267804 363788 267832
rect 304592 267792 304598 267804
rect 363782 267792 363788 267804
rect 363840 267792 363846 267844
rect 202782 267724 202788 267776
rect 202840 267764 202846 267776
rect 206554 267764 206560 267776
rect 202840 267736 206560 267764
rect 202840 267724 202846 267736
rect 206554 267724 206560 267736
rect 206612 267724 206618 267776
rect 206646 267724 206652 267776
rect 206704 267764 206710 267776
rect 212350 267764 212356 267776
rect 206704 267736 212356 267764
rect 206704 267724 206710 267736
rect 212350 267724 212356 267736
rect 212408 267724 212414 267776
rect 227622 267724 227628 267776
rect 227680 267764 227686 267776
rect 234154 267764 234160 267776
rect 227680 267736 234160 267764
rect 227680 267724 227686 267736
rect 234154 267724 234160 267736
rect 234212 267724 234218 267776
rect 234706 267724 234712 267776
rect 234764 267764 234770 267776
rect 237742 267764 237748 267776
rect 234764 267736 237748 267764
rect 234764 267724 234770 267736
rect 237742 267724 237748 267736
rect 237800 267724 237806 267776
rect 332502 267724 332508 267776
rect 332560 267764 332566 267776
rect 376754 267764 376760 267776
rect 332560 267736 376760 267764
rect 332560 267724 332566 267736
rect 376754 267724 376760 267736
rect 376812 267724 376818 267776
rect 660942 267724 660948 267776
rect 661000 267764 661006 267776
rect 676122 267764 676128 267776
rect 661000 267736 676128 267764
rect 661000 267724 661006 267736
rect 676122 267724 676128 267736
rect 676180 267724 676186 267776
rect 359734 267656 359740 267708
rect 359792 267696 359798 267708
rect 510338 267696 510344 267708
rect 359792 267668 510344 267696
rect 359792 267656 359798 267668
rect 510338 267656 510344 267668
rect 510396 267656 510402 267708
rect 674742 267656 674748 267708
rect 674800 267696 674806 267708
rect 676030 267696 676036 267708
rect 674800 267668 676036 267696
rect 674800 267656 674806 267668
rect 676030 267656 676036 267668
rect 676088 267656 676094 267708
rect 362402 267588 362408 267640
rect 362460 267628 362466 267640
rect 517422 267628 517428 267640
rect 362460 267600 517428 267628
rect 362460 267588 362466 267600
rect 517422 267588 517428 267600
rect 517480 267588 517486 267640
rect 365070 267520 365076 267572
rect 365128 267560 365134 267572
rect 524506 267560 524512 267572
rect 365128 267532 524512 267560
rect 365128 267520 365134 267532
rect 524506 267520 524512 267532
rect 524564 267520 524570 267572
rect 367738 267452 367744 267504
rect 367796 267492 367802 267504
rect 531590 267492 531596 267504
rect 367796 267464 531596 267492
rect 367796 267452 367802 267464
rect 531590 267452 531596 267464
rect 531648 267452 531654 267504
rect 672258 267452 672264 267504
rect 672316 267492 672322 267504
rect 675938 267492 675944 267504
rect 672316 267464 675944 267492
rect 672316 267452 672322 267464
rect 675938 267452 675944 267464
rect 675996 267452 676002 267504
rect 370498 267384 370504 267436
rect 370556 267424 370562 267436
rect 538766 267424 538772 267436
rect 370556 267396 538772 267424
rect 370556 267384 370562 267396
rect 538766 267384 538772 267396
rect 538824 267384 538830 267436
rect 373534 267316 373540 267368
rect 373592 267356 373598 267368
rect 547046 267356 547052 267368
rect 373592 267328 547052 267356
rect 373592 267316 373598 267328
rect 547046 267316 547052 267328
rect 547104 267316 547110 267368
rect 374454 267248 374460 267300
rect 374512 267288 374518 267300
rect 549346 267288 549352 267300
rect 374512 267260 549352 267288
rect 374512 267248 374518 267260
rect 549346 267248 549352 267260
rect 549404 267248 549410 267300
rect 376202 267180 376208 267232
rect 376260 267220 376266 267232
rect 554130 267220 554136 267232
rect 376260 267192 554136 267220
rect 376260 267180 376266 267192
rect 554130 267180 554136 267192
rect 554188 267180 554194 267232
rect 299658 267112 299664 267164
rect 299716 267152 299722 267164
rect 350718 267152 350724 267164
rect 299716 267124 350724 267152
rect 299716 267112 299722 267124
rect 350718 267112 350724 267124
rect 350776 267112 350782 267164
rect 375834 267112 375840 267164
rect 375892 267152 375898 267164
rect 552934 267152 552940 267164
rect 375892 267124 552940 267152
rect 375892 267112 375898 267124
rect 552934 267112 552940 267124
rect 552992 267112 552998 267164
rect 300946 267044 300952 267096
rect 301004 267084 301010 267096
rect 354306 267084 354312 267096
rect 301004 267056 354312 267084
rect 301004 267044 301010 267056
rect 354306 267044 354312 267056
rect 354364 267044 354370 267096
rect 377122 267044 377128 267096
rect 377180 267084 377186 267096
rect 556430 267084 556436 267096
rect 377180 267056 556436 267084
rect 377180 267044 377186 267056
rect 556430 267044 556436 267056
rect 556488 267044 556494 267096
rect 302326 266976 302332 267028
rect 302384 267016 302390 267028
rect 357894 267016 357900 267028
rect 302384 266988 357900 267016
rect 302384 266976 302390 266988
rect 357894 266976 357900 266988
rect 357952 266976 357958 267028
rect 378502 266976 378508 267028
rect 378560 267016 378566 267028
rect 560018 267016 560024 267028
rect 378560 266988 560024 267016
rect 378560 266976 378566 266988
rect 560018 266976 560024 266988
rect 560076 266976 560082 267028
rect 303706 266908 303712 266960
rect 303764 266948 303770 266960
rect 361390 266948 361396 266960
rect 303764 266920 361396 266948
rect 303764 266908 303770 266920
rect 361390 266908 361396 266920
rect 361448 266908 361454 266960
rect 378870 266908 378876 266960
rect 378928 266948 378934 266960
rect 561214 266948 561220 266960
rect 378928 266920 561220 266948
rect 378928 266908 378934 266920
rect 561214 266908 561220 266920
rect 561272 266908 561278 266960
rect 304994 266840 305000 266892
rect 305052 266880 305058 266892
rect 364978 266880 364984 266892
rect 305052 266852 364984 266880
rect 305052 266840 305058 266852
rect 364978 266840 364984 266852
rect 365036 266840 365042 266892
rect 379790 266840 379796 266892
rect 379848 266880 379854 266892
rect 563514 266880 563520 266892
rect 379848 266852 563520 266880
rect 379848 266840 379854 266852
rect 563514 266840 563520 266852
rect 563572 266840 563578 266892
rect 306374 266772 306380 266824
rect 306432 266812 306438 266824
rect 368474 266812 368480 266824
rect 306432 266784 368480 266812
rect 306432 266772 306438 266784
rect 368474 266772 368480 266784
rect 368532 266772 368538 266824
rect 381630 266772 381636 266824
rect 381688 266812 381694 266824
rect 568298 266812 568304 266824
rect 381688 266784 568304 266812
rect 381688 266772 381694 266784
rect 568298 266772 568304 266784
rect 568356 266772 568362 266824
rect 307662 266704 307668 266756
rect 307720 266744 307726 266756
rect 372062 266744 372068 266756
rect 307720 266716 372068 266744
rect 307720 266704 307726 266716
rect 372062 266704 372068 266716
rect 372120 266704 372126 266756
rect 381170 266704 381176 266756
rect 381228 266744 381234 266756
rect 567102 266744 567108 266756
rect 381228 266716 567108 266744
rect 381228 266704 381234 266716
rect 567102 266704 567108 266716
rect 567160 266704 567166 266756
rect 309042 266636 309048 266688
rect 309100 266676 309106 266688
rect 375558 266676 375564 266688
rect 309100 266648 375564 266676
rect 309100 266636 309106 266648
rect 375558 266636 375564 266648
rect 375616 266636 375622 266688
rect 382458 266636 382464 266688
rect 382516 266676 382522 266688
rect 570690 266676 570696 266688
rect 382516 266648 570696 266676
rect 382516 266636 382522 266648
rect 570690 266636 570696 266648
rect 570748 266636 570754 266688
rect 123754 266568 123760 266620
rect 123812 266608 123818 266620
rect 214190 266608 214196 266620
rect 123812 266580 214196 266608
rect 123812 266568 123818 266580
rect 214190 266568 214196 266580
rect 214248 266568 214254 266620
rect 310330 266568 310336 266620
rect 310388 266608 310394 266620
rect 379146 266608 379152 266620
rect 310388 266580 379152 266608
rect 310388 266568 310394 266580
rect 379146 266568 379152 266580
rect 379204 266568 379210 266620
rect 384298 266568 384304 266620
rect 384356 266608 384362 266620
rect 575382 266608 575388 266620
rect 384356 266580 575388 266608
rect 384356 266568 384362 266580
rect 575382 266568 575388 266580
rect 575440 266568 575446 266620
rect 116670 266500 116676 266552
rect 116728 266540 116734 266552
rect 211522 266540 211528 266552
rect 116728 266512 211528 266540
rect 116728 266500 116734 266512
rect 211522 266500 211528 266512
rect 211580 266500 211586 266552
rect 311710 266500 311716 266552
rect 311768 266540 311774 266552
rect 382642 266540 382648 266552
rect 311768 266512 382648 266540
rect 311768 266500 311774 266512
rect 382642 266500 382648 266512
rect 382700 266500 382706 266552
rect 383838 266500 383844 266552
rect 383896 266540 383902 266552
rect 574186 266540 574192 266552
rect 383896 266512 574192 266540
rect 383896 266500 383902 266512
rect 574186 266500 574192 266512
rect 574244 266500 574250 266552
rect 72970 266432 72976 266484
rect 73028 266472 73034 266484
rect 195054 266472 195060 266484
rect 73028 266444 195060 266472
rect 73028 266432 73034 266444
rect 195054 266432 195060 266444
rect 195112 266432 195118 266484
rect 312998 266432 313004 266484
rect 313056 266472 313062 266484
rect 386230 266472 386236 266484
rect 313056 266444 386236 266472
rect 313056 266432 313062 266444
rect 386230 266432 386236 266444
rect 386288 266432 386294 266484
rect 389174 266432 389180 266484
rect 389232 266472 389238 266484
rect 588354 266472 588360 266484
rect 389232 266444 588360 266472
rect 389232 266432 389238 266444
rect 588354 266432 588360 266444
rect 588412 266432 588418 266484
rect 113174 266364 113180 266416
rect 113232 266404 113238 266416
rect 210142 266404 210148 266416
rect 113232 266376 210148 266404
rect 113232 266364 113238 266376
rect 210142 266364 210148 266376
rect 210200 266364 210206 266416
rect 315666 266364 315672 266416
rect 315724 266404 315730 266416
rect 315724 266376 391934 266404
rect 315724 266364 315730 266376
rect 68186 266296 68192 266348
rect 68244 266336 68250 266348
rect 193214 266336 193220 266348
rect 68244 266308 193220 266336
rect 68244 266296 68250 266308
rect 193214 266296 193220 266308
rect 193272 266296 193278 266348
rect 317046 266296 317052 266348
rect 317104 266336 317110 266348
rect 382182 266336 382188 266348
rect 317104 266308 382188 266336
rect 317104 266296 317110 266308
rect 382182 266296 382188 266308
rect 382240 266296 382246 266348
rect 391906 266336 391934 266376
rect 392302 266364 392308 266416
rect 392360 266404 392366 266416
rect 596634 266404 596640 266416
rect 392360 266376 596640 266404
rect 392360 266364 392366 266376
rect 596634 266364 596640 266376
rect 596692 266364 596698 266416
rect 393314 266336 393320 266348
rect 391906 266308 393320 266336
rect 393314 266296 393320 266308
rect 393372 266296 393378 266348
rect 394970 266296 394976 266348
rect 395028 266336 395034 266348
rect 603718 266336 603724 266348
rect 395028 266308 603724 266336
rect 395028 266296 395034 266308
rect 603718 266296 603724 266308
rect 603776 266296 603782 266348
rect 652938 266296 652944 266348
rect 652996 266336 653002 266348
rect 675662 266336 675668 266348
rect 652996 266308 675668 266336
rect 652996 266296 653002 266308
rect 675662 266296 675668 266308
rect 675720 266296 675726 266348
rect 357066 266228 357072 266280
rect 357124 266268 357130 266280
rect 503254 266268 503260 266280
rect 357124 266240 503260 266268
rect 357124 266228 357130 266240
rect 503254 266228 503260 266240
rect 503312 266228 503318 266280
rect 353202 266160 353208 266212
rect 353260 266200 353266 266212
rect 492582 266200 492588 266212
rect 353260 266172 492588 266200
rect 353260 266160 353266 266172
rect 492582 266160 492588 266172
rect 492640 266160 492646 266212
rect 351730 266092 351736 266144
rect 351788 266132 351794 266144
rect 489086 266132 489092 266144
rect 351788 266104 489092 266132
rect 351788 266092 351794 266104
rect 489086 266092 489092 266104
rect 489144 266092 489150 266144
rect 671890 266092 671896 266144
rect 671948 266132 671954 266144
rect 676214 266132 676220 266144
rect 671948 266104 676220 266132
rect 671948 266092 671954 266104
rect 676214 266092 676220 266104
rect 676272 266092 676278 266144
rect 347774 266024 347780 266076
rect 347832 266064 347838 266076
rect 478414 266064 478420 266076
rect 347832 266036 478420 266064
rect 347832 266024 347838 266036
rect 478414 266024 478420 266036
rect 478472 266024 478478 266076
rect 346394 265956 346400 266008
rect 346452 265996 346458 266008
rect 474918 265996 474924 266008
rect 346452 265968 474924 265996
rect 346452 265956 346458 265968
rect 474918 265956 474924 265968
rect 474976 265956 474982 266008
rect 339770 265888 339776 265940
rect 339828 265928 339834 265940
rect 457162 265928 457168 265940
rect 339828 265900 457168 265928
rect 339828 265888 339834 265900
rect 457162 265888 457168 265900
rect 457220 265888 457226 265940
rect 338390 265820 338396 265872
rect 338448 265860 338454 265872
rect 453574 265860 453580 265872
rect 338448 265832 453580 265860
rect 338448 265820 338454 265832
rect 453574 265820 453580 265832
rect 453632 265820 453638 265872
rect 317506 265752 317512 265804
rect 317564 265792 317570 265804
rect 382090 265792 382096 265804
rect 317564 265764 382096 265792
rect 317564 265752 317570 265764
rect 382090 265752 382096 265764
rect 382148 265752 382154 265804
rect 382182 265752 382188 265804
rect 382240 265792 382246 265804
rect 396902 265792 396908 265804
rect 382240 265764 396908 265792
rect 382240 265752 382246 265764
rect 396902 265752 396908 265764
rect 396960 265752 396966 265804
rect 397638 265752 397644 265804
rect 397696 265792 397702 265804
rect 511626 265792 511632 265804
rect 397696 265764 511632 265792
rect 397696 265752 397702 265764
rect 511626 265752 511632 265764
rect 511684 265752 511690 265804
rect 329466 265684 329472 265736
rect 329524 265724 329530 265736
rect 429930 265724 429936 265736
rect 329524 265696 353294 265724
rect 329524 265684 329530 265696
rect 353266 265656 353294 265696
rect 382200 265696 429936 265724
rect 382200 265656 382228 265696
rect 429930 265684 429936 265696
rect 429988 265684 429994 265736
rect 353266 265628 382228 265656
rect 382274 265616 382280 265668
rect 382332 265656 382338 265668
rect 398006 265656 398012 265668
rect 382332 265628 398012 265656
rect 382332 265616 382338 265628
rect 398006 265616 398012 265628
rect 398064 265616 398070 265668
rect 400306 265616 400312 265668
rect 400364 265656 400370 265668
rect 498838 265656 498844 265668
rect 400364 265628 498844 265656
rect 400364 265616 400370 265628
rect 498838 265616 498844 265628
rect 498896 265616 498902 265668
rect 325510 265548 325516 265600
rect 325568 265588 325574 265600
rect 419350 265588 419356 265600
rect 325568 265560 419356 265588
rect 325568 265548 325574 265560
rect 419350 265548 419356 265560
rect 419408 265548 419414 265600
rect 324130 265480 324136 265532
rect 324188 265520 324194 265532
rect 415762 265520 415768 265532
rect 324188 265492 415768 265520
rect 324188 265480 324194 265492
rect 415762 265480 415768 265492
rect 415820 265480 415826 265532
rect 322842 265412 322848 265464
rect 322900 265452 322906 265464
rect 412266 265452 412272 265464
rect 322900 265424 412272 265452
rect 322900 265412 322906 265424
rect 412266 265412 412272 265424
rect 412324 265412 412330 265464
rect 321462 265344 321468 265396
rect 321520 265384 321526 265396
rect 408678 265384 408684 265396
rect 321520 265356 408684 265384
rect 321520 265344 321526 265356
rect 408678 265344 408684 265356
rect 408736 265344 408742 265396
rect 674742 265344 674748 265396
rect 674800 265384 674806 265396
rect 676030 265384 676036 265396
rect 674800 265356 676036 265384
rect 674800 265344 674806 265356
rect 676030 265344 676036 265356
rect 676088 265344 676094 265396
rect 318334 265276 318340 265328
rect 318392 265316 318398 265328
rect 400398 265316 400404 265328
rect 318392 265288 400404 265316
rect 318392 265276 318398 265288
rect 400398 265276 400404 265288
rect 400456 265276 400462 265328
rect 402974 265276 402980 265328
rect 403032 265316 403038 265328
rect 471974 265316 471980 265328
rect 403032 265288 471980 265316
rect 403032 265276 403038 265288
rect 471974 265276 471980 265288
rect 472032 265276 472038 265328
rect 314378 265208 314384 265260
rect 314436 265248 314442 265260
rect 389726 265248 389732 265260
rect 314436 265220 389732 265248
rect 314436 265208 314442 265220
rect 389726 265208 389732 265220
rect 389784 265208 389790 265260
rect 319714 265140 319720 265192
rect 319772 265180 319778 265192
rect 403986 265180 403992 265192
rect 319772 265152 403992 265180
rect 319772 265140 319778 265152
rect 403986 265140 403992 265152
rect 404044 265140 404050 265192
rect 675754 265044 675760 265056
rect 670666 265016 675760 265044
rect 658274 264936 658280 264988
rect 658332 264976 658338 264988
rect 670666 264976 670694 265016
rect 675754 265004 675760 265016
rect 675812 265004 675818 265056
rect 658332 264948 670694 264976
rect 658332 264936 658338 264948
rect 673178 264936 673184 264988
rect 673236 264976 673242 264988
rect 676214 264976 676220 264988
rect 673236 264948 676220 264976
rect 673236 264936 673242 264948
rect 676214 264936 676220 264948
rect 676272 264936 676278 264988
rect 674190 263032 674196 263084
rect 674248 263072 674254 263084
rect 676030 263072 676036 263084
rect 674248 263044 676036 263072
rect 674248 263032 674254 263044
rect 676030 263032 676036 263044
rect 676088 263032 676094 263084
rect 673730 262352 673736 262404
rect 673788 262392 673794 262404
rect 675938 262392 675944 262404
rect 673788 262364 675944 262392
rect 673788 262352 673794 262364
rect 675938 262352 675944 262364
rect 675996 262352 676002 262404
rect 674006 262284 674012 262336
rect 674064 262324 674070 262336
rect 676122 262324 676128 262336
rect 674064 262296 676128 262324
rect 674064 262284 674070 262296
rect 676122 262284 676128 262296
rect 676180 262284 676186 262336
rect 418062 262216 418068 262268
rect 418120 262256 418126 262268
rect 571702 262256 571708 262268
rect 418120 262228 571708 262256
rect 418120 262216 418126 262228
rect 571702 262216 571708 262228
rect 571760 262216 571766 262268
rect 674282 262216 674288 262268
rect 674340 262256 674346 262268
rect 676030 262256 676036 262268
rect 674340 262228 676036 262256
rect 674340 262216 674346 262228
rect 676030 262216 676036 262228
rect 676088 262216 676094 262268
rect 674098 261808 674104 261860
rect 674156 261848 674162 261860
rect 676030 261848 676036 261860
rect 674156 261820 676036 261848
rect 674156 261808 674162 261820
rect 676030 261808 676036 261820
rect 676088 261808 676094 261860
rect 673454 260176 673460 260228
rect 673512 260216 673518 260228
rect 675570 260216 675576 260228
rect 673512 260188 675576 260216
rect 673512 260176 673518 260188
rect 675570 260176 675576 260188
rect 675628 260176 675634 260228
rect 673546 259700 673552 259752
rect 673604 259740 673610 259752
rect 675570 259740 675576 259752
rect 673604 259712 675576 259740
rect 673604 259700 673610 259712
rect 675570 259700 675576 259712
rect 675628 259700 675634 259752
rect 674466 259632 674472 259684
rect 674524 259672 674530 259684
rect 676122 259672 676128 259684
rect 674524 259644 676128 259672
rect 674524 259632 674530 259644
rect 676122 259632 676128 259644
rect 676180 259632 676186 259684
rect 674374 259564 674380 259616
rect 674432 259604 674438 259616
rect 675938 259604 675944 259616
rect 674432 259576 675944 259604
rect 674432 259564 674438 259576
rect 675938 259564 675944 259576
rect 675996 259564 676002 259616
rect 675018 259496 675024 259548
rect 675076 259536 675082 259548
rect 676122 259536 676128 259548
rect 675076 259508 676128 259536
rect 675076 259496 675082 259508
rect 676122 259496 676128 259508
rect 676180 259496 676186 259548
rect 52270 259428 52276 259480
rect 52328 259468 52334 259480
rect 184934 259468 184940 259480
rect 52328 259440 184940 259468
rect 52328 259428 52334 259440
rect 184934 259428 184940 259440
rect 184992 259428 184998 259480
rect 417786 259428 417792 259480
rect 417844 259468 417850 259480
rect 571794 259468 571800 259480
rect 417844 259440 571800 259468
rect 417844 259428 417850 259440
rect 571794 259428 571800 259440
rect 571852 259428 571858 259480
rect 675202 259428 675208 259480
rect 675260 259468 675266 259480
rect 676030 259468 676036 259480
rect 675260 259440 676036 259468
rect 675260 259428 675266 259440
rect 676030 259428 676036 259440
rect 676088 259428 676094 259480
rect 41506 258340 41512 258392
rect 41564 258380 41570 258392
rect 48406 258380 48412 258392
rect 41564 258352 48412 258380
rect 41564 258340 41570 258352
rect 48406 258340 48412 258352
rect 48464 258340 48470 258392
rect 41782 257796 41788 257848
rect 41840 257836 41846 257848
rect 53926 257836 53932 257848
rect 41840 257808 53932 257836
rect 41840 257796 41846 257808
rect 53926 257796 53932 257808
rect 53984 257796 53990 257848
rect 41506 257524 41512 257576
rect 41564 257564 41570 257576
rect 50982 257564 50988 257576
rect 41564 257536 50988 257564
rect 41564 257524 41570 257536
rect 50982 257524 50988 257536
rect 51040 257524 51046 257576
rect 41782 256844 41788 256896
rect 41840 256884 41846 256896
rect 45830 256884 45836 256896
rect 41840 256856 45836 256884
rect 41840 256844 41846 256856
rect 45830 256844 45836 256856
rect 45888 256844 45894 256896
rect 672810 256844 672816 256896
rect 672868 256884 672874 256896
rect 678974 256884 678980 256896
rect 672868 256856 678980 256884
rect 672868 256844 672874 256856
rect 678974 256844 678980 256856
rect 679032 256844 679038 256896
rect 673638 256776 673644 256828
rect 673696 256816 673702 256828
rect 676122 256816 676128 256828
rect 673696 256788 676128 256816
rect 673696 256776 673702 256788
rect 676122 256776 676128 256788
rect 676180 256776 676186 256828
rect 418338 256708 418344 256760
rect 418396 256748 418402 256760
rect 571518 256748 571524 256760
rect 418396 256720 571524 256748
rect 418396 256708 418402 256720
rect 571518 256708 571524 256720
rect 571576 256708 571582 256760
rect 673822 256708 673828 256760
rect 673880 256748 673886 256760
rect 676030 256748 676036 256760
rect 673880 256720 676036 256748
rect 673880 256708 673886 256720
rect 676030 256708 676036 256720
rect 676088 256708 676094 256760
rect 674742 255280 674748 255332
rect 674800 255320 674806 255332
rect 675662 255320 675668 255332
rect 674800 255292 675668 255320
rect 674800 255280 674806 255292
rect 675662 255280 675668 255292
rect 675720 255280 675726 255332
rect 674650 255212 674656 255264
rect 674708 255252 674714 255264
rect 675754 255252 675760 255264
rect 674708 255224 675760 255252
rect 674708 255212 674714 255224
rect 675754 255212 675760 255224
rect 675812 255212 675818 255264
rect 416774 253920 416780 253972
rect 416832 253960 416838 253972
rect 574094 253960 574100 253972
rect 416832 253932 574100 253960
rect 416832 253920 416838 253932
rect 574094 253920 574100 253932
rect 574152 253920 574158 253972
rect 52178 251200 52184 251252
rect 52236 251240 52242 251252
rect 184934 251240 184940 251252
rect 52236 251212 184940 251240
rect 52236 251200 52242 251212
rect 184934 251200 184940 251212
rect 184992 251200 184998 251252
rect 416774 251200 416780 251252
rect 416832 251240 416838 251252
rect 572622 251240 572628 251252
rect 416832 251212 572628 251240
rect 416832 251200 416838 251212
rect 572622 251200 572628 251212
rect 572680 251200 572686 251252
rect 675754 251200 675760 251252
rect 675812 251200 675818 251252
rect 675772 250980 675800 251200
rect 675754 250928 675760 250980
rect 675812 250928 675818 250980
rect 675202 250384 675208 250436
rect 675260 250424 675266 250436
rect 675478 250424 675484 250436
rect 675260 250396 675484 250424
rect 675260 250384 675266 250396
rect 675478 250384 675484 250396
rect 675536 250384 675542 250436
rect 33042 249772 33048 249824
rect 33100 249812 33106 249824
rect 43622 249812 43628 249824
rect 33100 249784 43628 249812
rect 33100 249772 33106 249784
rect 43622 249772 43628 249784
rect 43680 249772 43686 249824
rect 674190 249568 674196 249620
rect 674248 249608 674254 249620
rect 675386 249608 675392 249620
rect 674248 249580 675392 249608
rect 674248 249568 674254 249580
rect 675386 249568 675392 249580
rect 675444 249568 675450 249620
rect 416774 248412 416780 248464
rect 416832 248452 416838 248464
rect 569862 248452 569868 248464
rect 416832 248424 569868 248452
rect 416832 248412 416838 248424
rect 569862 248412 569868 248424
rect 569920 248412 569926 248464
rect 674282 247868 674288 247920
rect 674340 247908 674346 247920
rect 675478 247908 675484 247920
rect 674340 247880 675484 247908
rect 674340 247868 674346 247880
rect 675478 247868 675484 247880
rect 675536 247868 675542 247920
rect 41506 247664 41512 247716
rect 41564 247704 41570 247716
rect 45922 247704 45928 247716
rect 41564 247676 45928 247704
rect 41564 247664 41570 247676
rect 45922 247664 45928 247676
rect 45980 247664 45986 247716
rect 41506 247256 41512 247308
rect 41564 247296 41570 247308
rect 45830 247296 45836 247308
rect 41564 247268 45836 247296
rect 41564 247256 41570 247268
rect 45830 247256 45836 247268
rect 45888 247256 45894 247308
rect 674466 247256 674472 247308
rect 674524 247296 674530 247308
rect 675386 247296 675392 247308
rect 674524 247268 675392 247296
rect 674524 247256 674530 247268
rect 675386 247256 675392 247268
rect 675444 247256 675450 247308
rect 674006 247120 674012 247172
rect 674064 247160 674070 247172
rect 674466 247160 674472 247172
rect 674064 247132 674472 247160
rect 674064 247120 674070 247132
rect 674466 247120 674472 247132
rect 674524 247120 674530 247172
rect 41506 246848 41512 246900
rect 41564 246888 41570 246900
rect 45738 246888 45744 246900
rect 41564 246860 45744 246888
rect 41564 246848 41570 246860
rect 45738 246848 45744 246860
rect 45796 246848 45802 246900
rect 674374 246508 674380 246560
rect 674432 246548 674438 246560
rect 675386 246548 675392 246560
rect 674432 246520 675392 246548
rect 674432 246508 674438 246520
rect 675386 246508 675392 246520
rect 675444 246508 675450 246560
rect 675110 246032 675116 246084
rect 675168 246072 675174 246084
rect 675386 246072 675392 246084
rect 675168 246044 675392 246072
rect 675168 246032 675174 246044
rect 675386 246032 675392 246044
rect 675444 246032 675450 246084
rect 43622 244740 43628 244792
rect 43680 244780 43686 244792
rect 43898 244780 43904 244792
rect 43680 244752 43904 244780
rect 43680 244740 43686 244752
rect 43898 244740 43904 244752
rect 43956 244740 43962 244792
rect 43346 244604 43352 244656
rect 43404 244644 43410 244656
rect 43622 244644 43628 244656
rect 43404 244616 43628 244644
rect 43404 244604 43410 244616
rect 43622 244604 43628 244616
rect 43680 244604 43686 244656
rect 42886 244536 42892 244588
rect 42944 244576 42950 244588
rect 43530 244576 43536 244588
rect 42944 244548 43536 244576
rect 42944 244536 42950 244548
rect 43530 244536 43536 244548
rect 43588 244536 43594 244588
rect 42702 244468 42708 244520
rect 42760 244508 42766 244520
rect 43346 244508 43352 244520
rect 42760 244480 43352 244508
rect 42760 244468 42766 244480
rect 43346 244468 43352 244480
rect 43404 244468 43410 244520
rect 33042 244400 33048 244452
rect 33100 244440 33106 244452
rect 42886 244440 42892 244452
rect 33100 244412 42892 244440
rect 33100 244400 33106 244412
rect 42886 244400 42892 244412
rect 42944 244400 42950 244452
rect 32858 244332 32864 244384
rect 32916 244372 32922 244384
rect 43162 244372 43168 244384
rect 32916 244344 43168 244372
rect 32916 244332 32922 244344
rect 43162 244332 43168 244344
rect 43220 244332 43226 244384
rect 32950 244264 32956 244316
rect 33008 244304 33014 244316
rect 42978 244304 42984 244316
rect 33008 244276 42984 244304
rect 33008 244264 33014 244276
rect 42978 244264 42984 244276
rect 43036 244264 43042 244316
rect 31662 244196 31668 244248
rect 31720 244236 31726 244248
rect 42702 244236 42708 244248
rect 31720 244208 42708 244236
rect 31720 244196 31726 244208
rect 42702 244196 42708 244208
rect 42760 244196 42766 244248
rect 673730 243584 673736 243636
rect 673788 243624 673794 243636
rect 675294 243624 675300 243636
rect 673788 243596 675300 243624
rect 673788 243584 673794 243596
rect 675294 243584 675300 243596
rect 675352 243584 675358 243636
rect 52086 242904 52092 242956
rect 52144 242944 52150 242956
rect 184934 242944 184940 242956
rect 52144 242916 184940 242944
rect 52144 242904 52150 242916
rect 184934 242904 184940 242916
rect 184992 242904 184998 242956
rect 673822 242904 673828 242956
rect 673880 242944 673886 242956
rect 675294 242944 675300 242956
rect 673880 242916 675300 242944
rect 673880 242904 673886 242916
rect 675294 242904 675300 242916
rect 675352 242904 675358 242956
rect 38286 242836 38292 242888
rect 38344 242876 38350 242888
rect 42794 242876 42800 242888
rect 38344 242848 42800 242876
rect 38344 242836 38350 242848
rect 42794 242836 42800 242848
rect 42852 242836 42858 242888
rect 673546 242156 673552 242208
rect 673604 242196 673610 242208
rect 675386 242196 675392 242208
rect 673604 242168 675392 242196
rect 673604 242156 673610 242168
rect 675386 242156 675392 242168
rect 675444 242156 675450 242208
rect 674466 241884 674472 241936
rect 674524 241924 674530 241936
rect 675294 241924 675300 241936
rect 674524 241896 675300 241924
rect 674524 241884 674530 241896
rect 675294 241884 675300 241896
rect 675352 241884 675358 241936
rect 673638 241544 673644 241596
rect 673696 241584 673702 241596
rect 675386 241584 675392 241596
rect 673696 241556 675392 241584
rect 673696 241544 673702 241556
rect 675386 241544 675392 241556
rect 675444 241544 675450 241596
rect 673454 240524 673460 240576
rect 673512 240564 673518 240576
rect 675386 240564 675392 240576
rect 673512 240536 675392 240564
rect 673512 240524 673518 240536
rect 675386 240524 675392 240536
rect 675444 240524 675450 240576
rect 42150 240320 42156 240372
rect 42208 240360 42214 240372
rect 43714 240360 43720 240372
rect 42208 240332 43720 240360
rect 42208 240320 42214 240332
rect 43714 240320 43720 240332
rect 43772 240320 43778 240372
rect 224126 238552 224132 238604
rect 224184 238552 224190 238604
rect 42150 238416 42156 238468
rect 42208 238456 42214 238468
rect 42702 238456 42708 238468
rect 42208 238428 42708 238456
rect 42208 238416 42214 238428
rect 42702 238416 42708 238428
rect 42760 238416 42766 238468
rect 224144 238400 224172 238552
rect 224126 238348 224132 238400
rect 224184 238348 224190 238400
rect 161382 237328 161388 237380
rect 161440 237368 161446 237380
rect 237190 237368 237196 237380
rect 161440 237340 237196 237368
rect 161440 237328 161446 237340
rect 237190 237328 237196 237340
rect 237248 237328 237254 237380
rect 238938 237328 238944 237380
rect 238996 237368 239002 237380
rect 266722 237368 266728 237380
rect 238996 237340 266728 237368
rect 238996 237328 239002 237340
rect 266722 237328 266728 237340
rect 266780 237328 266786 237380
rect 329190 237328 329196 237380
rect 329248 237368 329254 237380
rect 375742 237368 375748 237380
rect 329248 237340 375748 237368
rect 329248 237328 329254 237340
rect 375742 237328 375748 237340
rect 375800 237328 375806 237380
rect 395430 237328 395436 237380
rect 395488 237368 395494 237380
rect 533982 237368 533988 237380
rect 395488 237340 533988 237368
rect 395488 237328 395494 237340
rect 533982 237328 533988 237340
rect 534040 237328 534046 237380
rect 165430 237260 165436 237312
rect 165488 237300 165494 237312
rect 240410 237300 240416 237312
rect 165488 237272 240416 237300
rect 165488 237260 165494 237272
rect 240410 237260 240416 237272
rect 240468 237260 240474 237312
rect 241606 237260 241612 237312
rect 241664 237300 241670 237312
rect 269574 237300 269580 237312
rect 241664 237272 269580 237300
rect 241664 237260 241670 237272
rect 269574 237260 269580 237272
rect 269632 237260 269638 237312
rect 314930 237260 314936 237312
rect 314988 237300 314994 237312
rect 342714 237300 342720 237312
rect 314988 237272 342720 237300
rect 314988 237260 314994 237272
rect 342714 237260 342720 237272
rect 342772 237260 342778 237312
rect 397270 237260 397276 237312
rect 397328 237300 397334 237312
rect 535454 237300 535460 237312
rect 397328 237272 535460 237300
rect 397328 237260 397334 237272
rect 535454 237260 535460 237272
rect 535512 237260 535518 237312
rect 142154 237192 142160 237244
rect 142212 237232 142218 237244
rect 218974 237232 218980 237244
rect 142212 237204 218980 237232
rect 142212 237192 142218 237204
rect 218974 237192 218980 237204
rect 219032 237192 219038 237244
rect 254854 237192 254860 237244
rect 254912 237232 254918 237244
rect 263870 237232 263876 237244
rect 254912 237204 263876 237232
rect 254912 237192 254918 237204
rect 263870 237192 263876 237204
rect 263928 237192 263934 237244
rect 312078 237192 312084 237244
rect 312136 237232 312142 237244
rect 334434 237232 334440 237244
rect 312136 237204 334440 237232
rect 312136 237192 312142 237204
rect 334434 237192 334440 237204
rect 334492 237192 334498 237244
rect 399386 237192 399392 237244
rect 399444 237232 399450 237244
rect 539502 237232 539508 237244
rect 399444 237204 539508 237232
rect 399444 237192 399450 237204
rect 539502 237192 539508 237204
rect 539560 237192 539566 237244
rect 159818 237124 159824 237176
rect 159876 237164 159882 237176
rect 237558 237164 237564 237176
rect 159876 237136 237564 237164
rect 159876 237124 159882 237136
rect 237558 237124 237564 237136
rect 237616 237124 237622 237176
rect 238846 237124 238852 237176
rect 238904 237164 238910 237176
rect 265342 237164 265348 237176
rect 238904 237136 265348 237164
rect 238904 237124 238910 237136
rect 265342 237124 265348 237136
rect 265400 237124 265406 237176
rect 302418 237124 302424 237176
rect 302476 237164 302482 237176
rect 312814 237164 312820 237176
rect 302476 237136 312820 237164
rect 302476 237124 302482 237136
rect 312814 237124 312820 237136
rect 312872 237124 312878 237176
rect 317414 237124 317420 237176
rect 317472 237164 317478 237176
rect 329742 237164 329748 237176
rect 317472 237136 329748 237164
rect 317472 237124 317478 237136
rect 329742 237124 329748 237136
rect 329800 237124 329806 237176
rect 400490 237124 400496 237176
rect 400548 237164 400554 237176
rect 542262 237164 542268 237176
rect 400548 237136 542268 237164
rect 400548 237124 400554 237136
rect 542262 237124 542268 237136
rect 542320 237124 542326 237176
rect 153194 237056 153200 237108
rect 153252 237096 153258 237108
rect 234338 237096 234344 237108
rect 153252 237068 234344 237096
rect 153252 237056 153258 237068
rect 234338 237056 234344 237068
rect 234396 237056 234402 237108
rect 242802 237056 242808 237108
rect 242860 237096 242866 237108
rect 272150 237096 272156 237108
rect 242860 237068 272156 237096
rect 242860 237056 242866 237068
rect 272150 237056 272156 237068
rect 272208 237056 272214 237108
rect 401134 237056 401140 237108
rect 401192 237096 401198 237108
rect 545114 237096 545120 237108
rect 401192 237068 545120 237096
rect 401192 237056 401198 237068
rect 545114 237056 545120 237068
rect 545172 237056 545178 237108
rect 147582 236988 147588 237040
rect 147640 237028 147646 237040
rect 229002 237028 229008 237040
rect 147640 237000 229008 237028
rect 147640 236988 147646 237000
rect 229002 236988 229008 237000
rect 229060 236988 229066 237040
rect 245470 236988 245476 237040
rect 245528 237028 245534 237040
rect 273530 237028 273536 237040
rect 245528 237000 273536 237028
rect 245528 236988 245534 237000
rect 273530 236988 273536 237000
rect 273588 236988 273594 237040
rect 302786 236988 302792 237040
rect 302844 237028 302850 237040
rect 309778 237028 309784 237040
rect 302844 237000 309784 237028
rect 302844 236988 302850 237000
rect 309778 236988 309784 237000
rect 309836 236988 309842 237040
rect 405090 236988 405096 237040
rect 405148 237028 405154 237040
rect 413462 237028 413468 237040
rect 405148 237000 413468 237028
rect 405148 236988 405154 237000
rect 413462 236988 413468 237000
rect 413520 236988 413526 237040
rect 413554 236988 413560 237040
rect 413612 237028 413618 237040
rect 545022 237028 545028 237040
rect 413612 237000 545028 237028
rect 413612 236988 413618 237000
rect 545022 236988 545028 237000
rect 545080 236988 545086 237040
rect 136542 236920 136548 236972
rect 136600 236960 136606 236972
rect 216122 236960 216128 236972
rect 136600 236932 216128 236960
rect 136600 236920 136606 236932
rect 216122 236920 216128 236932
rect 216180 236920 216186 236972
rect 223482 236920 223488 236972
rect 223540 236960 223546 236972
rect 254854 236960 254860 236972
rect 223540 236932 254860 236960
rect 223540 236920 223546 236932
rect 254854 236920 254860 236932
rect 254912 236920 254918 236972
rect 258074 236920 258080 236972
rect 258132 236960 258138 236972
rect 258132 236932 258304 236960
rect 258132 236920 258138 236932
rect 128262 236852 128268 236904
rect 128320 236892 128326 236904
rect 197262 236892 197268 236904
rect 128320 236864 197268 236892
rect 128320 236852 128326 236864
rect 197262 236852 197268 236864
rect 197320 236852 197326 236904
rect 206370 236852 206376 236904
rect 206428 236892 206434 236904
rect 226150 236892 226156 236904
rect 206428 236864 226156 236892
rect 206428 236852 206434 236864
rect 226150 236852 226156 236864
rect 226208 236852 226214 236904
rect 226242 236852 226248 236904
rect 226300 236892 226306 236904
rect 258166 236892 258172 236904
rect 226300 236864 258172 236892
rect 226300 236852 226306 236864
rect 258166 236852 258172 236864
rect 258224 236852 258230 236904
rect 258276 236892 258304 236932
rect 264698 236920 264704 236972
rect 264756 236960 264762 236972
rect 280982 236960 280988 236972
rect 264756 236932 280988 236960
rect 264756 236920 264762 236932
rect 280982 236920 280988 236932
rect 281040 236920 281046 236972
rect 301682 236920 301688 236972
rect 301740 236960 301746 236972
rect 309962 236960 309968 236972
rect 301740 236932 309968 236960
rect 301740 236920 301746 236932
rect 309962 236920 309968 236932
rect 310020 236920 310026 236972
rect 325970 236920 325976 236972
rect 326028 236960 326034 236972
rect 343358 236960 343364 236972
rect 326028 236932 343364 236960
rect 326028 236920 326034 236932
rect 343358 236920 343364 236932
rect 343416 236920 343422 236972
rect 399018 236920 399024 236972
rect 399076 236960 399082 236972
rect 542354 236960 542360 236972
rect 399076 236932 542360 236960
rect 399076 236920 399082 236932
rect 542354 236920 542360 236932
rect 542412 236920 542418 236972
rect 277486 236892 277492 236904
rect 258276 236864 277492 236892
rect 277486 236852 277492 236864
rect 277544 236852 277550 236904
rect 318794 236852 318800 236904
rect 318852 236892 318858 236904
rect 338114 236892 338120 236904
rect 318852 236864 338120 236892
rect 318852 236852 318858 236864
rect 338114 236852 338120 236864
rect 338172 236852 338178 236904
rect 402974 236852 402980 236904
rect 403032 236892 403038 236904
rect 550358 236892 550364 236904
rect 403032 236864 550364 236892
rect 403032 236852 403038 236864
rect 550358 236852 550364 236864
rect 550416 236852 550422 236904
rect 674374 236852 674380 236904
rect 674432 236892 674438 236904
rect 675386 236892 675392 236904
rect 674432 236864 675392 236892
rect 674432 236852 674438 236864
rect 675386 236852 675392 236864
rect 675444 236852 675450 236904
rect 155862 236784 155868 236836
rect 155920 236824 155926 236836
rect 234706 236824 234712 236836
rect 155920 236796 234712 236824
rect 155920 236784 155926 236796
rect 234706 236784 234712 236796
rect 234764 236784 234770 236836
rect 241422 236784 241428 236836
rect 241480 236824 241486 236836
rect 271046 236824 271052 236836
rect 241480 236796 271052 236824
rect 241480 236784 241486 236796
rect 271046 236784 271052 236796
rect 271104 236784 271110 236836
rect 320266 236784 320272 236836
rect 320324 236824 320330 236836
rect 340874 236824 340880 236836
rect 320324 236796 340880 236824
rect 320324 236784 320330 236796
rect 340874 236784 340880 236796
rect 340932 236784 340938 236836
rect 403342 236784 403348 236836
rect 403400 236824 403406 236836
rect 550542 236824 550548 236836
rect 403400 236796 550548 236824
rect 403400 236784 403406 236796
rect 550542 236784 550548 236796
rect 550600 236784 550606 236836
rect 139302 236716 139308 236768
rect 139360 236756 139366 236768
rect 218606 236756 218612 236768
rect 139360 236728 218612 236756
rect 139360 236716 139366 236728
rect 218606 236716 218612 236728
rect 218664 236716 218670 236768
rect 220722 236716 220728 236768
rect 220780 236756 220786 236768
rect 264238 236756 264244 236768
rect 220780 236728 264244 236756
rect 220780 236716 220786 236728
rect 264238 236716 264244 236728
rect 264296 236716 264302 236768
rect 264882 236716 264888 236768
rect 264940 236756 264946 236768
rect 281718 236756 281724 236768
rect 264940 236728 281724 236756
rect 264940 236716 264946 236728
rect 281718 236716 281724 236728
rect 281776 236716 281782 236768
rect 324498 236716 324504 236768
rect 324556 236756 324562 236768
rect 343266 236756 343272 236768
rect 324556 236728 343272 236756
rect 324556 236716 324562 236728
rect 343266 236716 343272 236728
rect 343324 236716 343330 236768
rect 405458 236716 405464 236768
rect 405516 236756 405522 236768
rect 413646 236756 413652 236768
rect 405516 236728 413652 236756
rect 405516 236716 405522 236728
rect 413646 236716 413652 236728
rect 413704 236716 413710 236768
rect 413738 236716 413744 236768
rect 413796 236756 413802 236768
rect 547782 236756 547788 236768
rect 413796 236728 547788 236756
rect 413796 236716 413802 236728
rect 547782 236716 547788 236728
rect 547840 236716 547846 236768
rect 42150 236648 42156 236700
rect 42208 236688 42214 236700
rect 42886 236688 42892 236700
rect 42208 236660 42892 236688
rect 42208 236648 42214 236660
rect 42886 236648 42892 236660
rect 42944 236648 42950 236700
rect 117222 236648 117228 236700
rect 117280 236688 117286 236700
rect 199746 236688 199752 236700
rect 117280 236660 199752 236688
rect 117280 236648 117286 236660
rect 199746 236648 199752 236660
rect 199804 236648 199810 236700
rect 200850 236648 200856 236700
rect 200908 236688 200914 236700
rect 252462 236688 252468 236700
rect 200908 236660 252468 236688
rect 200908 236648 200914 236660
rect 252462 236648 252468 236660
rect 252520 236648 252526 236700
rect 253198 236648 253204 236700
rect 253256 236688 253262 236700
rect 263226 236688 263232 236700
rect 253256 236660 263232 236688
rect 253256 236648 253262 236660
rect 263226 236648 263232 236660
rect 263284 236648 263290 236700
rect 269298 236688 269304 236700
rect 264946 236660 269304 236688
rect 150342 236580 150348 236632
rect 150400 236620 150406 236632
rect 231854 236620 231860 236632
rect 150400 236592 231860 236620
rect 150400 236580 150406 236592
rect 231854 236580 231860 236592
rect 231912 236580 231918 236632
rect 237282 236580 237288 236632
rect 237340 236620 237346 236632
rect 264946 236620 264974 236660
rect 269298 236648 269304 236660
rect 269356 236648 269362 236700
rect 303154 236648 303160 236700
rect 303212 236688 303218 236700
rect 312630 236688 312636 236700
rect 303212 236660 312636 236688
rect 303212 236648 303218 236660
rect 312630 236648 312636 236660
rect 312688 236648 312694 236700
rect 404722 236648 404728 236700
rect 404780 236688 404786 236700
rect 552290 236688 552296 236700
rect 404780 236660 552296 236688
rect 404780 236648 404786 236660
rect 552290 236648 552296 236660
rect 552348 236648 552354 236700
rect 237340 236592 264974 236620
rect 237340 236580 237346 236592
rect 270402 236580 270408 236632
rect 270460 236620 270466 236632
rect 284570 236620 284576 236632
rect 270460 236592 284576 236620
rect 270460 236580 270466 236592
rect 284570 236580 284576 236592
rect 284628 236580 284634 236632
rect 406838 236580 406844 236632
rect 406896 236620 406902 236632
rect 557534 236620 557540 236632
rect 406896 236592 557540 236620
rect 406896 236580 406902 236592
rect 557534 236580 557540 236592
rect 557592 236580 557598 236632
rect 142062 236512 142068 236564
rect 142120 236552 142126 236564
rect 206370 236552 206376 236564
rect 142120 236524 206376 236552
rect 142120 236512 142126 236524
rect 206370 236512 206376 236524
rect 206428 236512 206434 236564
rect 206480 236524 226334 236552
rect 119982 236444 119988 236496
rect 120040 236484 120046 236496
rect 202598 236484 202604 236496
rect 120040 236456 202604 236484
rect 120040 236444 120046 236456
rect 202598 236444 202604 236456
rect 202656 236444 202662 236496
rect 203242 236444 203248 236496
rect 203300 236484 203306 236496
rect 206480 236484 206508 236524
rect 203300 236456 206508 236484
rect 203300 236444 203306 236456
rect 209682 236444 209688 236496
rect 209740 236484 209746 236496
rect 226150 236484 226156 236496
rect 209740 236456 226156 236484
rect 209740 236444 209746 236456
rect 226150 236444 226156 236456
rect 226208 236444 226214 236496
rect 226306 236484 226334 236524
rect 239950 236512 239956 236564
rect 240008 236552 240014 236564
rect 270678 236552 270684 236564
rect 240008 236524 270684 236552
rect 240008 236512 240014 236524
rect 270678 236512 270684 236524
rect 270736 236512 270742 236564
rect 407206 236512 407212 236564
rect 407264 236552 407270 236564
rect 413370 236552 413376 236564
rect 407264 236524 413376 236552
rect 407264 236512 407270 236524
rect 413370 236512 413376 236524
rect 413428 236512 413434 236564
rect 413462 236512 413468 236564
rect 413520 236552 413526 236564
rect 556154 236552 556160 236564
rect 413520 236524 556160 236552
rect 413520 236512 413526 236524
rect 556154 236512 556160 236524
rect 556212 236512 556218 236564
rect 255314 236484 255320 236496
rect 226306 236456 255320 236484
rect 255314 236444 255320 236456
rect 255372 236444 255378 236496
rect 259270 236444 259276 236496
rect 259328 236484 259334 236496
rect 279970 236484 279976 236496
rect 259328 236456 279976 236484
rect 259328 236444 259334 236456
rect 279970 236444 279976 236456
rect 280028 236444 280034 236496
rect 317782 236444 317788 236496
rect 317840 236484 317846 236496
rect 348142 236484 348148 236496
rect 317840 236456 348148 236484
rect 317840 236444 317846 236456
rect 348142 236444 348148 236456
rect 348200 236444 348206 236496
rect 407574 236444 407580 236496
rect 407632 236484 407638 236496
rect 413554 236484 413560 236496
rect 407632 236456 413560 236484
rect 407632 236444 407638 236456
rect 413554 236444 413560 236456
rect 413612 236444 413618 236496
rect 413646 236444 413652 236496
rect 413704 236484 413710 236496
rect 556062 236484 556068 236496
rect 413704 236456 556068 236484
rect 413704 236444 413710 236456
rect 556062 236444 556068 236456
rect 556120 236444 556126 236496
rect 125502 236376 125508 236428
rect 125560 236416 125566 236428
rect 215754 236416 215760 236428
rect 125560 236388 215760 236416
rect 125560 236376 125566 236388
rect 215754 236376 215760 236388
rect 215812 236376 215818 236428
rect 220630 236376 220636 236428
rect 220688 236416 220694 236428
rect 253198 236416 253204 236428
rect 220688 236388 253204 236416
rect 220688 236376 220694 236388
rect 253198 236376 253204 236388
rect 253256 236376 253262 236428
rect 261018 236416 261024 236428
rect 253308 236388 261024 236416
rect 122742 236308 122748 236360
rect 122800 236348 122806 236360
rect 213270 236348 213276 236360
rect 122800 236320 213276 236348
rect 122800 236308 122806 236320
rect 213270 236308 213276 236320
rect 213328 236308 213334 236360
rect 216674 236308 216680 236360
rect 216732 236348 216738 236360
rect 253308 236348 253336 236388
rect 261018 236376 261024 236388
rect 261076 236376 261082 236428
rect 264790 236376 264796 236428
rect 264848 236416 264854 236428
rect 282822 236416 282828 236428
rect 264848 236388 282828 236416
rect 264848 236376 264854 236388
rect 282822 236376 282828 236388
rect 282880 236376 282886 236428
rect 302050 236376 302056 236428
rect 302108 236416 302114 236428
rect 312262 236416 312268 236428
rect 302108 236388 312268 236416
rect 302108 236376 302114 236388
rect 312262 236376 312268 236388
rect 312320 236376 312326 236428
rect 316310 236376 316316 236428
rect 316368 236416 316374 236428
rect 345382 236416 345388 236428
rect 316368 236388 345388 236416
rect 316368 236376 316374 236388
rect 345382 236376 345388 236388
rect 345440 236376 345446 236428
rect 401502 236376 401508 236428
rect 401560 236416 401566 236428
rect 406378 236416 406384 236428
rect 401560 236388 406384 236416
rect 401560 236376 401566 236388
rect 406378 236376 406384 236388
rect 406436 236376 406442 236428
rect 409046 236376 409052 236428
rect 409104 236416 409110 236428
rect 563146 236416 563152 236428
rect 409104 236388 563152 236416
rect 409104 236376 409110 236388
rect 563146 236376 563152 236388
rect 563204 236376 563210 236428
rect 216732 236320 253336 236348
rect 216732 236308 216738 236320
rect 260834 236308 260840 236360
rect 260892 236348 260898 236360
rect 278866 236348 278872 236360
rect 260892 236320 278872 236348
rect 260892 236308 260898 236320
rect 278866 236308 278872 236320
rect 278924 236308 278930 236360
rect 303522 236308 303528 236360
rect 303580 236348 303586 236360
rect 315022 236348 315028 236360
rect 303580 236320 315028 236348
rect 303580 236308 303586 236320
rect 315022 236308 315028 236320
rect 315080 236308 315086 236360
rect 319162 236308 319168 236360
rect 319220 236348 319226 236360
rect 351086 236348 351092 236360
rect 319220 236320 351092 236348
rect 319220 236308 319226 236320
rect 351086 236308 351092 236320
rect 351144 236308 351150 236360
rect 396166 236308 396172 236360
rect 396224 236348 396230 236360
rect 399294 236348 399300 236360
rect 396224 236320 399300 236348
rect 396224 236308 396230 236320
rect 399294 236308 399300 236320
rect 399352 236308 399358 236360
rect 409322 236308 409328 236360
rect 409380 236348 409386 236360
rect 565538 236348 565544 236360
rect 409380 236320 565544 236348
rect 409380 236308 409386 236320
rect 565538 236308 565544 236320
rect 565596 236308 565602 236360
rect 103422 236240 103428 236292
rect 103480 236280 103486 236292
rect 196894 236280 196900 236292
rect 103480 236252 196900 236280
rect 103480 236240 103486 236252
rect 196894 236240 196900 236252
rect 196952 236240 196958 236292
rect 205726 236240 205732 236292
rect 205784 236280 205790 236292
rect 254302 236280 254308 236292
rect 205784 236252 254308 236280
rect 205784 236240 205790 236252
rect 254302 236240 254308 236252
rect 254360 236240 254366 236292
rect 256510 236240 256516 236292
rect 256568 236280 256574 236292
rect 278498 236280 278504 236292
rect 256568 236252 278504 236280
rect 256568 236240 256574 236252
rect 278498 236240 278504 236252
rect 278556 236240 278562 236292
rect 320634 236240 320640 236292
rect 320692 236280 320698 236292
rect 356422 236280 356428 236292
rect 320692 236252 356428 236280
rect 320692 236240 320698 236252
rect 356422 236240 356428 236252
rect 356480 236240 356486 236292
rect 387610 236240 387616 236292
rect 387668 236280 387674 236292
rect 401502 236280 401508 236292
rect 387668 236252 401508 236280
rect 387668 236240 387674 236252
rect 401502 236240 401508 236252
rect 401560 236240 401566 236292
rect 413370 236240 413376 236292
rect 413428 236280 413434 236292
rect 561582 236280 561588 236292
rect 413428 236252 561588 236280
rect 413428 236240 413434 236252
rect 561582 236240 561588 236252
rect 561640 236240 561646 236292
rect 111702 236172 111708 236224
rect 111760 236212 111766 236224
rect 197170 236212 197176 236224
rect 111760 236184 197176 236212
rect 111760 236172 111766 236184
rect 197170 236172 197176 236184
rect 197228 236172 197234 236224
rect 197262 236172 197268 236224
rect 197320 236212 197326 236224
rect 207198 236212 207204 236224
rect 197320 236184 207204 236212
rect 197320 236172 197326 236184
rect 207198 236172 207204 236184
rect 207256 236172 207262 236224
rect 210970 236172 210976 236224
rect 211028 236212 211034 236224
rect 260006 236212 260012 236224
rect 211028 236184 260012 236212
rect 211028 236172 211034 236184
rect 260006 236172 260012 236184
rect 260064 236172 260070 236224
rect 260742 236172 260748 236224
rect 260800 236212 260806 236224
rect 280338 236212 280344 236224
rect 260800 236184 280344 236212
rect 260800 236172 260806 236184
rect 280338 236172 280344 236184
rect 280396 236172 280402 236224
rect 303798 236172 303804 236224
rect 303856 236212 303862 236224
rect 317966 236212 317972 236224
rect 303856 236184 317972 236212
rect 303856 236172 303862 236184
rect 317966 236172 317972 236184
rect 318024 236172 318030 236224
rect 322014 236172 322020 236224
rect 322072 236212 322078 236224
rect 359182 236212 359188 236224
rect 322072 236184 359188 236212
rect 322072 236172 322078 236184
rect 359182 236172 359188 236184
rect 359240 236172 359246 236224
rect 379422 236172 379428 236224
rect 379480 236212 379486 236224
rect 390370 236212 390376 236224
rect 379480 236184 390376 236212
rect 379480 236172 379486 236184
rect 390370 236172 390376 236184
rect 390428 236172 390434 236224
rect 400766 236172 400772 236224
rect 400824 236212 400830 236224
rect 413278 236212 413284 236224
rect 400824 236184 413284 236212
rect 400824 236172 400830 236184
rect 413278 236172 413284 236184
rect 413336 236172 413342 236224
rect 413554 236172 413560 236224
rect 413612 236212 413618 236224
rect 561674 236212 561680 236224
rect 413612 236184 561680 236212
rect 413612 236172 413618 236184
rect 561674 236172 561680 236184
rect 561732 236172 561738 236224
rect 86862 236104 86868 236156
rect 86920 236144 86926 236156
rect 203334 236144 203340 236156
rect 86920 236116 203340 236144
rect 86920 236104 86926 236116
rect 203334 236104 203340 236116
rect 203392 236104 203398 236156
rect 204162 236104 204168 236156
rect 204220 236144 204226 236156
rect 257154 236144 257160 236156
rect 204220 236116 257160 236144
rect 204220 236104 204226 236116
rect 257154 236104 257160 236116
rect 257212 236104 257218 236156
rect 259362 236104 259368 236156
rect 259420 236144 259426 236156
rect 279234 236144 279240 236156
rect 259420 236116 279240 236144
rect 259420 236104 259426 236116
rect 279234 236104 279240 236116
rect 279292 236104 279298 236156
rect 309226 236104 309232 236156
rect 309284 236144 309290 236156
rect 328638 236144 328644 236156
rect 309284 236116 328644 236144
rect 309284 236104 309290 236116
rect 328638 236104 328644 236116
rect 328696 236104 328702 236156
rect 377950 236104 377956 236156
rect 378008 236144 378014 236156
rect 387610 236144 387616 236156
rect 378008 236116 387616 236144
rect 378008 236104 378014 236116
rect 387610 236104 387616 236116
rect 387668 236104 387674 236156
rect 390830 236104 390836 236156
rect 390888 236144 390894 236156
rect 401594 236144 401600 236156
rect 390888 236116 401600 236144
rect 390888 236104 390894 236116
rect 401594 236104 401600 236116
rect 401652 236104 401658 236156
rect 410058 236104 410064 236156
rect 410116 236144 410122 236156
rect 565814 236144 565820 236156
rect 410116 236116 565820 236144
rect 410116 236104 410122 236116
rect 565814 236104 565820 236116
rect 565872 236104 565878 236156
rect 67542 236036 67548 236088
rect 67600 236076 67606 236088
rect 192938 236076 192944 236088
rect 67600 236048 192944 236076
rect 67600 236036 67606 236048
rect 192938 236036 192944 236048
rect 192996 236036 193002 236088
rect 193030 236036 193036 236088
rect 193088 236076 193094 236088
rect 251818 236076 251824 236088
rect 193088 236048 251824 236076
rect 193088 236036 193094 236048
rect 251818 236036 251824 236048
rect 251876 236036 251882 236088
rect 253750 236036 253756 236088
rect 253808 236076 253814 236088
rect 276382 236076 276388 236088
rect 253808 236048 276388 236076
rect 253808 236036 253814 236048
rect 276382 236036 276388 236048
rect 276440 236036 276446 236088
rect 300946 236036 300952 236088
rect 301004 236076 301010 236088
rect 309410 236076 309416 236088
rect 301004 236048 309416 236076
rect 301004 236036 301010 236048
rect 309410 236036 309416 236048
rect 309468 236036 309474 236088
rect 330570 236036 330576 236088
rect 330628 236076 330634 236088
rect 378502 236076 378508 236088
rect 330628 236048 378508 236076
rect 330628 236036 330634 236048
rect 378502 236036 378508 236048
rect 378560 236036 378566 236088
rect 410426 236036 410432 236088
rect 410484 236076 410490 236088
rect 568022 236076 568028 236088
rect 410484 236048 568028 236076
rect 410484 236036 410490 236048
rect 568022 236036 568028 236048
rect 568080 236036 568086 236088
rect 73154 235968 73160 236020
rect 73212 236008 73218 236020
rect 200114 236008 200120 236020
rect 73212 235980 200120 236008
rect 73212 235968 73218 235980
rect 200114 235968 200120 235980
rect 200172 235968 200178 236020
rect 201402 235968 201408 236020
rect 201460 236008 201466 236020
rect 254670 236008 254676 236020
rect 201460 235980 254676 236008
rect 201460 235968 201466 235980
rect 254670 235968 254676 235980
rect 254728 235968 254734 236020
rect 255406 235968 255412 236020
rect 255464 236008 255470 236020
rect 277118 236008 277124 236020
rect 255464 235980 277124 236008
rect 255464 235968 255470 235980
rect 277118 235968 277124 235980
rect 277176 235968 277182 236020
rect 298094 235968 298100 236020
rect 298152 236008 298158 236020
rect 303798 236008 303804 236020
rect 298152 235980 303804 236008
rect 298152 235968 298158 235980
rect 303798 235968 303804 235980
rect 303856 235968 303862 236020
rect 313458 235968 313464 236020
rect 313516 236008 313522 236020
rect 337102 236008 337108 236020
rect 313516 235980 337108 236008
rect 313516 235968 313522 235980
rect 337102 235968 337108 235980
rect 337160 235968 337166 236020
rect 338390 235968 338396 236020
rect 338448 236008 338454 236020
rect 395154 236008 395160 236020
rect 338448 235980 395160 236008
rect 338448 235968 338454 235980
rect 395154 235968 395160 235980
rect 395212 235968 395218 236020
rect 410794 235968 410800 236020
rect 410852 236008 410858 236020
rect 569954 236008 569960 236020
rect 410852 235980 569960 236008
rect 410852 235968 410858 235980
rect 569954 235968 569960 235980
rect 570012 235968 570018 236020
rect 168098 235900 168104 235952
rect 168156 235940 168162 235952
rect 241146 235940 241152 235952
rect 168156 235912 241152 235940
rect 168156 235900 168162 235912
rect 241146 235900 241152 235912
rect 241204 235900 241210 235952
rect 245562 235900 245568 235952
rect 245620 235940 245626 235952
rect 245620 235900 245654 235940
rect 248322 235900 248328 235952
rect 248380 235940 248386 235952
rect 273898 235940 273904 235952
rect 248380 235912 273904 235940
rect 248380 235900 248386 235912
rect 273898 235900 273904 235912
rect 273956 235900 273962 235952
rect 310606 235900 310612 235952
rect 310664 235940 310670 235952
rect 331766 235940 331772 235952
rect 310664 235912 331772 235940
rect 310664 235900 310670 235912
rect 331766 235900 331772 235912
rect 331824 235900 331830 235952
rect 334526 235900 334532 235952
rect 334584 235940 334590 235952
rect 346486 235940 346492 235952
rect 334584 235912 346492 235940
rect 334584 235900 334590 235912
rect 346486 235900 346492 235912
rect 346544 235900 346550 235952
rect 397638 235900 397644 235952
rect 397696 235940 397702 235952
rect 536742 235940 536748 235952
rect 397696 235912 536748 235940
rect 397696 235900 397702 235912
rect 536742 235900 536748 235912
rect 536800 235900 536806 235952
rect 165338 235832 165344 235884
rect 165396 235872 165402 235884
rect 239766 235872 239772 235884
rect 165396 235844 239772 235872
rect 165396 235832 165402 235844
rect 239766 235832 239772 235844
rect 239824 235832 239830 235884
rect 245626 235872 245654 235900
rect 272426 235872 272432 235884
rect 245626 235844 272432 235872
rect 272426 235832 272432 235844
rect 272484 235832 272490 235884
rect 299934 235832 299940 235884
rect 299992 235872 299998 235884
rect 304074 235872 304080 235884
rect 299992 235844 304080 235872
rect 299992 235832 299998 235844
rect 304074 235832 304080 235844
rect 304132 235832 304138 235884
rect 393314 235832 393320 235884
rect 393372 235872 393378 235884
rect 528462 235872 528468 235884
rect 393372 235844 528468 235872
rect 393372 235832 393378 235844
rect 528462 235832 528468 235844
rect 528520 235832 528526 235884
rect 173710 235764 173716 235816
rect 173768 235804 173774 235816
rect 244274 235804 244280 235816
rect 173768 235776 244280 235804
rect 173768 235764 173774 235776
rect 244274 235764 244280 235776
rect 244332 235764 244338 235816
rect 250990 235764 250996 235816
rect 251048 235804 251054 235816
rect 275278 235804 275284 235816
rect 251048 235776 275284 235804
rect 251048 235764 251054 235776
rect 275278 235764 275284 235776
rect 275336 235764 275342 235816
rect 395062 235764 395068 235816
rect 395120 235804 395126 235816
rect 529934 235804 529940 235816
rect 395120 235776 529940 235804
rect 395120 235764 395126 235776
rect 529934 235764 529940 235776
rect 529992 235764 529998 235816
rect 173802 235696 173808 235748
rect 173860 235736 173866 235748
rect 243262 235736 243268 235748
rect 173860 235708 243268 235736
rect 173860 235696 173866 235708
rect 243262 235696 243268 235708
rect 243320 235696 243326 235748
rect 247310 235696 247316 235748
rect 247368 235736 247374 235748
rect 261386 235736 261392 235748
rect 247368 235708 261392 235736
rect 247368 235696 247374 235708
rect 261386 235696 261392 235708
rect 261444 235696 261450 235748
rect 267182 235696 267188 235748
rect 267240 235736 267246 235748
rect 281350 235736 281356 235748
rect 267240 235708 281356 235736
rect 267240 235696 267246 235708
rect 281350 235696 281356 235708
rect 281408 235696 281414 235748
rect 299198 235696 299204 235748
rect 299256 235736 299262 235748
rect 303706 235736 303712 235748
rect 299256 235708 303712 235736
rect 299256 235696 299262 235708
rect 303706 235696 303712 235708
rect 303764 235696 303770 235748
rect 307294 235736 307300 235748
rect 305472 235708 307300 235736
rect 197262 235628 197268 235680
rect 197320 235668 197326 235680
rect 246114 235668 246120 235680
rect 197320 235640 246120 235668
rect 197320 235628 197326 235640
rect 246114 235628 246120 235640
rect 246172 235628 246178 235680
rect 251082 235628 251088 235680
rect 251140 235668 251146 235680
rect 275002 235668 275008 235680
rect 251140 235640 275008 235668
rect 251140 235628 251146 235640
rect 275002 235628 275008 235640
rect 275060 235628 275066 235680
rect 301314 235628 301320 235680
rect 301372 235668 301378 235680
rect 305472 235668 305500 235708
rect 307294 235696 307300 235708
rect 307352 235696 307358 235748
rect 392946 235696 392952 235748
rect 393004 235736 393010 235748
rect 524414 235736 524420 235748
rect 393004 235708 524420 235736
rect 393004 235696 393010 235708
rect 524414 235696 524420 235708
rect 524472 235696 524478 235748
rect 301372 235640 305500 235668
rect 301372 235628 301378 235640
rect 306650 235628 306656 235680
rect 306708 235668 306714 235680
rect 308766 235668 308772 235680
rect 306708 235640 308772 235668
rect 306708 235628 306714 235640
rect 308766 235628 308772 235640
rect 308824 235628 308830 235680
rect 401594 235628 401600 235680
rect 401652 235668 401658 235680
rect 520182 235668 520188 235680
rect 401652 235640 520188 235668
rect 401652 235628 401658 235640
rect 520182 235628 520188 235640
rect 520240 235628 520246 235680
rect 158622 235560 158628 235612
rect 158680 235600 158686 235612
rect 208118 235600 208124 235612
rect 158680 235572 208124 235600
rect 158680 235560 158686 235572
rect 208118 235560 208124 235572
rect 208176 235560 208182 235612
rect 222930 235600 222936 235612
rect 208320 235572 222936 235600
rect 155954 235492 155960 235544
rect 156012 235532 156018 235544
rect 208320 235532 208348 235572
rect 222930 235560 222936 235572
rect 222988 235560 222994 235612
rect 224034 235560 224040 235612
rect 224092 235600 224098 235612
rect 224678 235600 224684 235612
rect 224092 235572 224684 235600
rect 224092 235560 224098 235572
rect 224678 235560 224684 235572
rect 224736 235560 224742 235612
rect 247126 235600 247132 235612
rect 233344 235572 247132 235600
rect 223298 235532 223304 235544
rect 156012 235504 208348 235532
rect 218026 235504 223304 235532
rect 156012 235492 156018 235504
rect 161566 235424 161572 235476
rect 161624 235464 161630 235476
rect 208210 235464 208216 235476
rect 161624 235436 208216 235464
rect 161624 235424 161630 235436
rect 208210 235424 208216 235436
rect 208268 235424 208274 235476
rect 218026 235464 218054 235504
rect 223298 235492 223304 235504
rect 223356 235492 223362 235544
rect 208320 235436 218054 235464
rect 42150 235356 42156 235408
rect 42208 235396 42214 235408
rect 42794 235396 42800 235408
rect 42208 235368 42800 235396
rect 42208 235356 42214 235368
rect 42794 235356 42800 235368
rect 42852 235356 42858 235408
rect 156046 235356 156052 235408
rect 156104 235396 156110 235408
rect 208320 235396 208348 235436
rect 156104 235368 208348 235396
rect 156104 235356 156110 235368
rect 208394 235356 208400 235408
rect 208452 235396 208458 235408
rect 231486 235396 231492 235408
rect 208452 235368 231492 235396
rect 208452 235356 208458 235368
rect 231486 235356 231492 235368
rect 231544 235356 231550 235408
rect 183462 235288 183468 235340
rect 183520 235328 183526 235340
rect 233344 235328 233372 235572
rect 247126 235560 247132 235572
rect 247184 235560 247190 235612
rect 259638 235600 259644 235612
rect 252664 235572 259644 235600
rect 244274 235492 244280 235544
rect 244332 235532 244338 235544
rect 249978 235532 249984 235544
rect 244332 235504 249984 235532
rect 244332 235492 244338 235504
rect 249978 235492 249984 235504
rect 250036 235492 250042 235544
rect 236086 235424 236092 235476
rect 236144 235464 236150 235476
rect 252664 235464 252692 235572
rect 259638 235560 259644 235572
rect 259696 235560 259702 235612
rect 261938 235560 261944 235612
rect 261996 235600 262002 235612
rect 279602 235600 279608 235612
rect 261996 235572 279608 235600
rect 261996 235560 262002 235572
rect 279602 235560 279608 235572
rect 279660 235560 279666 235612
rect 299566 235560 299572 235612
rect 299624 235600 299630 235612
rect 307202 235600 307208 235612
rect 299624 235572 307208 235600
rect 299624 235560 299630 235572
rect 307202 235560 307208 235572
rect 307260 235560 307266 235612
rect 331674 235560 331680 235612
rect 331732 235600 331738 235612
rect 346394 235600 346400 235612
rect 331732 235572 346400 235600
rect 331732 235560 331738 235572
rect 346394 235560 346400 235572
rect 346452 235560 346458 235612
rect 386230 235560 386236 235612
rect 386288 235600 386294 235612
rect 393774 235600 393780 235612
rect 386288 235572 393780 235600
rect 386288 235560 386294 235572
rect 393774 235560 393780 235572
rect 393832 235560 393838 235612
rect 393958 235560 393964 235612
rect 394016 235600 394022 235612
rect 511994 235600 512000 235612
rect 394016 235572 512000 235600
rect 394016 235560 394022 235572
rect 511994 235560 512000 235572
rect 512052 235560 512058 235612
rect 674742 235560 674748 235612
rect 674800 235600 674806 235612
rect 675662 235600 675668 235612
rect 674800 235572 675668 235600
rect 674800 235560 674806 235572
rect 675662 235560 675668 235572
rect 675720 235560 675726 235612
rect 258166 235492 258172 235544
rect 258224 235532 258230 235544
rect 276014 235532 276020 235544
rect 258224 235504 276020 235532
rect 258224 235492 258230 235504
rect 276014 235492 276020 235504
rect 276072 235492 276078 235544
rect 300302 235492 300308 235544
rect 300360 235532 300366 235544
rect 306650 235532 306656 235544
rect 300360 235504 306656 235532
rect 300360 235492 300366 235504
rect 306650 235492 306656 235504
rect 306708 235492 306714 235544
rect 394050 235492 394056 235544
rect 394108 235532 394114 235544
rect 401410 235532 401416 235544
rect 394108 235504 401416 235532
rect 394108 235492 394114 235504
rect 401410 235492 401416 235504
rect 401468 235492 401474 235544
rect 401502 235492 401508 235544
rect 401560 235532 401566 235544
rect 513466 235532 513472 235544
rect 401560 235504 513472 235532
rect 401560 235492 401566 235504
rect 513466 235492 513472 235504
rect 513524 235492 513530 235544
rect 674650 235492 674656 235544
rect 674708 235532 674714 235544
rect 675754 235532 675760 235544
rect 674708 235504 675760 235532
rect 674708 235492 674714 235504
rect 675754 235492 675760 235504
rect 675812 235492 675818 235544
rect 236144 235436 252692 235464
rect 236144 235424 236150 235436
rect 256602 235424 256608 235476
rect 256660 235464 256666 235476
rect 277854 235464 277860 235476
rect 256660 235436 277860 235464
rect 256660 235424 256666 235436
rect 277854 235424 277860 235436
rect 277912 235424 277918 235476
rect 388714 235424 388720 235476
rect 388772 235464 388778 235476
rect 511902 235464 511908 235476
rect 388772 235436 511908 235464
rect 388772 235424 388778 235436
rect 511902 235424 511908 235436
rect 511960 235424 511966 235476
rect 233418 235356 233424 235408
rect 233476 235396 233482 235408
rect 233476 235368 236224 235396
rect 233476 235356 233482 235368
rect 183520 235300 233372 235328
rect 236196 235328 236224 235368
rect 244182 235356 244188 235408
rect 244240 235396 244246 235408
rect 245746 235396 245752 235408
rect 244240 235368 245752 235396
rect 244240 235356 244246 235368
rect 245746 235356 245752 235368
rect 245804 235356 245810 235408
rect 255314 235356 255320 235408
rect 255372 235396 255378 235408
rect 274266 235396 274272 235408
rect 255372 235368 274272 235396
rect 255372 235356 255378 235368
rect 274266 235356 274272 235368
rect 274324 235356 274330 235408
rect 333054 235356 333060 235408
rect 333112 235396 333118 235408
rect 346210 235396 346216 235408
rect 333112 235368 346216 235396
rect 333112 235356 333118 235368
rect 346210 235356 346216 235368
rect 346268 235356 346274 235408
rect 385494 235356 385500 235408
rect 385552 235396 385558 235408
rect 507946 235396 507952 235408
rect 385552 235368 507952 235396
rect 385552 235356 385558 235368
rect 507946 235356 507952 235368
rect 508004 235356 508010 235408
rect 236196 235300 251588 235328
rect 183520 235288 183526 235300
rect 190362 235220 190368 235272
rect 190420 235260 190426 235272
rect 251450 235260 251456 235272
rect 190420 235232 251456 235260
rect 190420 235220 190426 235232
rect 251450 235220 251456 235232
rect 251508 235220 251514 235272
rect 251560 235260 251588 235300
rect 255222 235288 255228 235340
rect 255280 235328 255286 235340
rect 275646 235328 275652 235340
rect 255280 235300 275652 235328
rect 255280 235288 255286 235300
rect 275646 235288 275652 235300
rect 275704 235288 275710 235340
rect 306374 235288 306380 235340
rect 306432 235328 306438 235340
rect 321002 235328 321008 235340
rect 306432 235300 321008 235328
rect 306432 235288 306438 235300
rect 321002 235288 321008 235300
rect 321060 235288 321066 235340
rect 384022 235288 384028 235340
rect 384080 235328 384086 235340
rect 506382 235328 506388 235340
rect 384080 235300 506388 235328
rect 384080 235288 384086 235300
rect 506382 235288 506388 235300
rect 506440 235288 506446 235340
rect 256786 235260 256792 235272
rect 251560 235232 256792 235260
rect 256786 235220 256792 235232
rect 256844 235220 256850 235272
rect 262030 235220 262036 235272
rect 262088 235260 262094 235272
rect 267182 235260 267188 235272
rect 262088 235232 267188 235260
rect 262088 235220 262094 235232
rect 267182 235220 267188 235232
rect 267240 235220 267246 235272
rect 267274 235220 267280 235272
rect 267332 235260 267338 235272
rect 280706 235260 280712 235272
rect 267332 235232 280712 235260
rect 267332 235220 267338 235232
rect 280706 235220 280712 235232
rect 280764 235220 280770 235272
rect 304902 235220 304908 235272
rect 304960 235260 304966 235272
rect 317874 235260 317880 235272
rect 304960 235232 317880 235260
rect 304960 235220 304966 235232
rect 317874 235220 317880 235232
rect 317932 235220 317938 235272
rect 383378 235220 383384 235272
rect 383436 235260 383442 235272
rect 502794 235260 502800 235272
rect 383436 235232 502800 235260
rect 383436 235220 383442 235232
rect 502794 235220 502800 235232
rect 502852 235220 502858 235272
rect 187602 235152 187608 235204
rect 187660 235192 187666 235204
rect 187660 235164 235948 235192
rect 187660 235152 187666 235164
rect 169662 235084 169668 235136
rect 169720 235124 169726 235136
rect 208394 235124 208400 235136
rect 169720 235096 208400 235124
rect 169720 235084 169726 235096
rect 208394 235084 208400 235096
rect 208452 235084 208458 235136
rect 179322 235016 179328 235068
rect 179380 235056 179386 235068
rect 197262 235056 197268 235068
rect 179380 235028 197268 235056
rect 179380 235016 179386 235028
rect 197262 235016 197268 235028
rect 197320 235016 197326 235068
rect 235920 235056 235948 235164
rect 236270 235152 236276 235204
rect 236328 235192 236334 235204
rect 253934 235192 253940 235204
rect 236328 235164 253940 235192
rect 236328 235152 236334 235164
rect 253934 235152 253940 235164
rect 253992 235152 253998 235204
rect 259178 235152 259184 235204
rect 259236 235192 259242 235204
rect 278130 235192 278136 235204
rect 259236 235164 278136 235192
rect 259236 235152 259242 235164
rect 278130 235152 278136 235164
rect 278188 235152 278194 235204
rect 306006 235152 306012 235204
rect 306064 235192 306070 235204
rect 317782 235192 317788 235204
rect 306064 235164 317788 235192
rect 306064 235152 306070 235164
rect 317782 235152 317788 235164
rect 317840 235152 317846 235204
rect 381906 235152 381912 235204
rect 381964 235192 381970 235204
rect 500862 235192 500868 235204
rect 381964 235164 500868 235192
rect 381964 235152 381970 235164
rect 500862 235152 500868 235164
rect 500920 235152 500926 235204
rect 235994 235084 236000 235136
rect 236052 235124 236058 235136
rect 246942 235124 246948 235136
rect 236052 235096 246948 235124
rect 236052 235084 236058 235096
rect 246942 235084 246948 235096
rect 247000 235084 247006 235136
rect 247126 235084 247132 235136
rect 247184 235124 247190 235136
rect 258534 235124 258540 235136
rect 247184 235096 258540 235124
rect 247184 235084 247190 235096
rect 258534 235084 258540 235096
rect 258592 235084 258598 235136
rect 262122 235084 262128 235136
rect 262180 235124 262186 235136
rect 267274 235124 267280 235136
rect 262180 235096 267280 235124
rect 262180 235084 262186 235096
rect 267274 235084 267280 235096
rect 267332 235084 267338 235136
rect 267366 235084 267372 235136
rect 267424 235124 267430 235136
rect 276750 235124 276756 235136
rect 267424 235096 276756 235124
rect 267424 235084 267430 235096
rect 276750 235084 276756 235096
rect 276808 235084 276814 235136
rect 305638 235084 305644 235136
rect 305696 235124 305702 235136
rect 317690 235124 317696 235136
rect 305696 235096 317696 235124
rect 305696 235084 305702 235096
rect 317690 235084 317696 235096
rect 317748 235084 317754 235136
rect 379054 235084 379060 235136
rect 379112 235124 379118 235136
rect 495342 235124 495348 235136
rect 379112 235096 495348 235124
rect 379112 235084 379118 235096
rect 495342 235084 495348 235096
rect 495400 235084 495406 235136
rect 248966 235056 248972 235068
rect 197372 235028 226334 235056
rect 235920 235028 248972 235056
rect 161474 234948 161480 235000
rect 161532 234988 161538 235000
rect 161532 234960 168374 234988
rect 161532 234948 161538 234960
rect 168346 234852 168374 234960
rect 193030 234880 193036 234932
rect 193088 234920 193094 234932
rect 197372 234920 197400 235028
rect 193088 234892 197400 234920
rect 197464 234960 205956 234988
rect 193088 234880 193094 234892
rect 197464 234852 197492 234960
rect 198642 234880 198648 234932
rect 198700 234920 198706 234932
rect 205726 234920 205732 234932
rect 198700 234892 205732 234920
rect 198700 234880 198706 234892
rect 205726 234880 205732 234892
rect 205784 234880 205790 234932
rect 205928 234920 205956 234960
rect 208118 234948 208124 235000
rect 208176 234988 208182 235000
rect 225782 234988 225788 235000
rect 208176 234960 225788 234988
rect 208176 234948 208182 234960
rect 225782 234948 225788 234960
rect 225840 234948 225846 235000
rect 226306 234988 226334 235028
rect 248966 235016 248972 235028
rect 249024 235016 249030 235068
rect 257982 235016 257988 235068
rect 258040 235056 258046 235068
rect 274634 235056 274640 235068
rect 258040 235028 274640 235056
rect 258040 235016 258046 235028
rect 274634 235016 274640 235028
rect 274692 235016 274698 235068
rect 300670 235016 300676 235068
rect 300728 235056 300734 235068
rect 306742 235056 306748 235068
rect 300728 235028 306748 235056
rect 300728 235016 300734 235028
rect 306742 235016 306748 235028
rect 306800 235016 306806 235068
rect 307018 235016 307024 235068
rect 307076 235056 307082 235068
rect 320818 235056 320824 235068
rect 307076 235028 320824 235056
rect 307076 235016 307082 235028
rect 320818 235016 320824 235028
rect 320876 235016 320882 235068
rect 328822 235016 328828 235068
rect 328880 235056 328886 235068
rect 343634 235056 343640 235068
rect 328880 235028 343640 235056
rect 328880 235016 328886 235028
rect 343634 235016 343640 235028
rect 343692 235016 343698 235068
rect 380802 235016 380808 235068
rect 380860 235056 380866 235068
rect 489822 235056 489828 235068
rect 380860 235028 489828 235056
rect 380860 235016 380866 235028
rect 489822 235016 489828 235028
rect 489880 235016 489886 235068
rect 250806 234988 250812 235000
rect 226306 234960 250812 234988
rect 250806 234948 250812 234960
rect 250864 234948 250870 235000
rect 263502 234948 263508 235000
rect 263560 234988 263566 235000
rect 267458 234988 267464 235000
rect 263560 234960 267464 234988
rect 263560 234948 263566 234960
rect 267458 234948 267464 234960
rect 267516 234948 267522 235000
rect 304166 234948 304172 235000
rect 304224 234988 304230 235000
rect 315390 234988 315396 235000
rect 304224 234960 315396 234988
rect 304224 234948 304230 234960
rect 315390 234948 315396 234960
rect 315448 234948 315454 235000
rect 323118 234948 323124 235000
rect 323176 234988 323182 235000
rect 340782 234988 340788 235000
rect 323176 234960 340788 234988
rect 323176 234948 323182 234960
rect 340782 234948 340788 234960
rect 340840 234948 340846 235000
rect 376570 234948 376576 235000
rect 376628 234988 376634 235000
rect 481542 234988 481548 235000
rect 376628 234960 481548 234988
rect 376628 234948 376634 234960
rect 481542 234948 481548 234960
rect 481600 234948 481606 235000
rect 212902 234920 212908 234932
rect 205928 234892 212908 234920
rect 212902 234880 212908 234892
rect 212960 234880 212966 234932
rect 233142 234880 233148 234932
rect 233200 234920 233206 234932
rect 236270 234920 236276 234932
rect 233200 234892 236276 234920
rect 233200 234880 233206 234892
rect 236270 234880 236276 234892
rect 236328 234880 236334 234932
rect 249610 234920 249616 234932
rect 245626 234892 249616 234920
rect 168346 234824 197492 234852
rect 233234 234812 233240 234864
rect 233292 234852 233298 234864
rect 245626 234852 245654 234892
rect 249610 234880 249616 234892
rect 249668 234880 249674 234932
rect 255498 234880 255504 234932
rect 255556 234920 255562 234932
rect 273162 234920 273168 234932
rect 255556 234892 273168 234920
rect 255556 234880 255562 234892
rect 273162 234880 273168 234892
rect 273220 234880 273226 234932
rect 304534 234880 304540 234932
rect 304592 234920 304598 234932
rect 315298 234920 315304 234932
rect 304592 234892 315304 234920
rect 304592 234880 304598 234892
rect 315298 234880 315304 234892
rect 315356 234880 315362 234932
rect 336274 234880 336280 234932
rect 336332 234920 336338 234932
rect 336642 234920 336648 234932
rect 336332 234892 336648 234920
rect 336332 234880 336338 234892
rect 336642 234880 336648 234892
rect 336700 234880 336706 234932
rect 347038 234880 347044 234932
rect 347096 234920 347102 234932
rect 347682 234920 347688 234932
rect 347096 234892 347688 234920
rect 347096 234880 347102 234892
rect 347682 234880 347688 234892
rect 347740 234880 347746 234932
rect 402606 234880 402612 234932
rect 402664 234920 402670 234932
rect 413738 234920 413744 234932
rect 402664 234892 413744 234920
rect 402664 234880 402670 234892
rect 413738 234880 413744 234892
rect 413796 234880 413802 234932
rect 233292 234824 245654 234852
rect 233292 234812 233298 234824
rect 247034 234812 247040 234864
rect 247092 234852 247098 234864
rect 255682 234852 255688 234864
rect 247092 234824 255688 234852
rect 247092 234812 247098 234824
rect 255682 234812 255688 234824
rect 255740 234812 255746 234864
rect 272794 234852 272800 234864
rect 267384 234824 272800 234852
rect 210418 234784 210424 234796
rect 198706 234756 210424 234784
rect 197170 234676 197176 234728
rect 197228 234716 197234 234728
rect 198706 234716 198734 234756
rect 210418 234744 210424 234756
rect 210476 234744 210482 234796
rect 212534 234744 212540 234796
rect 212592 234784 212598 234796
rect 217226 234784 217232 234796
rect 212592 234756 217232 234784
rect 212592 234744 212598 234756
rect 217226 234744 217232 234756
rect 217284 234744 217290 234796
rect 246942 234744 246948 234796
rect 247000 234784 247006 234796
rect 247000 234756 248736 234784
rect 247000 234744 247006 234756
rect 197228 234688 198734 234716
rect 197228 234676 197234 234688
rect 208210 234676 208216 234728
rect 208268 234716 208274 234728
rect 228634 234716 228640 234728
rect 208268 234688 228640 234716
rect 208268 234676 208274 234688
rect 228634 234676 228640 234688
rect 228692 234676 228698 234728
rect 244458 234676 244464 234728
rect 244516 234716 244522 234728
rect 248598 234716 248604 234728
rect 244516 234688 248604 234716
rect 244516 234676 244522 234688
rect 248598 234676 248604 234688
rect 248656 234676 248662 234728
rect 248708 234716 248736 234756
rect 252554 234744 252560 234796
rect 252612 234784 252618 234796
rect 267384 234784 267412 234824
rect 272794 234812 272800 234824
rect 272852 234812 272858 234864
rect 297818 234812 297824 234864
rect 297876 234852 297882 234864
rect 300854 234852 300860 234864
rect 297876 234824 300860 234852
rect 297876 234812 297882 234824
rect 300854 234812 300860 234824
rect 300912 234812 300918 234864
rect 309502 234812 309508 234864
rect 309560 234852 309566 234864
rect 311710 234852 311716 234864
rect 309560 234824 311716 234852
rect 309560 234812 309566 234824
rect 311710 234812 311716 234824
rect 311768 234812 311774 234864
rect 312354 234812 312360 234864
rect 312412 234852 312418 234864
rect 314010 234852 314016 234864
rect 312412 234824 314016 234852
rect 312412 234812 312418 234824
rect 314010 234812 314016 234824
rect 314068 234812 314074 234864
rect 315206 234812 315212 234864
rect 315264 234852 315270 234864
rect 317138 234852 317144 234864
rect 315264 234824 317144 234852
rect 315264 234812 315270 234824
rect 317138 234812 317144 234824
rect 317196 234812 317202 234864
rect 320910 234812 320916 234864
rect 320968 234852 320974 234864
rect 322842 234852 322848 234864
rect 320968 234824 322848 234852
rect 320968 234812 320974 234824
rect 322842 234812 322848 234824
rect 322900 234812 322906 234864
rect 324130 234812 324136 234864
rect 324188 234852 324194 234864
rect 325510 234852 325516 234864
rect 324188 234824 325516 234852
rect 324188 234812 324194 234824
rect 325510 234812 325516 234824
rect 325568 234812 325574 234864
rect 326338 234812 326344 234864
rect 326396 234852 326402 234864
rect 328178 234852 328184 234864
rect 326396 234824 328184 234852
rect 326396 234812 326402 234824
rect 328178 234812 328184 234824
rect 328236 234812 328242 234864
rect 328454 234812 328460 234864
rect 328512 234852 328518 234864
rect 330846 234852 330852 234864
rect 328512 234824 330852 234852
rect 328512 234812 328518 234824
rect 330846 234812 330852 234824
rect 330904 234812 330910 234864
rect 331306 234812 331312 234864
rect 331364 234852 331370 234864
rect 333790 234852 333796 234864
rect 331364 234824 333796 234852
rect 331364 234812 331370 234824
rect 333790 234812 333796 234824
rect 333848 234812 333854 234864
rect 343082 234812 343088 234864
rect 343140 234852 343146 234864
rect 349062 234852 349068 234864
rect 343140 234824 349068 234852
rect 343140 234812 343146 234824
rect 349062 234812 349068 234824
rect 349120 234812 349126 234864
rect 386506 234812 386512 234864
rect 386564 234852 386570 234864
rect 390554 234852 390560 234864
rect 386564 234824 390560 234852
rect 386564 234812 386570 234824
rect 390554 234812 390560 234824
rect 390612 234812 390618 234864
rect 252612 234756 267412 234784
rect 252612 234744 252618 234756
rect 267458 234744 267464 234796
rect 267516 234784 267522 234796
rect 283190 234784 283196 234796
rect 267516 234756 283196 234784
rect 267516 234744 267522 234756
rect 283190 234744 283196 234756
rect 283248 234744 283254 234796
rect 296346 234744 296352 234796
rect 296404 234784 296410 234796
rect 298186 234784 298192 234796
rect 296404 234756 298192 234784
rect 296404 234744 296410 234756
rect 298186 234744 298192 234756
rect 298244 234744 298250 234796
rect 307386 234744 307392 234796
rect 307444 234784 307450 234796
rect 308950 234784 308956 234796
rect 307444 234756 308956 234784
rect 307444 234744 307450 234756
rect 308950 234744 308956 234756
rect 309008 234744 309014 234796
rect 309870 234744 309876 234796
rect 309928 234784 309934 234796
rect 311802 234784 311808 234796
rect 309928 234756 311808 234784
rect 309928 234744 309934 234756
rect 311802 234744 311808 234756
rect 311860 234744 311866 234796
rect 313090 234744 313096 234796
rect 313148 234784 313154 234796
rect 314470 234784 314476 234796
rect 313148 234756 314476 234784
rect 313148 234744 313154 234756
rect 314470 234744 314476 234756
rect 314528 234744 314534 234796
rect 315942 234744 315948 234796
rect 316000 234784 316006 234796
rect 317322 234784 317328 234796
rect 316000 234756 317328 234784
rect 316000 234744 316006 234756
rect 317322 234744 317328 234756
rect 317380 234744 317386 234796
rect 318058 234744 318064 234796
rect 318116 234784 318122 234796
rect 320082 234784 320088 234796
rect 318116 234756 320088 234784
rect 318116 234744 318122 234756
rect 320082 234744 320088 234756
rect 320140 234744 320146 234796
rect 321646 234744 321652 234796
rect 321704 234784 321710 234796
rect 322750 234784 322756 234796
rect 321704 234756 322756 234784
rect 321704 234744 321710 234756
rect 322750 234744 322756 234756
rect 322808 234744 322814 234796
rect 324866 234744 324872 234796
rect 324924 234784 324930 234796
rect 325602 234784 325608 234796
rect 324924 234756 325608 234784
rect 324924 234744 324930 234756
rect 325602 234744 325608 234756
rect 325660 234744 325666 234796
rect 326982 234744 326988 234796
rect 327040 234784 327046 234796
rect 328270 234784 328276 234796
rect 327040 234756 328276 234784
rect 327040 234744 327046 234756
rect 328270 234744 328276 234756
rect 328328 234744 328334 234796
rect 329466 234744 329472 234796
rect 329524 234784 329530 234796
rect 331122 234784 331128 234796
rect 329524 234756 331128 234784
rect 329524 234744 329530 234756
rect 331122 234744 331128 234756
rect 331180 234744 331186 234796
rect 332686 234744 332692 234796
rect 332744 234784 332750 234796
rect 333882 234784 333888 234796
rect 332744 234756 333888 234784
rect 332744 234744 332750 234756
rect 333882 234744 333888 234756
rect 333940 234744 333946 234796
rect 337010 234744 337016 234796
rect 337068 234784 337074 234796
rect 339218 234784 339224 234796
rect 337068 234756 339224 234784
rect 337068 234744 337074 234756
rect 339218 234744 339224 234756
rect 339276 234744 339282 234796
rect 339494 234744 339500 234796
rect 339552 234784 339558 234796
rect 341794 234784 341800 234796
rect 339552 234756 341800 234784
rect 339552 234744 339558 234756
rect 341794 234744 341800 234756
rect 341852 234744 341858 234796
rect 342346 234744 342352 234796
rect 342404 234784 342410 234796
rect 344370 234784 344376 234796
rect 342404 234756 344376 234784
rect 342404 234744 342410 234756
rect 344370 234744 344376 234756
rect 344428 234744 344434 234796
rect 345198 234744 345204 234796
rect 345256 234784 345262 234796
rect 347130 234784 347136 234796
rect 345256 234756 347136 234784
rect 345256 234744 345262 234756
rect 347130 234744 347136 234756
rect 347188 234744 347194 234796
rect 347314 234744 347320 234796
rect 347372 234784 347378 234796
rect 347682 234784 347688 234796
rect 347372 234756 347688 234784
rect 347372 234744 347378 234756
rect 347682 234744 347688 234756
rect 347740 234744 347746 234796
rect 348050 234744 348056 234796
rect 348108 234784 348114 234796
rect 349890 234784 349896 234796
rect 348108 234756 349896 234784
rect 348108 234744 348114 234756
rect 349890 234744 349896 234756
rect 349948 234744 349954 234796
rect 350902 234744 350908 234796
rect 350960 234784 350966 234796
rect 353018 234784 353024 234796
rect 350960 234756 353024 234784
rect 350960 234744 350966 234756
rect 353018 234744 353024 234756
rect 353076 234744 353082 234796
rect 353386 234744 353392 234796
rect 353444 234784 353450 234796
rect 355778 234784 355784 234796
rect 353444 234756 355784 234784
rect 353444 234744 353450 234756
rect 355778 234744 355784 234756
rect 355836 234744 355842 234796
rect 356238 234744 356244 234796
rect 356296 234784 356302 234796
rect 358538 234784 358544 234796
rect 356296 234756 358544 234784
rect 356296 234744 356302 234756
rect 358538 234744 358544 234756
rect 358596 234744 358602 234796
rect 359090 234744 359096 234796
rect 359148 234784 359154 234796
rect 361206 234784 361212 234796
rect 359148 234756 361212 234784
rect 359148 234744 359154 234756
rect 361206 234744 361212 234756
rect 361264 234744 361270 234796
rect 384390 234744 384396 234796
rect 384448 234784 384454 234796
rect 387794 234784 387800 234796
rect 384448 234756 387800 234784
rect 384448 234744 384454 234756
rect 387794 234744 387800 234756
rect 387852 234744 387858 234796
rect 248708 234688 252968 234716
rect 42150 234608 42156 234660
rect 42208 234648 42214 234660
rect 43254 234648 43260 234660
rect 42208 234620 43260 234648
rect 42208 234608 42214 234620
rect 43254 234608 43260 234620
rect 43312 234608 43318 234660
rect 215294 234608 215300 234660
rect 215352 234648 215358 234660
rect 220078 234648 220084 234660
rect 215352 234620 220084 234648
rect 215352 234608 215358 234620
rect 220078 234608 220084 234620
rect 220136 234608 220142 234660
rect 241790 234608 241796 234660
rect 241848 234648 241854 234660
rect 242894 234648 242900 234660
rect 241848 234620 242900 234648
rect 241848 234608 241854 234620
rect 242894 234608 242900 234620
rect 242952 234608 242958 234660
rect 246942 234608 246948 234660
rect 247000 234648 247006 234660
rect 252830 234648 252836 234660
rect 247000 234620 252836 234648
rect 247000 234608 247006 234620
rect 252830 234608 252836 234620
rect 252888 234608 252894 234660
rect 252940 234648 252968 234688
rect 253842 234676 253848 234728
rect 253900 234716 253906 234728
rect 267366 234716 267372 234728
rect 253900 234688 267372 234716
rect 253900 234676 253906 234688
rect 267366 234676 267372 234688
rect 267424 234676 267430 234728
rect 267550 234676 267556 234728
rect 267608 234716 267614 234728
rect 282454 234716 282460 234728
rect 267608 234688 282460 234716
rect 267608 234676 267614 234688
rect 282454 234676 282460 234688
rect 282512 234676 282518 234728
rect 292574 234676 292580 234728
rect 292632 234716 292638 234728
rect 294598 234716 294604 234728
rect 292632 234688 294604 234716
rect 292632 234676 292638 234688
rect 294598 234676 294604 234688
rect 294656 234676 294662 234728
rect 295242 234676 295248 234728
rect 295300 234716 295306 234728
rect 295886 234716 295892 234728
rect 295300 234688 295892 234716
rect 295300 234676 295306 234688
rect 295886 234676 295892 234688
rect 295944 234676 295950 234728
rect 296714 234676 296720 234728
rect 296772 234716 296778 234728
rect 298278 234716 298284 234728
rect 296772 234688 298284 234716
rect 296772 234676 296778 234688
rect 298278 234676 298284 234688
rect 298336 234676 298342 234728
rect 298462 234676 298468 234728
rect 298520 234716 298526 234728
rect 301038 234716 301044 234728
rect 298520 234688 301044 234716
rect 298520 234676 298526 234688
rect 301038 234676 301044 234688
rect 301096 234676 301102 234728
rect 308122 234676 308128 234728
rect 308180 234716 308186 234728
rect 308858 234716 308864 234728
rect 308180 234688 308864 234716
rect 308180 234676 308186 234688
rect 308858 234676 308864 234688
rect 308916 234676 308922 234728
rect 310238 234676 310244 234728
rect 310296 234716 310302 234728
rect 311434 234716 311440 234728
rect 310296 234688 311440 234716
rect 310296 234676 310302 234688
rect 311434 234676 311440 234688
rect 311492 234676 311498 234728
rect 312722 234676 312728 234728
rect 312780 234716 312786 234728
rect 314102 234716 314108 234728
rect 312780 234688 314108 234716
rect 312780 234676 312786 234688
rect 314102 234676 314108 234688
rect 314160 234676 314166 234728
rect 314194 234676 314200 234728
rect 314252 234716 314258 234728
rect 314562 234716 314568 234728
rect 314252 234688 314568 234716
rect 314252 234676 314258 234688
rect 314562 234676 314568 234688
rect 314620 234676 314626 234728
rect 316678 234676 316684 234728
rect 316736 234716 316742 234728
rect 317230 234716 317236 234728
rect 316736 234688 317236 234716
rect 316736 234676 316742 234688
rect 317230 234676 317236 234688
rect 317288 234676 317294 234728
rect 318426 234676 318432 234728
rect 318484 234716 318490 234728
rect 319898 234716 319904 234728
rect 318484 234688 319904 234716
rect 318484 234676 318490 234688
rect 319898 234676 319904 234688
rect 319956 234676 319962 234728
rect 321278 234676 321284 234728
rect 321336 234716 321342 234728
rect 322474 234716 322480 234728
rect 321336 234688 322480 234716
rect 321336 234676 321342 234688
rect 322474 234676 322480 234688
rect 322532 234676 322538 234728
rect 323762 234676 323768 234728
rect 323820 234716 323826 234728
rect 325326 234716 325332 234728
rect 323820 234688 325332 234716
rect 323820 234676 323826 234688
rect 325326 234676 325332 234688
rect 325384 234676 325390 234728
rect 327350 234676 327356 234728
rect 327408 234716 327414 234728
rect 328362 234716 328368 234728
rect 327408 234688 328368 234716
rect 327408 234676 327414 234688
rect 328362 234676 328368 234688
rect 328420 234676 328426 234728
rect 330202 234676 330208 234728
rect 330260 234716 330266 234728
rect 331030 234716 331036 234728
rect 330260 234688 331036 234716
rect 330260 234676 330266 234688
rect 331030 234676 331036 234688
rect 331088 234676 331094 234728
rect 332042 234676 332048 234728
rect 332100 234716 332106 234728
rect 333514 234716 333520 234728
rect 332100 234688 333520 234716
rect 332100 234676 332106 234688
rect 333514 234676 333520 234688
rect 333572 234676 333578 234728
rect 334158 234676 334164 234728
rect 334216 234716 334222 234728
rect 336090 234716 336096 234728
rect 334216 234688 336096 234716
rect 334216 234676 334222 234688
rect 336090 234676 336096 234688
rect 336148 234676 336154 234728
rect 337378 234676 337384 234728
rect 337436 234716 337442 234728
rect 338850 234716 338856 234728
rect 337436 234688 338856 234716
rect 337436 234676 337442 234688
rect 338850 234676 338856 234688
rect 338908 234676 338914 234728
rect 340598 234676 340604 234728
rect 340656 234716 340662 234728
rect 341978 234716 341984 234728
rect 340656 234688 341984 234716
rect 340656 234676 340662 234688
rect 341978 234676 341984 234688
rect 342036 234676 342042 234728
rect 343450 234676 343456 234728
rect 343508 234716 343514 234728
rect 344646 234716 344652 234728
rect 343508 234688 344652 234716
rect 343508 234676 343514 234688
rect 344646 234676 344652 234688
rect 344704 234676 344710 234728
rect 346302 234676 346308 234728
rect 346360 234716 346366 234728
rect 347590 234716 347596 234728
rect 346360 234688 347596 234716
rect 346360 234676 346366 234688
rect 347590 234676 347596 234688
rect 347648 234676 347654 234728
rect 349154 234676 349160 234728
rect 349212 234716 349218 234728
rect 350258 234716 350264 234728
rect 349212 234688 350264 234716
rect 349212 234676 349218 234688
rect 350258 234676 350264 234688
rect 350316 234676 350322 234728
rect 350534 234676 350540 234728
rect 350592 234716 350598 234728
rect 352558 234716 352564 234728
rect 350592 234688 352564 234716
rect 350592 234676 350598 234688
rect 352558 234676 352564 234688
rect 352616 234676 352622 234728
rect 353754 234676 353760 234728
rect 353812 234716 353818 234728
rect 355410 234716 355416 234728
rect 353812 234688 355416 234716
rect 353812 234676 353818 234688
rect 355410 234676 355416 234688
rect 355468 234676 355474 234728
rect 356606 234676 356612 234728
rect 356664 234716 356670 234728
rect 358078 234716 358084 234728
rect 356664 234688 358084 234716
rect 356664 234676 356670 234688
rect 358078 234676 358084 234688
rect 358136 234676 358142 234728
rect 359458 234676 359464 234728
rect 359516 234716 359522 234728
rect 361390 234716 361396 234728
rect 359516 234688 361396 234716
rect 359516 234676 359522 234688
rect 361390 234676 361396 234688
rect 361448 234676 361454 234728
rect 362310 234676 362316 234728
rect 362368 234716 362374 234728
rect 364058 234716 364064 234728
rect 362368 234688 364064 234716
rect 362368 234676 362374 234688
rect 364058 234676 364064 234688
rect 364116 234676 364122 234728
rect 375466 234676 375472 234728
rect 375524 234716 375530 234728
rect 379422 234716 379428 234728
rect 375524 234688 379428 234716
rect 375524 234676 375530 234688
rect 379422 234676 379428 234688
rect 379480 234676 379486 234728
rect 384758 234676 384764 234728
rect 384816 234716 384822 234728
rect 386230 234716 386236 234728
rect 384816 234688 386236 234716
rect 384816 234676 384822 234688
rect 386230 234676 386236 234688
rect 386288 234676 386294 234728
rect 387242 234676 387248 234728
rect 387300 234716 387306 234728
rect 389082 234716 389088 234728
rect 387300 234688 389088 234716
rect 387300 234676 387306 234688
rect 389082 234676 389088 234688
rect 389140 234676 389146 234728
rect 398282 234676 398288 234728
rect 398340 234716 398346 234728
rect 403802 234716 403808 234728
rect 398340 234688 403808 234716
rect 398340 234676 398346 234688
rect 403802 234676 403808 234688
rect 403860 234676 403866 234728
rect 411530 234676 411536 234728
rect 411588 234716 411594 234728
rect 413830 234716 413836 234728
rect 411588 234688 413836 234716
rect 411588 234676 411594 234688
rect 413830 234676 413836 234688
rect 413888 234676 413894 234728
rect 262490 234648 262496 234660
rect 252940 234620 262496 234648
rect 262490 234608 262496 234620
rect 262548 234608 262554 234660
rect 267642 234608 267648 234660
rect 267700 234648 267706 234660
rect 282086 234648 282092 234660
rect 267700 234620 282092 234648
rect 267700 234608 267706 234620
rect 282086 234608 282092 234620
rect 282144 234608 282150 234660
rect 289814 234608 289820 234660
rect 289872 234648 289878 234660
rect 292390 234648 292396 234660
rect 289872 234620 292396 234648
rect 289872 234608 289878 234620
rect 292390 234608 292396 234620
rect 292448 234608 292454 234660
rect 292666 234608 292672 234660
rect 292724 234648 292730 234660
rect 293862 234648 293868 234660
rect 292724 234620 293868 234648
rect 292724 234608 292730 234620
rect 293862 234608 293868 234620
rect 293920 234608 293926 234660
rect 294966 234608 294972 234660
rect 295024 234648 295030 234660
rect 295426 234648 295432 234660
rect 295024 234620 295432 234648
rect 295024 234608 295030 234620
rect 295426 234608 295432 234620
rect 295484 234608 295490 234660
rect 295794 234608 295800 234660
rect 295852 234648 295858 234660
rect 297082 234648 297088 234660
rect 295852 234620 297088 234648
rect 295852 234608 295858 234620
rect 297082 234608 297088 234620
rect 297140 234608 297146 234660
rect 298830 234608 298836 234660
rect 298888 234648 298894 234660
rect 300946 234648 300952 234660
rect 298888 234620 300952 234648
rect 298888 234608 298894 234620
rect 300946 234608 300952 234620
rect 301004 234608 301010 234660
rect 305270 234608 305276 234660
rect 305328 234648 305334 234660
rect 306282 234648 306288 234660
rect 305328 234620 306288 234648
rect 305328 234608 305334 234620
rect 306282 234608 306288 234620
rect 306340 234608 306346 234660
rect 307754 234608 307760 234660
rect 307812 234648 307818 234660
rect 308490 234648 308496 234660
rect 307812 234620 308496 234648
rect 307812 234608 307818 234620
rect 308490 234608 308496 234620
rect 308548 234608 308554 234660
rect 310974 234608 310980 234660
rect 311032 234648 311038 234660
rect 311618 234648 311624 234660
rect 311032 234620 311624 234648
rect 311032 234608 311038 234620
rect 311618 234608 311624 234620
rect 311676 234608 311682 234660
rect 313826 234608 313832 234660
rect 313884 234648 313890 234660
rect 314378 234648 314384 234660
rect 313884 234620 314384 234648
rect 313884 234608 313890 234620
rect 314378 234608 314384 234620
rect 314436 234608 314442 234660
rect 315574 234608 315580 234660
rect 315632 234648 315638 234660
rect 316954 234648 316960 234660
rect 315632 234620 316960 234648
rect 315632 234608 315638 234620
rect 316954 234608 316960 234620
rect 317012 234608 317018 234660
rect 319530 234608 319536 234660
rect 319588 234648 319594 234660
rect 319990 234648 319996 234660
rect 319588 234620 319996 234648
rect 319588 234608 319594 234620
rect 319990 234608 319996 234620
rect 320048 234608 320054 234660
rect 322382 234608 322388 234660
rect 322440 234648 322446 234660
rect 322658 234648 322664 234660
rect 322440 234620 322664 234648
rect 322440 234608 322446 234620
rect 322658 234608 322664 234620
rect 322716 234608 322722 234660
rect 323486 234608 323492 234660
rect 323544 234648 323550 234660
rect 325142 234648 325148 234660
rect 323544 234620 325148 234648
rect 323544 234608 323550 234620
rect 325142 234608 325148 234620
rect 325200 234608 325206 234660
rect 326614 234608 326620 234660
rect 326672 234648 326678 234660
rect 327902 234648 327908 234660
rect 326672 234620 327908 234648
rect 326672 234608 326678 234620
rect 327902 234608 327908 234620
rect 327960 234608 327966 234660
rect 329834 234608 329840 234660
rect 329892 234648 329898 234660
rect 330754 234648 330760 234660
rect 329892 234620 330760 234648
rect 329892 234608 329898 234620
rect 330754 234608 330760 234620
rect 330812 234608 330818 234660
rect 332318 234608 332324 234660
rect 332376 234648 332382 234660
rect 333606 234648 333612 234660
rect 332376 234620 333612 234648
rect 332376 234608 332382 234620
rect 333606 234608 333612 234620
rect 333664 234608 333670 234660
rect 335538 234608 335544 234660
rect 335596 234648 335602 234660
rect 336458 234648 336464 234660
rect 335596 234620 336464 234648
rect 335596 234608 335602 234620
rect 336458 234608 336464 234620
rect 336516 234608 336522 234660
rect 338022 234608 338028 234660
rect 338080 234648 338086 234660
rect 338942 234648 338948 234660
rect 338080 234620 338948 234648
rect 338080 234608 338086 234620
rect 338942 234608 338948 234620
rect 339000 234608 339006 234660
rect 340230 234608 340236 234660
rect 340288 234648 340294 234660
rect 341610 234648 341616 234660
rect 340288 234620 341616 234648
rect 340288 234608 340294 234620
rect 341610 234608 341616 234620
rect 341668 234608 341674 234660
rect 343726 234608 343732 234660
rect 343784 234648 343790 234660
rect 344830 234648 344836 234660
rect 343784 234620 344836 234648
rect 343784 234608 343790 234620
rect 344830 234608 344836 234620
rect 344888 234608 344894 234660
rect 346578 234608 346584 234660
rect 346636 234648 346642 234660
rect 347498 234648 347504 234660
rect 346636 234620 347504 234648
rect 346636 234608 346642 234620
rect 347498 234608 347504 234620
rect 347556 234608 347562 234660
rect 349430 234608 349436 234660
rect 349488 234648 349494 234660
rect 350350 234648 350356 234660
rect 349488 234620 350356 234648
rect 349488 234608 349494 234620
rect 350350 234608 350356 234620
rect 350408 234608 350414 234660
rect 352006 234608 352012 234660
rect 352064 234648 352070 234660
rect 352650 234648 352656 234660
rect 352064 234620 352656 234648
rect 352064 234608 352070 234620
rect 352650 234608 352656 234620
rect 352708 234608 352714 234660
rect 354858 234608 354864 234660
rect 354916 234648 354922 234660
rect 355686 234648 355692 234660
rect 354916 234620 355692 234648
rect 354916 234608 354922 234620
rect 355686 234608 355692 234620
rect 355744 234608 355750 234660
rect 357710 234608 357716 234660
rect 357768 234648 357774 234660
rect 358446 234648 358452 234660
rect 357768 234620 358452 234648
rect 357768 234608 357774 234620
rect 358446 234608 358452 234620
rect 358504 234608 358510 234660
rect 360562 234608 360568 234660
rect 360620 234648 360626 234660
rect 361298 234648 361304 234660
rect 360620 234620 361304 234648
rect 360620 234608 360626 234620
rect 361298 234608 361304 234620
rect 361356 234608 361362 234660
rect 361942 234608 361948 234660
rect 362000 234648 362006 234660
rect 363506 234648 363512 234660
rect 362000 234620 363512 234648
rect 362000 234608 362006 234620
rect 363506 234608 363512 234620
rect 363564 234608 363570 234660
rect 364794 234608 364800 234660
rect 364852 234648 364858 234660
rect 367002 234648 367008 234660
rect 364852 234620 367008 234648
rect 364852 234608 364858 234620
rect 367002 234608 367008 234620
rect 367060 234608 367066 234660
rect 367646 234608 367652 234660
rect 367704 234648 367710 234660
rect 369118 234648 369124 234660
rect 367704 234620 369124 234648
rect 367704 234608 367710 234620
rect 369118 234608 369124 234620
rect 369176 234608 369182 234660
rect 370498 234608 370504 234660
rect 370556 234648 370562 234660
rect 371970 234648 371976 234660
rect 370556 234620 371976 234648
rect 370556 234608 370562 234620
rect 371970 234608 371976 234620
rect 372028 234608 372034 234660
rect 373350 234608 373356 234660
rect 373408 234648 373414 234660
rect 374730 234648 374736 234660
rect 373408 234620 374736 234648
rect 373408 234608 373414 234620
rect 374730 234608 374736 234620
rect 374788 234608 374794 234660
rect 376938 234608 376944 234660
rect 376996 234648 377002 234660
rect 377950 234648 377956 234660
rect 376996 234620 377956 234648
rect 376996 234608 377002 234620
rect 377950 234608 377956 234620
rect 378008 234608 378014 234660
rect 379790 234608 379796 234660
rect 379848 234648 379854 234660
rect 380618 234648 380624 234660
rect 379848 234620 380624 234648
rect 379848 234608 379854 234620
rect 380618 234608 380624 234620
rect 380676 234608 380682 234660
rect 382274 234608 382280 234660
rect 382332 234648 382338 234660
rect 384942 234648 384948 234660
rect 382332 234620 384948 234648
rect 382332 234608 382338 234620
rect 384942 234608 384948 234620
rect 385000 234608 385006 234660
rect 385126 234608 385132 234660
rect 385184 234648 385190 234660
rect 386322 234648 386328 234660
rect 385184 234620 386328 234648
rect 385184 234608 385190 234620
rect 386322 234608 386328 234620
rect 386380 234608 386386 234660
rect 386874 234608 386880 234660
rect 386932 234648 386938 234660
rect 388990 234648 388996 234660
rect 386932 234620 388996 234648
rect 386932 234608 386938 234620
rect 388990 234608 388996 234620
rect 389048 234608 389054 234660
rect 390094 234608 390100 234660
rect 390152 234648 390158 234660
rect 391842 234648 391848 234660
rect 390152 234620 391848 234648
rect 390152 234608 390158 234620
rect 391842 234608 391848 234620
rect 391900 234608 391906 234660
rect 391934 234608 391940 234660
rect 391992 234648 391998 234660
rect 403066 234648 403072 234660
rect 391992 234620 403072 234648
rect 391992 234608 391998 234620
rect 403066 234608 403072 234620
rect 403124 234608 403130 234660
rect 403618 234608 403624 234660
rect 403676 234648 403682 234660
rect 407390 234648 407396 234660
rect 403676 234620 407396 234648
rect 403676 234608 403682 234620
rect 407390 234608 407396 234620
rect 407448 234608 407454 234660
rect 411898 234608 411904 234660
rect 411956 234648 411962 234660
rect 413922 234648 413928 234660
rect 411956 234620 413928 234648
rect 411956 234608 411962 234620
rect 413922 234608 413928 234620
rect 413980 234608 413986 234660
rect 42150 234200 42156 234252
rect 42208 234240 42214 234252
rect 43070 234240 43076 234252
rect 42208 234212 43076 234240
rect 42208 234200 42214 234212
rect 43070 234200 43076 234212
rect 43128 234200 43134 234252
rect 389726 233724 389732 233776
rect 389784 233764 389790 233776
rect 401318 233764 401324 233776
rect 389784 233736 401324 233764
rect 389784 233724 389790 233736
rect 401318 233724 401324 233736
rect 401376 233724 401382 233776
rect 377674 233452 377680 233504
rect 377732 233492 377738 233504
rect 489914 233492 489920 233504
rect 377732 233464 489920 233492
rect 377732 233452 377738 233464
rect 489914 233452 489920 233464
rect 489972 233452 489978 233504
rect 393682 233384 393688 233436
rect 393740 233424 393746 233436
rect 528554 233424 528560 233436
rect 393740 233396 528560 233424
rect 393740 233384 393746 233396
rect 528554 233384 528560 233396
rect 528612 233384 528618 233436
rect 42150 233316 42156 233368
rect 42208 233356 42214 233368
rect 43898 233356 43904 233368
rect 42208 233328 43904 233356
rect 42208 233316 42214 233328
rect 43898 233316 43904 233328
rect 43956 233316 43962 233368
rect 396902 233316 396908 233368
rect 396960 233356 396966 233368
rect 536834 233356 536840 233368
rect 396960 233328 536840 233356
rect 396960 233316 396966 233328
rect 536834 233316 536840 233328
rect 536892 233316 536898 233368
rect 397914 233248 397920 233300
rect 397972 233288 397978 233300
rect 539594 233288 539600 233300
rect 397972 233260 539600 233288
rect 397972 233248 397978 233260
rect 539594 233248 539600 233260
rect 539652 233248 539658 233300
rect 287238 233180 287244 233232
rect 287296 233220 287302 233232
rect 287882 233220 287888 233232
rect 287296 233192 287888 233220
rect 287296 233180 287302 233192
rect 287882 233180 287888 233192
rect 287940 233180 287946 233232
rect 400122 233180 400128 233232
rect 400180 233220 400186 233232
rect 542446 233220 542452 233232
rect 400180 233192 542452 233220
rect 400180 233180 400186 233192
rect 542446 233180 542452 233192
rect 542504 233180 542510 233232
rect 284386 233112 284392 233164
rect 284444 233152 284450 233164
rect 285030 233152 285036 233164
rect 284444 233124 285036 233152
rect 284444 233112 284450 233124
rect 285030 233112 285036 233124
rect 285088 233112 285094 233164
rect 287054 233112 287060 233164
rect 287112 233152 287118 233164
rect 287606 233152 287612 233164
rect 287112 233124 287612 233152
rect 287112 233112 287118 233124
rect 287606 233112 287612 233124
rect 287664 233112 287670 233164
rect 193674 233044 193680 233096
rect 193732 233084 193738 233096
rect 195514 233084 195520 233096
rect 193732 233056 195520 233084
rect 193732 233044 193738 233056
rect 195514 233044 195520 233056
rect 195572 233044 195578 233096
rect 196158 233044 196164 233096
rect 196216 233084 196222 233096
rect 198366 233084 198372 233096
rect 196216 233056 198372 233084
rect 196216 233044 196222 233056
rect 198366 233044 198372 233056
rect 198424 233044 198430 233096
rect 226610 233044 226616 233096
rect 226668 233084 226674 233096
rect 227622 233084 227628 233096
rect 226668 233056 227628 233084
rect 226668 233044 226674 233056
rect 227622 233044 227628 233056
rect 227680 233044 227686 233096
rect 229278 233044 229284 233096
rect 229336 233084 229342 233096
rect 230474 233084 230480 233096
rect 229336 233056 230480 233084
rect 229336 233044 229342 233056
rect 230474 233044 230480 233056
rect 230532 233044 230538 233096
rect 232038 233044 232044 233096
rect 232096 233084 232102 233096
rect 233326 233084 233332 233096
rect 232096 233056 233332 233084
rect 232096 233044 232102 233056
rect 233326 233044 233332 233056
rect 233384 233044 233390 233096
rect 234798 233044 234804 233096
rect 234856 233084 234862 233096
rect 236178 233084 236184 233096
rect 234856 233056 236184 233084
rect 234856 233044 234862 233056
rect 236178 233044 236184 233056
rect 236236 233044 236242 233096
rect 240318 233044 240324 233096
rect 240376 233084 240382 233096
rect 241882 233084 241888 233096
rect 240376 233056 241888 233084
rect 240376 233044 240382 233056
rect 241882 233044 241888 233056
rect 241940 233044 241946 233096
rect 243078 233044 243084 233096
rect 243136 233084 243142 233096
rect 244734 233084 244740 233096
rect 243136 233056 244740 233084
rect 243136 233044 243142 233056
rect 244734 233044 244740 233056
rect 244792 233044 244798 233096
rect 245838 233044 245844 233096
rect 245896 233084 245902 233096
rect 247586 233084 247592 233096
rect 245896 233056 247592 233084
rect 245896 233044 245902 233056
rect 247586 233044 247592 233056
rect 247644 233044 247650 233096
rect 251358 233044 251364 233096
rect 251416 233084 251422 233096
rect 253290 233084 253296 233096
rect 251416 233056 253296 233084
rect 251416 233044 251422 233056
rect 253290 233044 253296 233056
rect 253348 233044 253354 233096
rect 281718 233044 281724 233096
rect 281776 233084 281782 233096
rect 283282 233084 283288 233096
rect 281776 233056 283288 233084
rect 281776 233044 281782 233056
rect 283282 233044 283288 233056
rect 283340 233044 283346 233096
rect 290274 233044 290280 233096
rect 290332 233084 290338 233096
rect 291102 233084 291108 233096
rect 290332 233056 291108 233084
rect 290332 233044 290338 233056
rect 291102 233044 291108 233056
rect 291160 233044 291166 233096
rect 190638 232976 190644 233028
rect 190696 233016 190702 233028
rect 192386 233016 192392 233028
rect 190696 232988 192392 233016
rect 190696 232976 190702 232988
rect 192386 232976 192392 232988
rect 192444 232976 192450 233028
rect 193490 232976 193496 233028
rect 193548 233016 193554 233028
rect 194870 233016 194876 233028
rect 193548 232988 194876 233016
rect 193548 232976 193554 232988
rect 194870 232976 194876 232988
rect 194928 232976 194934 233028
rect 196342 232976 196348 233028
rect 196400 233016 196406 233028
rect 198090 233016 198096 233028
rect 196400 232988 198096 233016
rect 196400 232976 196406 232988
rect 198090 232976 198096 232988
rect 198148 232976 198154 233028
rect 218422 232976 218428 233028
rect 218480 233016 218486 233028
rect 220170 233016 220176 233028
rect 218480 232988 220176 233016
rect 218480 232976 218486 232988
rect 220170 232976 220176 232988
rect 220228 232976 220234 233028
rect 221090 232976 221096 233028
rect 221148 233016 221154 233028
rect 221918 233016 221924 233028
rect 221148 232988 221924 233016
rect 221148 232976 221154 232988
rect 221918 232976 221924 232988
rect 221976 232976 221982 233028
rect 223758 232976 223764 233028
rect 223816 233016 223822 233028
rect 224770 233016 224776 233028
rect 223816 232988 224776 233016
rect 223816 232976 223822 232988
rect 224770 232976 224776 232988
rect 224828 232976 224834 233028
rect 226794 232976 226800 233028
rect 226852 233016 226858 233028
rect 227254 233016 227260 233028
rect 226852 232988 227260 233016
rect 226852 232976 226858 232988
rect 227254 232976 227260 232988
rect 227312 232976 227318 233028
rect 229186 232976 229192 233028
rect 229244 233016 229250 233028
rect 230106 233016 230112 233028
rect 229244 232988 230112 233016
rect 229244 232976 229250 232988
rect 230106 232976 230112 232988
rect 230164 232976 230170 233028
rect 232314 232976 232320 233028
rect 232372 233016 232378 233028
rect 232958 233016 232964 233028
rect 232372 232988 232964 233016
rect 232372 232976 232378 232988
rect 232958 232976 232964 232988
rect 233016 232976 233022 233028
rect 235166 232976 235172 233028
rect 235224 233016 235230 233028
rect 235810 233016 235816 233028
rect 235224 232988 235816 233016
rect 235224 232976 235230 232988
rect 235810 232976 235816 232988
rect 235868 232976 235874 233028
rect 237742 232976 237748 233028
rect 237800 233016 237806 233028
rect 238662 233016 238668 233028
rect 237800 232988 238668 233016
rect 237800 232976 237806 232988
rect 238662 232976 238668 232988
rect 238720 232976 238726 233028
rect 240502 232976 240508 233028
rect 240560 233016 240566 233028
rect 241514 233016 241520 233028
rect 240560 232988 241520 233016
rect 240560 232976 240566 232988
rect 241514 232976 241520 232988
rect 241572 232976 241578 233028
rect 243262 232976 243268 233028
rect 243320 233016 243326 233028
rect 244366 233016 244372 233028
rect 243320 232988 244372 233016
rect 243320 232976 243326 232988
rect 244366 232976 244372 232988
rect 244424 232976 244430 233028
rect 246022 232976 246028 233028
rect 246080 233016 246086 233028
rect 247218 233016 247224 233028
rect 246080 232988 247224 233016
rect 246080 232976 246086 232988
rect 247218 232976 247224 232988
rect 247276 232976 247282 233028
rect 248598 232976 248604 233028
rect 248656 233016 248662 233028
rect 250438 233016 250444 233028
rect 248656 232988 250444 233016
rect 248656 232976 248662 232988
rect 250438 232976 250444 232988
rect 250496 232976 250502 233028
rect 251450 232976 251456 233028
rect 251508 233016 251514 233028
rect 252922 233016 252928 233028
rect 251508 232988 252928 233016
rect 251508 232976 251514 232988
rect 252922 232976 252928 232988
rect 252980 232976 252986 233028
rect 254210 232976 254216 233028
rect 254268 233016 254274 233028
rect 255774 233016 255780 233028
rect 254268 232988 255780 233016
rect 254268 232976 254274 232988
rect 255774 232976 255780 232988
rect 255832 232976 255838 233028
rect 257062 232976 257068 233028
rect 257120 233016 257126 233028
rect 258626 233016 258632 233028
rect 257120 232988 258632 233016
rect 257120 232976 257126 232988
rect 258626 232976 258632 232988
rect 258684 232976 258690 233028
rect 259822 232976 259828 233028
rect 259880 233016 259886 233028
rect 261478 233016 261484 233028
rect 259880 232988 261484 233016
rect 259880 232976 259886 232988
rect 261478 232976 261484 232988
rect 261536 232976 261542 233028
rect 262582 232976 262588 233028
rect 262640 233016 262646 233028
rect 264330 233016 264336 233028
rect 262640 232988 264336 233016
rect 262640 232976 262646 232988
rect 264330 232976 264336 232988
rect 264388 232976 264394 233028
rect 268194 232976 268200 233028
rect 268252 233016 268258 233028
rect 270034 233016 270040 233028
rect 268252 232988 270040 233016
rect 268252 232976 268258 232988
rect 270034 232976 270040 232988
rect 270092 232976 270098 233028
rect 281994 232976 282000 233028
rect 282052 233016 282058 233028
rect 283650 233016 283656 233028
rect 282052 232988 283656 233016
rect 282052 232976 282058 232988
rect 283650 232976 283656 232988
rect 283708 232976 283714 233028
rect 284478 232976 284484 233028
rect 284536 233016 284542 233028
rect 286502 233016 286508 233028
rect 284536 232988 286508 233016
rect 284536 232976 284542 232988
rect 286502 232976 286508 232988
rect 286560 232976 286566 233028
rect 287882 232976 287888 233028
rect 287940 233016 287946 233028
rect 289354 233016 289360 233028
rect 287940 232988 289360 233016
rect 287940 232976 287946 232988
rect 289354 232976 289360 232988
rect 289412 232976 289418 233028
rect 290366 232976 290372 233028
rect 290424 233016 290430 233028
rect 291470 233016 291476 233028
rect 290424 232988 291476 233016
rect 290424 232976 290430 232988
rect 291470 232976 291476 232988
rect 291528 232976 291534 233028
rect 292758 232976 292764 233028
rect 292816 233016 292822 233028
rect 293954 233016 293960 233028
rect 292816 232988 293960 233016
rect 292816 232976 292822 232988
rect 293954 232976 293960 232988
rect 294012 232976 294018 233028
rect 196434 232908 196440 232960
rect 196492 232948 196498 232960
rect 197722 232948 197728 232960
rect 196492 232920 197728 232948
rect 196492 232908 196498 232920
rect 197722 232908 197728 232920
rect 197780 232908 197786 232960
rect 237650 232908 237656 232960
rect 237708 232948 237714 232960
rect 239030 232948 239036 232960
rect 237708 232920 239036 232948
rect 237708 232908 237714 232920
rect 239030 232908 239036 232920
rect 239088 232908 239094 232960
rect 281810 232908 281816 232960
rect 281868 232948 281874 232960
rect 283926 232948 283932 232960
rect 281868 232920 283932 232948
rect 281868 232908 281874 232920
rect 283926 232908 283932 232920
rect 283984 232908 283990 232960
rect 287422 232908 287428 232960
rect 287480 232948 287486 232960
rect 288618 232948 288624 232960
rect 287480 232920 288624 232948
rect 287480 232908 287486 232920
rect 288618 232908 288624 232920
rect 288676 232908 288682 232960
rect 290182 232908 290188 232960
rect 290240 232948 290246 232960
rect 291838 232948 291844 232960
rect 290240 232920 291844 232948
rect 290240 232908 290246 232920
rect 291838 232908 291844 232920
rect 291896 232908 291902 232960
rect 314010 232908 314016 232960
rect 314068 232948 314074 232960
rect 314470 232948 314476 232960
rect 314068 232920 314476 232948
rect 314068 232908 314074 232920
rect 314470 232908 314476 232920
rect 314528 232908 314534 232960
rect 335446 232908 335452 232960
rect 335504 232948 335510 232960
rect 336366 232948 336372 232960
rect 335504 232920 336372 232948
rect 335504 232908 335510 232920
rect 336366 232908 336372 232920
rect 336424 232908 336430 232960
rect 196250 232840 196256 232892
rect 196308 232880 196314 232892
rect 196618 232880 196624 232892
rect 196308 232852 196624 232880
rect 196308 232840 196314 232852
rect 196618 232840 196624 232852
rect 196676 232840 196682 232892
rect 287146 232840 287152 232892
rect 287204 232880 287210 232892
rect 288250 232880 288256 232892
rect 287204 232852 288256 232880
rect 287204 232840 287210 232852
rect 288250 232840 288256 232852
rect 288308 232840 288314 232892
rect 284846 232636 284852 232688
rect 284904 232676 284910 232688
rect 286134 232676 286140 232688
rect 284904 232648 286140 232676
rect 284904 232636 284910 232648
rect 286134 232636 286140 232648
rect 286192 232636 286198 232688
rect 341702 231752 341708 231804
rect 341760 231792 341766 231804
rect 403618 231792 403624 231804
rect 341760 231764 403624 231792
rect 341760 231752 341766 231764
rect 403618 231752 403624 231764
rect 403676 231752 403682 231804
rect 363046 231684 363052 231736
rect 363104 231724 363110 231736
rect 454126 231724 454132 231736
rect 363104 231696 454132 231724
rect 363104 231684 363110 231696
rect 454126 231684 454132 231696
rect 454184 231684 454190 231736
rect 364426 231616 364432 231668
rect 364484 231656 364490 231668
rect 457438 231656 457444 231668
rect 364484 231628 457444 231656
rect 364484 231616 364490 231628
rect 457438 231616 457444 231628
rect 457496 231616 457502 231668
rect 367278 231548 367284 231600
rect 367336 231588 367342 231600
rect 464246 231588 464252 231600
rect 367336 231560 464252 231588
rect 367336 231548 367342 231560
rect 464246 231548 464252 231560
rect 464304 231548 464310 231600
rect 287790 231480 287796 231532
rect 287848 231520 287854 231532
rect 288986 231520 288992 231532
rect 287848 231492 288992 231520
rect 287848 231480 287854 231492
rect 288986 231480 288992 231492
rect 289044 231480 289050 231532
rect 365898 231480 365904 231532
rect 365956 231520 365962 231532
rect 460934 231520 460940 231532
rect 365956 231492 460940 231520
rect 365956 231480 365962 231492
rect 460934 231480 460940 231492
rect 460992 231480 460998 231532
rect 370130 231412 370136 231464
rect 370188 231452 370194 231464
rect 470962 231452 470968 231464
rect 370188 231424 470968 231452
rect 370188 231412 370194 231424
rect 470962 231412 470968 231424
rect 471020 231412 471026 231464
rect 368750 231344 368756 231396
rect 368808 231384 368814 231396
rect 467558 231384 467564 231396
rect 368808 231356 467564 231384
rect 368808 231344 368814 231356
rect 467558 231344 467564 231356
rect 467616 231344 467622 231396
rect 371602 231276 371608 231328
rect 371660 231316 371666 231328
rect 474274 231316 474280 231328
rect 371660 231288 474280 231316
rect 371660 231276 371666 231288
rect 474274 231276 474280 231288
rect 474332 231276 474338 231328
rect 372982 231208 372988 231260
rect 373040 231248 373046 231260
rect 477678 231248 477684 231260
rect 373040 231220 477684 231248
rect 373040 231208 373046 231220
rect 477678 231208 477684 231220
rect 477736 231208 477742 231260
rect 374454 231140 374460 231192
rect 374512 231180 374518 231192
rect 480990 231180 480996 231192
rect 374512 231152 480996 231180
rect 374512 231140 374518 231152
rect 480990 231140 480996 231152
rect 481048 231140 481054 231192
rect 42150 231072 42156 231124
rect 42208 231112 42214 231124
rect 43622 231112 43628 231124
rect 42208 231084 43628 231112
rect 42208 231072 42214 231084
rect 43622 231072 43628 231084
rect 43680 231072 43686 231124
rect 374546 231072 374552 231124
rect 374604 231112 374610 231124
rect 483014 231112 483020 231124
rect 374604 231084 483020 231112
rect 374604 231072 374610 231084
rect 483014 231072 483020 231084
rect 483072 231072 483078 231124
rect 186406 231004 186412 231056
rect 186464 231044 186470 231056
rect 248230 231044 248236 231056
rect 186464 231016 248236 231044
rect 186464 231004 186470 231016
rect 248230 231004 248236 231016
rect 248288 231004 248294 231056
rect 376202 231004 376208 231056
rect 376260 231044 376266 231056
rect 487154 231044 487160 231056
rect 376260 231016 487160 231044
rect 376260 231004 376266 231016
rect 487154 231004 487160 231016
rect 487212 231004 487218 231056
rect 179690 230936 179696 230988
rect 179748 230976 179754 230988
rect 245378 230976 245384 230988
rect 179748 230948 245384 230976
rect 179748 230936 179754 230948
rect 245378 230936 245384 230948
rect 245436 230936 245442 230988
rect 389358 230936 389364 230988
rect 389416 230976 389422 230988
rect 389416 230948 401548 230976
rect 389416 230936 389422 230948
rect 183094 230868 183100 230920
rect 183152 230908 183158 230920
rect 246758 230908 246764 230920
rect 183152 230880 246764 230908
rect 183152 230868 183158 230880
rect 246758 230868 246764 230880
rect 246816 230868 246822 230920
rect 390462 230868 390468 230920
rect 390520 230908 390526 230920
rect 401520 230908 401548 230948
rect 401594 230936 401600 230988
rect 401652 230976 401658 230988
rect 515490 230976 515496 230988
rect 401652 230948 515496 230976
rect 401652 230936 401658 230948
rect 515490 230936 515496 230948
rect 515548 230936 515554 230988
rect 518066 230908 518072 230920
rect 390520 230880 401456 230908
rect 401520 230880 518072 230908
rect 390520 230868 390526 230880
rect 172974 230800 172980 230852
rect 173032 230840 173038 230852
rect 242526 230840 242532 230852
rect 173032 230812 242532 230840
rect 173032 230800 173038 230812
rect 242526 230800 242532 230812
rect 242584 230800 242590 230852
rect 391566 230800 391572 230852
rect 391624 230840 391630 230852
rect 401428 230840 401456 230880
rect 518066 230868 518072 230880
rect 518124 230868 518130 230920
rect 518986 230840 518992 230852
rect 391624 230812 391934 230840
rect 401428 230812 518992 230840
rect 391624 230800 391630 230812
rect 176378 230732 176384 230784
rect 176436 230772 176442 230784
rect 243906 230772 243912 230784
rect 176436 230744 243912 230772
rect 176436 230732 176442 230744
rect 243906 230732 243912 230744
rect 243964 230732 243970 230784
rect 391906 230772 391934 230812
rect 518986 230800 518992 230812
rect 519044 230800 519050 230852
rect 523402 230772 523408 230784
rect 391906 230744 523408 230772
rect 523402 230732 523408 230744
rect 523460 230732 523466 230784
rect 166258 230664 166264 230716
rect 166316 230704 166322 230716
rect 239674 230704 239680 230716
rect 166316 230676 239680 230704
rect 166316 230664 166322 230676
rect 239674 230664 239680 230676
rect 239732 230664 239738 230716
rect 334894 230664 334900 230716
rect 334952 230704 334958 230716
rect 389358 230704 389364 230716
rect 334952 230676 389364 230704
rect 334952 230664 334958 230676
rect 389358 230664 389364 230676
rect 389416 230664 389422 230716
rect 392578 230664 392584 230716
rect 392636 230704 392642 230716
rect 525886 230704 525892 230716
rect 392636 230676 525892 230704
rect 392636 230664 392642 230676
rect 525886 230664 525892 230676
rect 525944 230664 525950 230716
rect 169570 230596 169576 230648
rect 169628 230636 169634 230648
rect 241054 230636 241060 230648
rect 169628 230608 241060 230636
rect 169628 230596 169634 230608
rect 241054 230596 241060 230608
rect 241112 230596 241118 230648
rect 336642 230596 336648 230648
rect 336700 230636 336706 230648
rect 392670 230636 392676 230648
rect 336700 230608 392676 230636
rect 336700 230596 336706 230608
rect 392670 230596 392676 230608
rect 392728 230596 392734 230648
rect 394786 230596 394792 230648
rect 394844 230636 394850 230648
rect 530946 230636 530952 230648
rect 394844 230608 530952 230636
rect 394844 230596 394850 230608
rect 530946 230596 530952 230608
rect 531004 230596 531010 230648
rect 42150 230528 42156 230580
rect 42208 230568 42214 230580
rect 42978 230568 42984 230580
rect 42208 230540 42984 230568
rect 42208 230528 42214 230540
rect 42978 230528 42984 230540
rect 43036 230528 43042 230580
rect 162762 230528 162768 230580
rect 162820 230568 162826 230580
rect 238202 230568 238208 230580
rect 162820 230540 238208 230568
rect 162820 230528 162826 230540
rect 238202 230528 238208 230540
rect 238260 230528 238266 230580
rect 337746 230528 337752 230580
rect 337804 230568 337810 230580
rect 395706 230568 395712 230580
rect 337804 230540 395712 230568
rect 337804 230528 337810 230540
rect 395706 230528 395712 230540
rect 395764 230528 395770 230580
rect 395798 230528 395804 230580
rect 395856 230568 395862 230580
rect 533154 230568 533160 230580
rect 395856 230540 533160 230568
rect 395856 230528 395862 230540
rect 533154 230528 533160 230540
rect 533212 230528 533218 230580
rect 46842 230460 46848 230512
rect 46900 230500 46906 230512
rect 662874 230500 662880 230512
rect 46900 230472 662880 230500
rect 46900 230460 46906 230472
rect 662874 230460 662880 230472
rect 662932 230460 662938 230512
rect 46382 230392 46388 230444
rect 46440 230432 46446 230444
rect 662782 230432 662788 230444
rect 46440 230404 662788 230432
rect 46440 230392 46446 230404
rect 662782 230392 662788 230404
rect 662840 230392 662846 230444
rect 339402 230324 339408 230376
rect 339460 230364 339466 230376
rect 399478 230364 399484 230376
rect 339460 230336 399484 230364
rect 339460 230324 339466 230336
rect 399478 230324 399484 230336
rect 399536 230324 399542 230376
rect 388346 230256 388352 230308
rect 388404 230296 388410 230308
rect 401594 230296 401600 230308
rect 388404 230268 401600 230296
rect 388404 230256 388410 230268
rect 401594 230256 401600 230268
rect 401652 230256 401658 230308
rect 42150 229848 42156 229900
rect 42208 229888 42214 229900
rect 43162 229888 43168 229900
rect 42208 229860 43168 229888
rect 42208 229848 42214 229860
rect 43162 229848 43168 229860
rect 43220 229848 43226 229900
rect 42150 229032 42156 229084
rect 42208 229072 42214 229084
rect 43530 229072 43536 229084
rect 42208 229044 43536 229072
rect 42208 229032 42214 229044
rect 43530 229032 43536 229044
rect 43588 229032 43594 229084
rect 353110 229032 353116 229084
rect 353168 229072 353174 229084
rect 428918 229072 428924 229084
rect 353168 229044 428924 229072
rect 353168 229032 353174 229044
rect 428918 229032 428924 229044
rect 428976 229032 428982 229084
rect 159542 228964 159548 229016
rect 159600 229004 159606 229016
rect 236822 229004 236828 229016
rect 159600 228976 236828 229004
rect 159600 228964 159606 228976
rect 236822 228964 236828 228976
rect 236880 228964 236886 229016
rect 354122 228964 354128 229016
rect 354180 229004 354186 229016
rect 432230 229004 432236 229016
rect 354180 228976 432236 229004
rect 354180 228964 354186 228976
rect 432230 228964 432236 228976
rect 432288 228964 432294 229016
rect 156138 228896 156144 228948
rect 156196 228936 156202 228948
rect 235350 228936 235356 228948
rect 156196 228908 235356 228936
rect 156196 228896 156202 228908
rect 235350 228896 235356 228908
rect 235408 228896 235414 228948
rect 355502 228896 355508 228948
rect 355560 228936 355566 228948
rect 435634 228936 435640 228948
rect 355560 228908 435640 228936
rect 355560 228896 355566 228908
rect 435634 228896 435640 228908
rect 435692 228896 435698 228948
rect 152826 228828 152832 228880
rect 152884 228868 152890 228880
rect 233970 228868 233976 228880
rect 152884 228840 233976 228868
rect 152884 228828 152890 228840
rect 233970 228828 233976 228840
rect 234028 228828 234034 228880
rect 354490 228828 354496 228880
rect 354548 228868 354554 228880
rect 433886 228868 433892 228880
rect 354548 228840 433892 228868
rect 354548 228828 354554 228840
rect 433886 228828 433892 228840
rect 433944 228828 433950 228880
rect 149422 228760 149428 228812
rect 149480 228800 149486 228812
rect 232498 228800 232504 228812
rect 149480 228772 232504 228800
rect 149480 228760 149486 228772
rect 232498 228760 232504 228772
rect 232556 228760 232562 228812
rect 353202 228760 353208 228812
rect 353260 228800 353266 228812
rect 430574 228800 430580 228812
rect 353260 228772 430580 228800
rect 353260 228760 353266 228772
rect 430574 228760 430580 228772
rect 430632 228760 430638 228812
rect 146018 228692 146024 228744
rect 146076 228732 146082 228744
rect 231118 228732 231124 228744
rect 146076 228704 231124 228732
rect 146076 228692 146082 228704
rect 231118 228692 231124 228704
rect 231176 228692 231182 228744
rect 357342 228692 357348 228744
rect 357400 228732 357406 228744
rect 440694 228732 440700 228744
rect 357400 228704 440700 228732
rect 357400 228692 357406 228704
rect 440694 228692 440700 228704
rect 440752 228692 440758 228744
rect 142706 228624 142712 228676
rect 142764 228664 142770 228676
rect 229646 228664 229652 228676
rect 142764 228636 229652 228664
rect 142764 228624 142770 228636
rect 229646 228624 229652 228636
rect 229704 228624 229710 228676
rect 355870 228624 355876 228676
rect 355928 228664 355934 228676
rect 437290 228664 437296 228676
rect 355928 228636 437296 228664
rect 355928 228624 355934 228636
rect 437290 228624 437296 228636
rect 437348 228624 437354 228676
rect 139210 228556 139216 228608
rect 139268 228596 139274 228608
rect 228266 228596 228272 228608
rect 139268 228568 228272 228596
rect 139268 228556 139274 228568
rect 228266 228556 228272 228568
rect 228324 228556 228330 228608
rect 356974 228556 356980 228608
rect 357032 228596 357038 228608
rect 438946 228596 438952 228608
rect 357032 228568 438952 228596
rect 357032 228556 357038 228568
rect 438946 228556 438952 228568
rect 439004 228556 439010 228608
rect 135990 228488 135996 228540
rect 136048 228528 136054 228540
rect 226702 228528 226708 228540
rect 136048 228500 226708 228528
rect 136048 228488 136054 228500
rect 226702 228488 226708 228500
rect 226760 228488 226766 228540
rect 358354 228488 358360 228540
rect 358412 228528 358418 228540
rect 442350 228528 442356 228540
rect 358412 228500 442356 228528
rect 358412 228488 358418 228500
rect 442350 228488 442356 228500
rect 442408 228488 442414 228540
rect 132402 228420 132408 228472
rect 132460 228460 132466 228472
rect 225414 228460 225420 228472
rect 132460 228432 225420 228460
rect 132460 228420 132466 228432
rect 225414 228420 225420 228432
rect 225472 228420 225478 228472
rect 359826 228420 359832 228472
rect 359884 228460 359890 228472
rect 445662 228460 445668 228472
rect 359884 228432 445668 228460
rect 359884 228420 359890 228432
rect 445662 228420 445668 228432
rect 445720 228420 445726 228472
rect 129274 228352 129280 228404
rect 129332 228392 129338 228404
rect 223942 228392 223948 228404
rect 129332 228364 223948 228392
rect 129332 228352 129338 228364
rect 223942 228352 223948 228364
rect 224000 228352 224006 228404
rect 358722 228352 358728 228404
rect 358780 228392 358786 228404
rect 444374 228392 444380 228404
rect 358780 228364 444380 228392
rect 358780 228352 358786 228364
rect 444374 228352 444380 228364
rect 444432 228352 444438 228404
rect 125870 228284 125876 228336
rect 125928 228324 125934 228336
rect 222562 228324 222568 228336
rect 125928 228296 222568 228324
rect 125928 228284 125934 228296
rect 222562 228284 222568 228296
rect 222620 228284 222626 228336
rect 360194 228284 360200 228336
rect 360252 228324 360258 228336
rect 447410 228324 447416 228336
rect 360252 228296 447416 228324
rect 360252 228284 360258 228296
rect 447410 228284 447416 228296
rect 447468 228284 447474 228336
rect 122466 228216 122472 228268
rect 122524 228256 122530 228268
rect 221182 228256 221188 228268
rect 122524 228228 221188 228256
rect 122524 228216 122530 228228
rect 221182 228216 221188 228228
rect 221240 228216 221246 228268
rect 361482 228216 361488 228268
rect 361540 228256 361546 228268
rect 449066 228256 449072 228268
rect 361540 228228 449072 228256
rect 361540 228216 361546 228228
rect 449066 228216 449072 228228
rect 449124 228216 449130 228268
rect 119154 228148 119160 228200
rect 119212 228188 119218 228200
rect 219710 228188 219716 228200
rect 119212 228160 219716 228188
rect 119212 228148 119218 228160
rect 219710 228148 219716 228160
rect 219768 228148 219774 228200
rect 361574 228148 361580 228200
rect 361632 228188 361638 228200
rect 450722 228188 450728 228200
rect 361632 228160 450728 228188
rect 361632 228148 361638 228160
rect 450722 228148 450728 228160
rect 450780 228148 450786 228200
rect 97258 228080 97264 228132
rect 97316 228120 97322 228132
rect 210786 228120 210792 228132
rect 97316 228092 210792 228120
rect 97316 228080 97322 228092
rect 210786 228080 210792 228092
rect 210844 228080 210850 228132
rect 248782 228080 248788 228132
rect 248840 228120 248846 228132
rect 250070 228120 250076 228132
rect 248840 228092 250076 228120
rect 248840 228080 248846 228092
rect 250070 228080 250076 228092
rect 250128 228080 250134 228132
rect 362678 228080 362684 228132
rect 362736 228120 362742 228132
rect 452654 228120 452660 228132
rect 362736 228092 452660 228120
rect 362736 228080 362742 228092
rect 452654 228080 452660 228092
rect 452712 228080 452718 228132
rect 93762 228012 93768 228064
rect 93820 228052 93826 228064
rect 209406 228052 209412 228064
rect 93820 228024 209412 228052
rect 93820 228012 93826 228024
rect 209406 228012 209412 228024
rect 209464 228012 209470 228064
rect 221734 228012 221740 228064
rect 221792 228052 221798 228064
rect 263594 228052 263600 228064
rect 221792 228024 263600 228052
rect 221792 228012 221798 228024
rect 263594 228012 263600 228024
rect 263652 228012 263658 228064
rect 365530 228012 365536 228064
rect 365588 228052 365594 228064
rect 459186 228052 459192 228064
rect 365588 228024 459192 228052
rect 365588 228012 365594 228024
rect 459186 228012 459192 228024
rect 459244 228012 459250 228064
rect 87138 227944 87144 227996
rect 87196 227984 87202 227996
rect 206554 227984 206560 227996
rect 87196 227956 206560 227984
rect 87196 227944 87202 227956
rect 206554 227944 206560 227956
rect 206612 227944 206618 227996
rect 218330 227944 218336 227996
rect 218388 227984 218394 227996
rect 261846 227984 261852 227996
rect 218388 227956 261852 227984
rect 218388 227944 218394 227956
rect 261846 227944 261852 227956
rect 261904 227944 261910 227996
rect 364242 227944 364248 227996
rect 364300 227984 364306 227996
rect 455782 227984 455788 227996
rect 364300 227956 455788 227984
rect 364300 227944 364306 227956
rect 455782 227944 455788 227956
rect 455840 227944 455846 227996
rect 90542 227876 90548 227928
rect 90600 227916 90606 227928
rect 207934 227916 207940 227928
rect 90600 227888 207940 227916
rect 90600 227876 90606 227888
rect 207934 227876 207940 227888
rect 207992 227876 207998 227928
rect 215018 227876 215024 227928
rect 215076 227916 215082 227928
rect 260466 227916 260472 227928
rect 215076 227888 260472 227916
rect 215076 227876 215082 227888
rect 260466 227876 260472 227888
rect 260524 227876 260530 227928
rect 363966 227876 363972 227928
rect 364024 227916 364030 227928
rect 458358 227916 458364 227928
rect 364024 227888 458364 227916
rect 364024 227876 364030 227888
rect 458358 227876 458364 227888
rect 458416 227876 458422 227928
rect 61930 227808 61936 227860
rect 61988 227848 61994 227860
rect 195422 227848 195428 227860
rect 61988 227820 195428 227848
rect 61988 227808 61994 227820
rect 195422 227808 195428 227820
rect 195480 227808 195486 227860
rect 211706 227808 211712 227860
rect 211764 227848 211770 227860
rect 258994 227848 259000 227860
rect 211764 227820 259000 227848
rect 211764 227808 211770 227820
rect 258994 227808 259000 227820
rect 259052 227808 259058 227860
rect 368382 227808 368388 227860
rect 368440 227848 368446 227860
rect 465902 227848 465908 227860
rect 368440 227820 465908 227848
rect 368440 227808 368446 227820
rect 465902 227808 465908 227820
rect 465960 227808 465966 227860
rect 58618 227740 58624 227792
rect 58676 227780 58682 227792
rect 194042 227780 194048 227792
rect 58676 227752 194048 227780
rect 58676 227740 58682 227752
rect 194042 227740 194048 227752
rect 194100 227740 194106 227792
rect 204898 227740 204904 227792
rect 204956 227780 204962 227792
rect 256418 227780 256424 227792
rect 204956 227752 256424 227780
rect 204956 227740 204962 227752
rect 256418 227740 256424 227752
rect 256476 227740 256482 227792
rect 365162 227740 365168 227792
rect 365220 227780 365226 227792
rect 461670 227780 461676 227792
rect 365220 227752 461676 227780
rect 365220 227740 365226 227752
rect 461670 227740 461676 227752
rect 461728 227740 461734 227792
rect 53558 227672 53564 227724
rect 53616 227712 53622 227724
rect 192294 227712 192300 227724
rect 53616 227684 192300 227712
rect 53616 227672 53622 227684
rect 192294 227672 192300 227684
rect 192352 227672 192358 227724
rect 208486 227672 208492 227724
rect 208544 227712 208550 227724
rect 257890 227712 257896 227724
rect 208544 227684 257896 227712
rect 208544 227672 208550 227684
rect 257890 227672 257896 227684
rect 257948 227672 257954 227724
rect 366910 227672 366916 227724
rect 366968 227712 366974 227724
rect 462498 227712 462504 227724
rect 366968 227684 462504 227712
rect 366968 227672 366974 227684
rect 462498 227672 462504 227684
rect 462556 227672 462562 227724
rect 349798 227604 349804 227656
rect 349856 227644 349862 227656
rect 422294 227644 422300 227656
rect 349856 227616 422300 227644
rect 349856 227604 349862 227616
rect 422294 227604 422300 227616
rect 422352 227604 422358 227656
rect 351638 227536 351644 227588
rect 351696 227576 351702 227588
rect 427170 227576 427176 227588
rect 351696 227548 427176 227576
rect 351696 227536 351702 227548
rect 427170 227536 427176 227548
rect 427228 227536 427234 227588
rect 350166 227468 350172 227520
rect 350224 227508 350230 227520
rect 423858 227508 423864 227520
rect 350224 227480 423864 227508
rect 350224 227468 350230 227480
rect 423858 227468 423864 227480
rect 423916 227468 423922 227520
rect 42058 227400 42064 227452
rect 42116 227440 42122 227452
rect 43346 227440 43352 227452
rect 42116 227412 43352 227440
rect 42116 227400 42122 227412
rect 43346 227400 43352 227412
rect 43404 227400 43410 227452
rect 351270 227400 351276 227452
rect 351328 227440 351334 227452
rect 425514 227440 425520 227452
rect 351328 227412 425520 227440
rect 351328 227400 351334 227412
rect 425514 227400 425520 227412
rect 425572 227400 425578 227452
rect 348786 227332 348792 227384
rect 348844 227372 348850 227384
rect 420454 227372 420460 227384
rect 348844 227344 420460 227372
rect 348844 227332 348850 227344
rect 420454 227332 420460 227344
rect 420512 227332 420518 227384
rect 347682 227264 347688 227316
rect 347740 227304 347746 227316
rect 417142 227304 417148 227316
rect 347740 227276 417148 227304
rect 347740 227264 347746 227276
rect 417142 227264 417148 227276
rect 417200 227264 417206 227316
rect 345934 227196 345940 227248
rect 345992 227236 345998 227248
rect 414014 227236 414020 227248
rect 345992 227208 414020 227236
rect 345992 227196 345998 227208
rect 414014 227196 414020 227208
rect 414072 227196 414078 227248
rect 289998 227128 290004 227180
rect 290056 227168 290062 227180
rect 290734 227168 290740 227180
rect 290056 227140 290740 227168
rect 290056 227128 290062 227140
rect 290734 227128 290740 227140
rect 290792 227128 290798 227180
rect 348418 227128 348424 227180
rect 348476 227168 348482 227180
rect 418798 227168 418804 227180
rect 348476 227140 418804 227168
rect 348476 227128 348482 227140
rect 418798 227128 418804 227140
rect 418856 227128 418862 227180
rect 346946 227060 346952 227112
rect 347004 227100 347010 227112
rect 415394 227100 415400 227112
rect 347004 227072 415400 227100
rect 347004 227060 347010 227072
rect 415394 227060 415400 227072
rect 415452 227060 415458 227112
rect 344462 226992 344468 227044
rect 344520 227032 344526 227044
rect 410334 227032 410340 227044
rect 344520 227004 410340 227032
rect 344520 226992 344526 227004
rect 410334 226992 410340 227004
rect 410392 226992 410398 227044
rect 345566 226924 345572 226976
rect 345624 226964 345630 226976
rect 412082 226964 412088 226976
rect 345624 226936 412088 226964
rect 345624 226924 345630 226936
rect 412082 226924 412088 226936
rect 412140 226924 412146 226976
rect 344094 226856 344100 226908
rect 344152 226896 344158 226908
rect 408678 226896 408684 226908
rect 344152 226868 408684 226896
rect 344152 226856 344158 226868
rect 408678 226856 408684 226868
rect 408736 226856 408742 226908
rect 42150 226788 42156 226840
rect 42208 226828 42214 226840
rect 43806 226828 43812 226840
rect 42208 226800 43812 226828
rect 42208 226788 42214 226800
rect 43806 226788 43812 226800
rect 43864 226788 43870 226840
rect 342990 226788 342996 226840
rect 343048 226828 343054 226840
rect 405734 226828 405740 226840
rect 343048 226800 405740 226828
rect 343048 226788 343054 226800
rect 405734 226788 405740 226800
rect 405792 226788 405798 226840
rect 341242 226720 341248 226772
rect 341300 226760 341306 226772
rect 401962 226760 401968 226772
rect 341300 226732 401968 226760
rect 341300 226720 341306 226732
rect 401962 226720 401968 226732
rect 402020 226720 402026 226772
rect 339862 226652 339868 226704
rect 339920 226692 339926 226704
rect 398558 226692 398564 226704
rect 339920 226664 398564 226692
rect 339920 226652 339926 226664
rect 398558 226652 398564 226664
rect 398616 226652 398622 226704
rect 137646 226244 137652 226296
rect 137704 226284 137710 226296
rect 226610 226284 226616 226296
rect 137704 226256 226616 226284
rect 137704 226244 137710 226256
rect 226610 226244 226616 226256
rect 226668 226244 226674 226296
rect 349890 226244 349896 226296
rect 349948 226284 349954 226296
rect 421282 226284 421288 226296
rect 349948 226256 421288 226284
rect 349948 226244 349954 226256
rect 421282 226244 421288 226256
rect 421340 226244 421346 226296
rect 134242 226176 134248 226228
rect 134300 226216 134306 226228
rect 226518 226216 226524 226228
rect 134300 226188 226524 226216
rect 134300 226176 134306 226188
rect 226518 226176 226524 226188
rect 226576 226176 226582 226228
rect 347406 226176 347412 226228
rect 347464 226216 347470 226228
rect 418246 226216 418252 226228
rect 347464 226188 418252 226216
rect 347464 226176 347470 226188
rect 418246 226176 418252 226188
rect 418304 226176 418310 226228
rect 130930 226108 130936 226160
rect 130988 226148 130994 226160
rect 223758 226148 223764 226160
rect 130988 226120 223764 226148
rect 130988 226108 130994 226120
rect 223758 226108 223764 226120
rect 223816 226108 223822 226160
rect 347038 226108 347044 226160
rect 347096 226148 347102 226160
rect 419718 226148 419724 226160
rect 347096 226120 419724 226148
rect 347096 226108 347102 226120
rect 419718 226108 419724 226120
rect 419776 226108 419782 226160
rect 127526 226040 127532 226092
rect 127584 226080 127590 226092
rect 223850 226080 223856 226092
rect 127584 226052 223856 226080
rect 127584 226040 127590 226052
rect 223850 226040 223856 226052
rect 223908 226040 223914 226092
rect 352558 226040 352564 226092
rect 352616 226080 352622 226092
rect 426342 226080 426348 226092
rect 352616 226052 426348 226080
rect 352616 226040 352622 226052
rect 426342 226040 426348 226052
rect 426400 226040 426406 226092
rect 124122 225972 124128 226024
rect 124180 226012 124186 226024
rect 221090 226012 221096 226024
rect 124180 225984 221096 226012
rect 124180 225972 124186 225984
rect 221090 225972 221096 225984
rect 221148 225972 221154 226024
rect 350258 225972 350264 226024
rect 350316 226012 350322 226024
rect 423030 226012 423036 226024
rect 350316 225984 423036 226012
rect 350316 225972 350322 225984
rect 423030 225972 423036 225984
rect 423088 225972 423094 226024
rect 114094 225904 114100 225956
rect 114152 225944 114158 225956
rect 217594 225944 217600 225956
rect 114152 225916 217600 225944
rect 114152 225904 114158 225916
rect 217594 225904 217600 225916
rect 217652 225904 217658 225956
rect 352650 225904 352656 225956
rect 352708 225944 352714 225956
rect 429746 225944 429752 225956
rect 352708 225916 429752 225944
rect 352708 225904 352714 225916
rect 429746 225904 429752 225916
rect 429804 225904 429810 225956
rect 117498 225836 117504 225888
rect 117556 225876 117562 225888
rect 219066 225876 219072 225888
rect 117556 225848 219072 225876
rect 117556 225836 117562 225848
rect 219066 225836 219072 225848
rect 219124 225836 219130 225888
rect 353018 225836 353024 225888
rect 353076 225876 353082 225888
rect 427998 225876 428004 225888
rect 353076 225848 428004 225876
rect 353076 225836 353082 225848
rect 427998 225836 428004 225848
rect 428056 225836 428062 225888
rect 120810 225768 120816 225820
rect 120868 225808 120874 225820
rect 220998 225808 221004 225820
rect 120868 225780 221004 225808
rect 120868 225768 120874 225780
rect 220998 225768 221004 225780
rect 221056 225768 221062 225820
rect 350350 225768 350356 225820
rect 350408 225808 350414 225820
rect 425054 225808 425060 225820
rect 350408 225780 425060 225808
rect 350408 225768 350414 225780
rect 425054 225768 425060 225780
rect 425112 225768 425118 225820
rect 110690 225700 110696 225752
rect 110748 225740 110754 225752
rect 216214 225740 216220 225752
rect 110748 225712 216220 225740
rect 110748 225700 110754 225712
rect 216214 225700 216220 225712
rect 216272 225700 216278 225752
rect 355778 225700 355784 225752
rect 355836 225740 355842 225752
rect 433334 225740 433340 225752
rect 355836 225712 433340 225740
rect 355836 225700 355842 225712
rect 433334 225700 433340 225712
rect 433392 225700 433398 225752
rect 115750 225632 115756 225684
rect 115808 225672 115814 225684
rect 218238 225672 218244 225684
rect 115808 225644 218244 225672
rect 115808 225632 115814 225644
rect 218238 225632 218244 225644
rect 218296 225632 218302 225684
rect 355410 225632 355416 225684
rect 355468 225672 355474 225684
rect 434806 225672 434812 225684
rect 355468 225644 434812 225672
rect 355468 225632 355474 225644
rect 434806 225632 434812 225644
rect 434864 225632 434870 225684
rect 112438 225564 112444 225616
rect 112496 225604 112502 225616
rect 216582 225604 216588 225616
rect 112496 225576 216588 225604
rect 112496 225564 112502 225576
rect 216582 225564 216588 225576
rect 216640 225564 216646 225616
rect 352926 225564 352932 225616
rect 352984 225604 352990 225616
rect 431402 225604 431408 225616
rect 352984 225576 431408 225604
rect 352984 225564 352990 225576
rect 431402 225564 431408 225576
rect 431460 225564 431466 225616
rect 109034 225496 109040 225548
rect 109092 225536 109098 225548
rect 215662 225536 215668 225548
rect 109092 225508 215668 225536
rect 109092 225496 109098 225508
rect 215662 225496 215668 225508
rect 215720 225496 215726 225548
rect 355318 225496 355324 225548
rect 355376 225536 355382 225548
rect 438118 225536 438124 225548
rect 355376 225508 438124 225536
rect 355376 225496 355382 225508
rect 438118 225496 438124 225508
rect 438176 225496 438182 225548
rect 105722 225428 105728 225480
rect 105780 225468 105786 225480
rect 213730 225468 213736 225480
rect 105780 225440 213736 225468
rect 105780 225428 105786 225440
rect 213730 225428 213736 225440
rect 213788 225428 213794 225480
rect 358538 225428 358544 225480
rect 358596 225468 358602 225480
rect 439774 225468 439780 225480
rect 358596 225440 439780 225468
rect 358596 225428 358602 225440
rect 439774 225428 439780 225440
rect 439832 225428 439838 225480
rect 107378 225360 107384 225412
rect 107436 225400 107442 225412
rect 214834 225400 214840 225412
rect 107436 225372 214840 225400
rect 107436 225360 107442 225372
rect 214834 225360 214840 225372
rect 214892 225360 214898 225412
rect 355686 225360 355692 225412
rect 355744 225400 355750 225412
rect 436462 225400 436468 225412
rect 355744 225372 436468 225400
rect 355744 225360 355750 225372
rect 436462 225360 436468 225372
rect 436520 225360 436526 225412
rect 100662 225292 100668 225344
rect 100720 225332 100726 225344
rect 211982 225332 211988 225344
rect 100720 225304 211988 225332
rect 100720 225292 100726 225304
rect 211982 225292 211988 225304
rect 212040 225292 212046 225344
rect 228450 225292 228456 225344
rect 228508 225332 228514 225344
rect 266170 225332 266176 225344
rect 228508 225304 266176 225332
rect 228508 225292 228514 225304
rect 266170 225292 266176 225304
rect 266228 225292 266234 225344
rect 358078 225292 358084 225344
rect 358136 225332 358142 225344
rect 441614 225332 441620 225344
rect 358136 225304 441620 225332
rect 358136 225292 358142 225304
rect 441614 225292 441620 225304
rect 441672 225292 441678 225344
rect 103974 225224 103980 225276
rect 104032 225264 104038 225276
rect 213362 225264 213368 225276
rect 104032 225236 213368 225264
rect 104032 225224 104038 225236
rect 213362 225224 213368 225236
rect 213420 225224 213426 225276
rect 231762 225224 231768 225276
rect 231820 225264 231826 225276
rect 267826 225264 267832 225276
rect 231820 225236 267832 225264
rect 231820 225224 231826 225236
rect 267826 225224 267832 225236
rect 267884 225224 267890 225276
rect 361206 225224 361212 225276
rect 361264 225264 361270 225276
rect 446582 225264 446588 225276
rect 361264 225236 446588 225264
rect 361264 225224 361270 225236
rect 446582 225224 446588 225236
rect 446640 225224 446646 225276
rect 95602 225156 95608 225208
rect 95660 225196 95666 225208
rect 209498 225196 209504 225208
rect 95660 225168 209504 225196
rect 95660 225156 95666 225168
rect 209498 225156 209504 225168
rect 209556 225156 209562 225208
rect 225138 225156 225144 225208
rect 225196 225196 225202 225208
rect 265250 225196 265256 225208
rect 225196 225168 265256 225196
rect 225196 225156 225202 225168
rect 265250 225156 265256 225168
rect 265308 225156 265314 225208
rect 358446 225156 358452 225208
rect 358504 225196 358510 225208
rect 443178 225196 443184 225208
rect 358504 225168 443184 225196
rect 358504 225156 358510 225168
rect 443178 225156 443184 225168
rect 443236 225156 443242 225208
rect 73706 225088 73712 225140
rect 73764 225128 73770 225140
rect 200574 225128 200580 225140
rect 73764 225100 200580 225128
rect 73764 225088 73770 225100
rect 200574 225088 200580 225100
rect 200632 225088 200638 225140
rect 201310 225088 201316 225140
rect 201368 225128 201374 225140
rect 254762 225128 254768 225140
rect 201368 225100 254768 225128
rect 201368 225088 201374 225100
rect 254762 225088 254768 225100
rect 254820 225088 254826 225140
rect 358170 225088 358176 225140
rect 358228 225128 358234 225140
rect 444834 225128 444840 225140
rect 358228 225100 444840 225128
rect 358228 225088 358234 225100
rect 444834 225088 444840 225100
rect 444892 225088 444898 225140
rect 66990 225020 66996 225072
rect 67048 225060 67054 225072
rect 196434 225060 196440 225072
rect 67048 225032 196440 225060
rect 67048 225020 67054 225032
rect 196434 225020 196440 225032
rect 196492 225020 196498 225072
rect 198182 225020 198188 225072
rect 198240 225060 198246 225072
rect 251358 225060 251364 225072
rect 198240 225032 251364 225060
rect 198240 225020 198246 225032
rect 251358 225020 251364 225032
rect 251416 225020 251422 225072
rect 361390 225020 361396 225072
rect 361448 225060 361454 225072
rect 448238 225060 448244 225072
rect 361448 225032 448244 225060
rect 361448 225020 361454 225032
rect 448238 225020 448244 225032
rect 448296 225020 448302 225072
rect 60274 224952 60280 225004
rect 60332 224992 60338 225004
rect 193490 224992 193496 225004
rect 60332 224964 193496 224992
rect 60332 224952 60338 224964
rect 193490 224952 193496 224964
rect 193548 224952 193554 225004
rect 194870 224952 194876 225004
rect 194928 224992 194934 225004
rect 251910 224992 251916 225004
rect 194928 224964 251916 224992
rect 194928 224952 194934 224964
rect 251910 224952 251916 224964
rect 251968 224952 251974 225004
rect 363506 224952 363512 225004
rect 363564 224992 363570 225004
rect 453298 224992 453304 225004
rect 363564 224964 453304 224992
rect 363564 224952 363570 224964
rect 453298 224952 453304 224964
rect 453356 224952 453362 225004
rect 55122 224884 55128 224936
rect 55180 224924 55186 224936
rect 190638 224924 190644 224936
rect 55180 224896 190644 224924
rect 55180 224884 55186 224896
rect 190638 224884 190644 224896
rect 190696 224884 190702 224936
rect 191466 224884 191472 224936
rect 191524 224924 191530 224936
rect 248598 224924 248604 224936
rect 191524 224896 248604 224924
rect 191524 224884 191530 224896
rect 248598 224884 248604 224896
rect 248656 224884 248662 224936
rect 361298 224884 361304 224936
rect 361356 224924 361362 224936
rect 449894 224924 449900 224936
rect 361356 224896 449900 224924
rect 361356 224884 361362 224896
rect 449894 224884 449900 224896
rect 449952 224884 449958 224936
rect 141050 224816 141056 224868
rect 141108 224856 141114 224868
rect 229370 224856 229376 224868
rect 141108 224828 229376 224856
rect 141108 224816 141114 224828
rect 229370 224816 229376 224828
rect 229428 224816 229434 224868
rect 347590 224816 347596 224868
rect 347648 224856 347654 224868
rect 416222 224856 416228 224868
rect 347648 224828 416228 224856
rect 347648 224816 347654 224828
rect 416222 224816 416228 224828
rect 416280 224816 416286 224868
rect 144362 224748 144368 224800
rect 144420 224788 144426 224800
rect 229278 224788 229284 224800
rect 144420 224760 229284 224788
rect 144420 224748 144426 224760
rect 229278 224748 229284 224760
rect 229336 224748 229342 224800
rect 344830 224748 344836 224800
rect 344888 224788 344894 224800
rect 411254 224788 411260 224800
rect 344888 224760 411260 224788
rect 344888 224748 344894 224760
rect 411254 224748 411260 224760
rect 411312 224748 411318 224800
rect 147766 224680 147772 224732
rect 147824 224720 147830 224732
rect 232130 224720 232136 224732
rect 147824 224692 232136 224720
rect 147824 224680 147830 224692
rect 232130 224680 232136 224692
rect 232188 224680 232194 224732
rect 344738 224680 344744 224732
rect 344796 224720 344802 224732
rect 412910 224720 412916 224732
rect 344796 224692 412916 224720
rect 344796 224680 344802 224692
rect 412910 224680 412916 224692
rect 412968 224680 412974 224732
rect 154482 224612 154488 224664
rect 154540 224652 154546 224664
rect 234890 224652 234896 224664
rect 154540 224624 234896 224652
rect 154540 224612 154546 224624
rect 234890 224612 234896 224624
rect 234948 224612 234954 224664
rect 347130 224612 347136 224664
rect 347188 224652 347194 224664
rect 414566 224652 414572 224664
rect 347188 224624 414572 224652
rect 347188 224612 347194 224624
rect 414566 224612 414572 224624
rect 414624 224612 414630 224664
rect 151078 224544 151084 224596
rect 151136 224584 151142 224596
rect 232038 224584 232044 224596
rect 151136 224556 232044 224584
rect 151136 224544 151142 224556
rect 232038 224544 232044 224556
rect 232096 224544 232102 224596
rect 344646 224544 344652 224596
rect 344704 224584 344710 224596
rect 409506 224584 409512 224596
rect 344704 224556 409512 224584
rect 344704 224544 344710 224556
rect 409506 224544 409512 224556
rect 409564 224544 409570 224596
rect 161198 224476 161204 224528
rect 161256 224516 161262 224528
rect 237558 224516 237564 224528
rect 161256 224488 237564 224516
rect 161256 224476 161262 224488
rect 237558 224476 237564 224488
rect 237616 224476 237622 224528
rect 341886 224476 341892 224528
rect 341944 224516 341950 224528
rect 406194 224516 406200 224528
rect 341944 224488 406200 224516
rect 341944 224476 341950 224488
rect 406194 224476 406200 224488
rect 406252 224476 406258 224528
rect 703998 224476 704004 224528
rect 704056 224516 704062 224528
rect 708874 224516 708880 224528
rect 704056 224488 708880 224516
rect 704056 224476 704062 224488
rect 708874 224476 708880 224488
rect 708932 224476 708938 224528
rect 157794 224408 157800 224460
rect 157852 224448 157858 224460
rect 234798 224448 234804 224460
rect 157852 224420 234804 224448
rect 157852 224408 157858 224420
rect 234798 224408 234804 224420
rect 234856 224408 234862 224460
rect 341978 224408 341984 224460
rect 342036 224448 342042 224460
rect 402974 224448 402980 224460
rect 342036 224420 402980 224448
rect 342036 224408 342042 224420
rect 402974 224408 402980 224420
rect 403032 224408 403038 224460
rect 704458 224408 704464 224460
rect 704516 224448 704522 224460
rect 708414 224448 708420 224460
rect 704516 224420 708420 224448
rect 704516 224408 704522 224420
rect 708414 224408 708420 224420
rect 708472 224408 708478 224460
rect 164602 224340 164608 224392
rect 164660 224380 164666 224392
rect 237650 224380 237656 224392
rect 164660 224352 237656 224380
rect 164660 224340 164666 224352
rect 237650 224340 237656 224352
rect 237708 224340 237714 224392
rect 341150 224340 341156 224392
rect 341208 224380 341214 224392
rect 404446 224380 404452 224392
rect 341208 224352 404452 224380
rect 341208 224340 341214 224352
rect 404446 224340 404452 224352
rect 404504 224340 404510 224392
rect 707494 224380 707500 224392
rect 705304 224352 707500 224380
rect 167914 224272 167920 224324
rect 167972 224312 167978 224324
rect 240594 224312 240600 224324
rect 167972 224284 240600 224312
rect 167972 224272 167978 224284
rect 240594 224272 240600 224284
rect 240652 224272 240658 224324
rect 344370 224272 344376 224324
rect 344428 224312 344434 224324
rect 407850 224312 407856 224324
rect 344428 224284 407856 224312
rect 344428 224272 344434 224284
rect 407850 224272 407856 224284
rect 407908 224272 407914 224324
rect 705304 224256 705332 224352
rect 707494 224340 707500 224352
rect 707552 224340 707558 224392
rect 707034 224312 707040 224324
rect 705764 224284 707040 224312
rect 705764 224256 705792 224284
rect 707034 224272 707040 224284
rect 707092 224272 707098 224324
rect 171042 224204 171048 224256
rect 171100 224244 171106 224256
rect 240318 224244 240324 224256
rect 171100 224216 240324 224244
rect 171100 224204 171106 224216
rect 240318 224204 240324 224216
rect 240376 224204 240382 224256
rect 336274 224204 336280 224256
rect 336332 224244 336338 224256
rect 394694 224244 394700 224256
rect 336332 224216 394700 224244
rect 336332 224204 336338 224216
rect 394694 224204 394700 224216
rect 394752 224204 394758 224256
rect 705286 224204 705292 224256
rect 705344 224204 705350 224256
rect 705746 224204 705752 224256
rect 705804 224204 705810 224256
rect 706206 224204 706212 224256
rect 706264 224244 706270 224256
rect 706574 224244 706580 224256
rect 706264 224216 706580 224244
rect 706264 224204 706270 224216
rect 706574 224204 706580 224216
rect 706632 224204 706638 224256
rect 174630 224136 174636 224188
rect 174688 224176 174694 224188
rect 243446 224176 243452 224188
rect 174688 224148 243452 224176
rect 174688 224136 174694 224148
rect 243446 224136 243452 224148
rect 243504 224136 243510 224188
rect 339126 224136 339132 224188
rect 339184 224176 339190 224188
rect 397730 224176 397736 224188
rect 339184 224148 397736 224176
rect 339184 224136 339190 224148
rect 397730 224136 397736 224148
rect 397788 224136 397794 224188
rect 705838 224136 705844 224188
rect 705896 224176 705902 224188
rect 707034 224176 707040 224188
rect 705896 224148 707040 224176
rect 705896 224136 705902 224148
rect 707034 224136 707040 224148
rect 707092 224136 707098 224188
rect 178034 224068 178040 224120
rect 178092 224108 178098 224120
rect 243078 224108 243084 224120
rect 178092 224080 243084 224108
rect 178092 224068 178098 224080
rect 243078 224068 243084 224080
rect 243136 224068 243142 224120
rect 341794 224068 341800 224120
rect 341852 224108 341858 224120
rect 401134 224108 401140 224120
rect 341852 224080 401140 224108
rect 341852 224068 341858 224080
rect 401134 224068 401140 224080
rect 401192 224068 401198 224120
rect 706298 224068 706304 224120
rect 706356 224108 706362 224120
rect 706574 224108 706580 224120
rect 706356 224080 706580 224108
rect 706356 224068 706362 224080
rect 706574 224068 706580 224080
rect 706632 224068 706638 224120
rect 181346 224000 181352 224052
rect 181404 224040 181410 224052
rect 246206 224040 246212 224052
rect 181404 224012 246212 224040
rect 181404 224000 181410 224012
rect 246206 224000 246212 224012
rect 246264 224000 246270 224052
rect 336366 224000 336372 224052
rect 336424 224040 336430 224052
rect 391014 224040 391020 224052
rect 336424 224012 391020 224040
rect 336424 224000 336430 224012
rect 391014 224000 391020 224012
rect 391072 224000 391078 224052
rect 705378 224000 705384 224052
rect 705436 224040 705442 224052
rect 707494 224040 707500 224052
rect 705436 224012 707500 224040
rect 705436 224000 705442 224012
rect 707494 224000 707500 224012
rect 707552 224000 707558 224052
rect 708046 224000 708052 224052
rect 708104 224000 708110 224052
rect 184750 223932 184756 223984
rect 184808 223972 184814 223984
rect 245838 223972 245844 223984
rect 184808 223944 245844 223972
rect 184808 223932 184814 223944
rect 245838 223932 245844 223944
rect 245896 223932 245902 223984
rect 333422 223932 333428 223984
rect 333480 223972 333486 223984
rect 385954 223972 385960 223984
rect 333480 223944 385960 223972
rect 333480 223932 333486 223944
rect 385954 223932 385960 223944
rect 386012 223932 386018 223984
rect 704918 223932 704924 223984
rect 704976 223972 704982 223984
rect 707954 223972 707960 223984
rect 704976 223944 707960 223972
rect 704976 223932 704982 223944
rect 707954 223932 707960 223944
rect 708012 223932 708018 223984
rect 188154 223864 188160 223916
rect 188212 223904 188218 223916
rect 249058 223904 249064 223916
rect 188212 223876 249064 223904
rect 188212 223864 188218 223876
rect 249058 223864 249064 223876
rect 249116 223864 249122 223916
rect 333514 223864 333520 223916
rect 333572 223904 333578 223916
rect 382642 223904 382648 223916
rect 333572 223876 382648 223904
rect 333572 223864 333578 223876
rect 382642 223864 382648 223876
rect 382700 223864 382706 223916
rect 704826 223864 704832 223916
rect 704884 223904 704890 223916
rect 708064 223904 708092 224000
rect 704884 223876 708092 223904
rect 704884 223864 704890 223876
rect 113082 223524 113088 223576
rect 113140 223564 113146 223576
rect 139302 223564 139308 223576
rect 113140 223536 139308 223564
rect 113140 223524 113146 223536
rect 139302 223524 139308 223536
rect 139360 223524 139366 223576
rect 141878 223524 141884 223576
rect 141936 223564 141942 223576
rect 229186 223564 229192 223576
rect 141936 223536 229192 223564
rect 141936 223524 141942 223536
rect 229186 223524 229192 223536
rect 229244 223524 229250 223576
rect 272242 223524 272248 223576
rect 272300 223564 272306 223576
rect 284570 223564 284576 223576
rect 272300 223536 284576 223564
rect 272300 223524 272306 223536
rect 284570 223524 284576 223536
rect 284628 223524 284634 223576
rect 325510 223524 325516 223576
rect 325568 223564 325574 223576
rect 361758 223564 361764 223576
rect 325568 223536 361764 223564
rect 325568 223524 325574 223536
rect 361758 223524 361764 223536
rect 361816 223524 361822 223576
rect 494330 223524 494336 223576
rect 494388 223564 494394 223576
rect 495342 223564 495348 223576
rect 494388 223536 495348 223564
rect 494388 223524 494394 223536
rect 495342 223524 495348 223536
rect 495400 223564 495406 223576
rect 607582 223564 607588 223576
rect 495400 223536 607588 223564
rect 495400 223524 495406 223536
rect 607582 223524 607588 223536
rect 607640 223524 607646 223576
rect 108206 223456 108212 223508
rect 108264 223496 108270 223508
rect 136542 223496 136548 223508
rect 108264 223468 136548 223496
rect 108264 223456 108270 223468
rect 136542 223456 136548 223468
rect 136600 223456 136606 223508
rect 140130 223456 140136 223508
rect 140188 223496 140194 223508
rect 229738 223496 229744 223508
rect 140188 223468 229744 223496
rect 140188 223456 140194 223468
rect 229738 223456 229744 223468
rect 229796 223456 229802 223508
rect 230934 223456 230940 223508
rect 230992 223496 230998 223508
rect 244274 223496 244280 223508
rect 230992 223468 244280 223496
rect 230992 223456 230998 223468
rect 244274 223456 244280 223468
rect 244332 223456 244338 223508
rect 244458 223456 244464 223508
rect 244516 223456 244522 223508
rect 273070 223456 273076 223508
rect 273128 223496 273134 223508
rect 284754 223496 284760 223508
rect 273128 223468 284760 223496
rect 273128 223456 273134 223468
rect 284754 223456 284760 223468
rect 284812 223456 284818 223508
rect 325142 223456 325148 223508
rect 325200 223496 325206 223508
rect 362402 223496 362408 223508
rect 325200 223468 362408 223496
rect 325200 223456 325206 223468
rect 362402 223456 362408 223468
rect 362460 223456 362466 223508
rect 499482 223456 499488 223508
rect 499540 223496 499546 223508
rect 608042 223496 608048 223508
rect 499540 223468 608048 223496
rect 499540 223456 499546 223468
rect 608042 223456 608048 223468
rect 608100 223456 608106 223508
rect 106550 223388 106556 223440
rect 106608 223428 106614 223440
rect 125502 223428 125508 223440
rect 106608 223400 125508 223428
rect 106608 223388 106614 223400
rect 125502 223388 125508 223400
rect 125560 223388 125566 223440
rect 135162 223388 135168 223440
rect 135220 223428 135226 223440
rect 226794 223428 226800 223440
rect 135220 223400 226800 223428
rect 135220 223388 135226 223400
rect 226794 223388 226800 223400
rect 226852 223388 226858 223440
rect 227530 223388 227536 223440
rect 227588 223428 227594 223440
rect 244476 223428 244504 223456
rect 227588 223400 244504 223428
rect 227588 223388 227594 223400
rect 278682 223388 278688 223440
rect 278740 223428 278746 223440
rect 287330 223428 287336 223440
rect 278740 223400 287336 223428
rect 278740 223388 278746 223400
rect 287330 223388 287336 223400
rect 287388 223388 287394 223440
rect 314194 223388 314200 223440
rect 314252 223428 314258 223440
rect 339678 223428 339684 223440
rect 314252 223400 339684 223428
rect 314252 223388 314258 223400
rect 339678 223388 339684 223400
rect 339736 223388 339742 223440
rect 346210 223388 346216 223440
rect 346268 223428 346274 223440
rect 383654 223428 383660 223440
rect 346268 223400 383660 223428
rect 346268 223388 346274 223400
rect 383654 223388 383660 223400
rect 383712 223388 383718 223440
rect 403802 223388 403808 223440
rect 403860 223428 403866 223440
rect 539042 223428 539048 223440
rect 403860 223400 539048 223428
rect 403860 223388 403866 223400
rect 539042 223388 539048 223400
rect 539100 223388 539106 223440
rect 546034 223388 546040 223440
rect 546092 223428 546098 223440
rect 616874 223428 616880 223440
rect 546092 223400 616880 223428
rect 546092 223388 546098 223400
rect 616874 223388 616880 223400
rect 616932 223388 616938 223440
rect 86310 223320 86316 223372
rect 86368 223360 86374 223372
rect 128262 223360 128268 223372
rect 86368 223332 128268 223360
rect 86368 223320 86374 223332
rect 128262 223320 128268 223332
rect 128320 223320 128326 223372
rect 198706 223332 198964 223360
rect 101490 223252 101496 223304
rect 101548 223292 101554 223304
rect 122742 223292 122748 223304
rect 101548 223264 122748 223292
rect 101548 223252 101554 223264
rect 122742 223252 122748 223264
rect 122800 223252 122806 223304
rect 128354 223252 128360 223304
rect 128412 223292 128418 223304
rect 198706 223292 198734 223332
rect 128412 223264 198734 223292
rect 198936 223292 198964 223332
rect 199010 223320 199016 223372
rect 199068 223360 199074 223372
rect 224126 223360 224132 223372
rect 199068 223332 224132 223360
rect 199068 223320 199074 223332
rect 224126 223320 224132 223332
rect 224184 223320 224190 223372
rect 229278 223320 229284 223372
rect 229336 223360 229342 223372
rect 244182 223360 244188 223372
rect 229336 223332 244188 223360
rect 229336 223320 229342 223332
rect 244182 223320 244188 223332
rect 244240 223320 244246 223372
rect 244458 223320 244464 223372
rect 244516 223360 244522 223372
rect 255314 223360 255320 223372
rect 244516 223332 255320 223360
rect 244516 223320 244522 223332
rect 255314 223320 255320 223332
rect 255372 223320 255378 223372
rect 278130 223320 278136 223372
rect 278188 223360 278194 223372
rect 287146 223360 287152 223372
rect 278188 223332 287152 223360
rect 278188 223320 278194 223332
rect 287146 223320 287152 223332
rect 287204 223320 287210 223372
rect 328178 223320 328184 223372
rect 328236 223360 328242 223372
rect 369118 223360 369124 223372
rect 328236 223332 369124 223360
rect 328236 223320 328242 223332
rect 369118 223320 369124 223332
rect 369176 223320 369182 223372
rect 500862 223320 500868 223372
rect 500920 223360 500926 223372
rect 608502 223360 608508 223372
rect 500920 223332 608508 223360
rect 500920 223320 500926 223332
rect 608502 223320 608508 223332
rect 608560 223320 608566 223372
rect 224034 223292 224040 223304
rect 198936 223264 224040 223292
rect 128412 223252 128418 223264
rect 224034 223252 224040 223264
rect 224092 223252 224098 223304
rect 241146 223252 241152 223304
rect 241204 223292 241210 223304
rect 252554 223292 252560 223304
rect 241204 223264 252560 223292
rect 241204 223252 241210 223264
rect 252554 223252 252560 223264
rect 252612 223252 252618 223304
rect 328270 223252 328276 223304
rect 328328 223292 328334 223304
rect 368290 223292 368296 223304
rect 328328 223264 368296 223292
rect 328328 223252 328334 223264
rect 368290 223252 368296 223264
rect 368348 223252 368354 223304
rect 394510 223252 394516 223304
rect 394568 223292 394574 223304
rect 530026 223292 530032 223304
rect 394568 223264 530032 223292
rect 394568 223252 394574 223264
rect 530026 223252 530032 223264
rect 530084 223252 530090 223304
rect 538858 223252 538864 223304
rect 538916 223292 538922 223304
rect 539594 223292 539600 223304
rect 538916 223264 539600 223292
rect 538916 223252 538922 223264
rect 539594 223252 539600 223264
rect 539652 223292 539658 223304
rect 539652 223264 546908 223292
rect 539652 223252 539658 223264
rect 78766 223184 78772 223236
rect 78824 223224 78830 223236
rect 119982 223224 119988 223236
rect 78824 223196 119988 223224
rect 78824 223184 78830 223196
rect 119982 223184 119988 223196
rect 120040 223184 120046 223236
rect 126698 223184 126704 223236
rect 126756 223224 126762 223236
rect 198826 223224 198832 223236
rect 126756 223196 198832 223224
rect 126756 223184 126762 223196
rect 198826 223184 198832 223196
rect 198884 223184 198890 223236
rect 198918 223184 198924 223236
rect 198976 223224 198982 223236
rect 207934 223224 207940 223236
rect 198976 223196 207940 223224
rect 198976 223184 198982 223196
rect 207934 223184 207940 223196
rect 207992 223184 207998 223236
rect 215294 223224 215300 223236
rect 208228 223196 215300 223224
rect 94774 223116 94780 223168
rect 94832 223156 94838 223168
rect 111702 223156 111708 223168
rect 94832 223128 111708 223156
rect 94832 223116 94838 223128
rect 111702 223116 111708 223128
rect 111760 223116 111766 223168
rect 116578 223116 116584 223168
rect 116636 223156 116642 223168
rect 208228 223156 208256 223196
rect 215294 223184 215300 223196
rect 215352 223184 215358 223236
rect 221274 223224 221280 223236
rect 218026 223196 221280 223224
rect 218026 223156 218054 223196
rect 221274 223184 221280 223196
rect 221332 223184 221338 223236
rect 237742 223184 237748 223236
rect 237800 223224 237806 223236
rect 252462 223224 252468 223236
rect 237800 223196 252468 223224
rect 237800 223184 237806 223196
rect 252462 223184 252468 223196
rect 252520 223184 252526 223236
rect 325602 223184 325608 223236
rect 325660 223224 325666 223236
rect 365806 223224 365812 223236
rect 325660 223196 365812 223224
rect 325660 223184 325666 223196
rect 365806 223184 365812 223196
rect 365864 223184 365870 223236
rect 398650 223184 398656 223236
rect 398708 223224 398714 223236
rect 539870 223224 539876 223236
rect 398708 223196 539876 223224
rect 398708 223184 398714 223196
rect 539870 223184 539876 223196
rect 539928 223184 539934 223236
rect 542446 223184 542452 223236
rect 542504 223224 542510 223236
rect 543642 223224 543648 223236
rect 542504 223196 543648 223224
rect 542504 223184 542510 223196
rect 543642 223184 543648 223196
rect 543700 223224 543706 223236
rect 546880 223224 546908 223264
rect 546954 223252 546960 223304
rect 547012 223292 547018 223304
rect 615034 223292 615040 223304
rect 547012 223264 615040 223292
rect 547012 223252 547018 223264
rect 615034 223252 615040 223264
rect 615092 223252 615098 223304
rect 615494 223224 615500 223236
rect 543700 223196 546816 223224
rect 546880 223196 615500 223224
rect 543700 223184 543706 223196
rect 116636 223128 208256 223156
rect 208320 223128 218054 223156
rect 116636 223116 116642 223128
rect 72050 223048 72056 223100
rect 72108 223088 72114 223100
rect 117222 223088 117228 223100
rect 72108 223060 117228 223088
rect 72108 223048 72114 223060
rect 117222 223048 117228 223060
rect 117280 223048 117286 223100
rect 119982 223048 119988 223100
rect 120040 223088 120046 223100
rect 208320 223088 208348 223128
rect 220078 223116 220084 223168
rect 220136 223156 220142 223168
rect 235902 223156 235908 223168
rect 220136 223128 235908 223156
rect 220136 223116 220142 223128
rect 235902 223116 235908 223128
rect 235960 223116 235966 223168
rect 242710 223116 242716 223168
rect 242768 223156 242774 223168
rect 255498 223156 255504 223168
rect 242768 223128 255504 223156
rect 242768 223116 242774 223128
rect 255498 223116 255504 223128
rect 255556 223116 255562 223168
rect 308950 223116 308956 223168
rect 309008 223156 309014 223168
rect 323118 223156 323124 223168
rect 309008 223128 323124 223156
rect 309008 223116 309014 223128
rect 323118 223116 323124 223128
rect 323176 223116 323182 223168
rect 325418 223116 325424 223168
rect 325476 223156 325482 223168
rect 364978 223156 364984 223168
rect 325476 223128 364984 223156
rect 325476 223116 325482 223128
rect 364978 223116 364984 223128
rect 365036 223116 365042 223168
rect 406378 223116 406384 223168
rect 406436 223156 406442 223168
rect 546678 223156 546684 223168
rect 406436 223128 546684 223156
rect 406436 223116 406442 223128
rect 546678 223116 546684 223128
rect 546736 223116 546742 223168
rect 546788 223156 546816 223196
rect 615494 223184 615500 223196
rect 615552 223184 615558 223236
rect 616414 223156 616420 223168
rect 546788 223128 616420 223156
rect 616414 223116 616420 223128
rect 616472 223116 616478 223168
rect 218422 223088 218428 223100
rect 120040 223060 208348 223088
rect 218026 223060 218428 223088
rect 120040 223048 120046 223060
rect 88058 222980 88064 223032
rect 88116 223020 88122 223032
rect 106182 223020 106188 223032
rect 88116 222992 106188 223020
rect 88116 222980 88122 222992
rect 106182 222980 106188 222992
rect 106240 222980 106246 223032
rect 118326 222980 118332 223032
rect 118384 223020 118390 223032
rect 218026 223020 218054 223060
rect 218422 223048 218428 223060
rect 218480 223048 218486 223100
rect 226610 223048 226616 223100
rect 226668 223088 226674 223100
rect 230934 223088 230940 223100
rect 226668 223060 230940 223088
rect 226668 223048 226674 223060
rect 230934 223048 230940 223060
rect 230992 223048 230998 223100
rect 231026 223048 231032 223100
rect 231084 223088 231090 223100
rect 249886 223088 249892 223100
rect 231084 223060 249892 223088
rect 231084 223048 231090 223060
rect 249886 223048 249892 223060
rect 249944 223048 249950 223100
rect 311710 223048 311716 223100
rect 311768 223088 311774 223100
rect 330478 223088 330484 223100
rect 311768 223060 330484 223088
rect 311768 223048 311774 223060
rect 330478 223048 330484 223060
rect 330536 223048 330542 223100
rect 330846 223048 330852 223100
rect 330904 223088 330910 223100
rect 371694 223088 371700 223100
rect 330904 223060 371700 223088
rect 330904 223048 330910 223060
rect 371694 223048 371700 223060
rect 371752 223048 371758 223100
rect 400030 223048 400036 223100
rect 400088 223088 400094 223100
rect 542170 223088 542176 223100
rect 400088 223060 542176 223088
rect 400088 223048 400094 223060
rect 542170 223048 542176 223060
rect 542228 223048 542234 223100
rect 542354 223048 542360 223100
rect 542412 223088 542418 223100
rect 615954 223088 615960 223100
rect 542412 223060 615960 223088
rect 542412 223048 542418 223060
rect 615954 223048 615960 223060
rect 616012 223048 616018 223100
rect 118384 222992 218054 223020
rect 118384 222980 118390 222992
rect 224310 222980 224316 223032
rect 224368 223020 224374 223032
rect 250162 223020 250168 223032
rect 224368 222992 250168 223020
rect 224368 222980 224374 222992
rect 250162 222980 250168 222992
rect 250220 222980 250226 223032
rect 308766 222980 308772 223032
rect 308824 223020 308830 223032
rect 323762 223020 323768 223032
rect 308824 222992 323768 223020
rect 308824 222980 308830 222992
rect 323762 222980 323768 222992
rect 323820 222980 323826 223032
rect 325326 222980 325332 223032
rect 325384 223020 325390 223032
rect 364334 223020 364340 223032
rect 325384 222992 364340 223020
rect 325384 222980 325390 222992
rect 364334 222980 364340 222992
rect 364392 222980 364398 223032
rect 401870 222980 401876 223032
rect 401928 223020 401934 223032
rect 544930 223020 544936 223032
rect 401928 222992 544936 223020
rect 401928 222980 401934 222992
rect 544930 222980 544936 222992
rect 544988 222980 544994 223032
rect 545114 222980 545120 223032
rect 545172 223020 545178 223032
rect 546034 223020 546040 223032
rect 545172 222992 546040 223020
rect 545172 222980 545178 222992
rect 546034 222980 546040 222992
rect 546092 222980 546098 223032
rect 65334 222912 65340 222964
rect 65392 222952 65398 222964
rect 103422 222952 103428 222964
rect 65392 222924 103428 222952
rect 65392 222912 65398 222924
rect 103422 222912 103428 222924
rect 103480 222912 103486 222964
rect 109862 222912 109868 222964
rect 109920 222952 109926 222964
rect 198918 222952 198924 222964
rect 109920 222924 198924 222952
rect 109920 222912 109926 222924
rect 198918 222912 198924 222924
rect 198976 222912 198982 222964
rect 199010 222912 199016 222964
rect 199068 222952 199074 222964
rect 201402 222952 201408 222964
rect 199068 222924 201408 222952
rect 199068 222912 199074 222924
rect 201402 222912 201408 222924
rect 201460 222912 201466 222964
rect 207934 222912 207940 222964
rect 207992 222952 207998 222964
rect 212534 222952 212540 222964
rect 207992 222924 212540 222952
rect 207992 222912 207998 222924
rect 212534 222912 212540 222924
rect 212592 222912 212598 222964
rect 229370 222912 229376 222964
rect 229428 222952 229434 222964
rect 229428 222924 236040 222952
rect 229428 222912 229434 222924
rect 82722 222844 82728 222896
rect 82780 222884 82786 222896
rect 97902 222884 97908 222896
rect 82780 222856 97908 222884
rect 82780 222844 82786 222856
rect 97902 222844 97908 222856
rect 97960 222844 97966 222896
rect 103146 222844 103152 222896
rect 103204 222884 103210 222896
rect 214098 222884 214104 222896
rect 103204 222856 214104 222884
rect 103204 222844 103210 222856
rect 214098 222844 214104 222856
rect 214156 222844 214162 222896
rect 214190 222844 214196 222896
rect 214248 222884 214254 222896
rect 236012 222884 236040 222924
rect 236086 222912 236092 222964
rect 236144 222952 236150 222964
rect 268194 222952 268200 222964
rect 236144 222924 268200 222952
rect 236144 222912 236150 222924
rect 268194 222912 268200 222924
rect 268252 222912 268258 222964
rect 317230 222912 317236 222964
rect 317288 222952 317294 222964
rect 347314 222952 347320 222964
rect 317288 222924 347320 222952
rect 317288 222912 317294 222924
rect 347314 222912 347320 222924
rect 347372 222912 347378 222964
rect 347406 222912 347412 222964
rect 347464 222952 347470 222964
rect 386782 222952 386788 222964
rect 347464 222924 386788 222952
rect 347464 222912 347470 222924
rect 386782 222912 386788 222924
rect 386840 222912 386846 222964
rect 402514 222912 402520 222964
rect 402572 222952 402578 222964
rect 536282 222952 536288 222964
rect 402572 222924 536288 222952
rect 402572 222912 402578 222924
rect 536282 222912 536288 222924
rect 536340 222912 536346 222964
rect 536374 222912 536380 222964
rect 536432 222952 536438 222964
rect 536834 222952 536840 222964
rect 536432 222924 536840 222952
rect 536432 222912 536438 222924
rect 536834 222912 536840 222924
rect 536892 222952 536898 222964
rect 546954 222952 546960 222964
rect 536892 222924 546960 222952
rect 536892 222912 536898 222924
rect 546954 222912 546960 222924
rect 547012 222912 547018 222964
rect 550542 222912 550548 222964
rect 550600 222952 550606 222964
rect 551462 222952 551468 222964
rect 550600 222924 551468 222952
rect 550600 222912 550606 222924
rect 551462 222912 551468 222924
rect 551520 222952 551526 222964
rect 617794 222952 617800 222964
rect 551520 222924 617800 222952
rect 551520 222912 551526 222924
rect 617794 222912 617800 222924
rect 617852 222912 617858 222964
rect 263502 222884 263508 222896
rect 214248 222856 235948 222884
rect 236012 222856 263508 222884
rect 214248 222844 214254 222856
rect 98086 222776 98092 222828
rect 98144 222816 98150 222828
rect 211614 222816 211620 222828
rect 98144 222788 211620 222816
rect 98144 222776 98150 222788
rect 211614 222776 211620 222788
rect 211672 222776 211678 222828
rect 215846 222776 215852 222828
rect 215904 222816 215910 222828
rect 235810 222816 235816 222828
rect 215904 222788 235816 222816
rect 215904 222776 215910 222788
rect 235810 222776 235816 222788
rect 235868 222776 235874 222828
rect 235920 222816 235948 222856
rect 263502 222844 263508 222856
rect 263560 222844 263566 222896
rect 309042 222844 309048 222896
rect 309100 222884 309106 222896
rect 326246 222884 326252 222896
rect 309100 222856 326252 222884
rect 309100 222844 309106 222856
rect 326246 222844 326252 222856
rect 326304 222844 326310 222896
rect 328362 222844 328368 222896
rect 328420 222884 328426 222896
rect 370038 222884 370044 222896
rect 328420 222856 370044 222884
rect 328420 222844 328426 222856
rect 370038 222844 370044 222856
rect 370096 222844 370102 222896
rect 407390 222844 407396 222896
rect 407448 222884 407454 222896
rect 552014 222884 552020 222896
rect 407448 222856 552020 222884
rect 407448 222844 407454 222856
rect 552014 222844 552020 222856
rect 552072 222844 552078 222896
rect 557902 222884 557908 222896
rect 555160 222856 557908 222884
rect 247310 222816 247316 222828
rect 235920 222788 247316 222816
rect 247310 222776 247316 222788
rect 247368 222776 247374 222828
rect 308674 222776 308680 222828
rect 308732 222816 308738 222828
rect 324590 222816 324596 222828
rect 308732 222788 324596 222816
rect 308732 222776 308738 222788
rect 324590 222776 324596 222788
rect 324648 222776 324654 222828
rect 325234 222776 325240 222828
rect 325292 222816 325298 222828
rect 367462 222816 367468 222828
rect 325292 222788 367468 222816
rect 325292 222776 325298 222788
rect 367462 222776 367468 222788
rect 367520 222776 367526 222828
rect 405826 222776 405832 222828
rect 405884 222816 405890 222828
rect 405884 222788 554774 222816
rect 405884 222776 405890 222788
rect 62758 222708 62764 222760
rect 62816 222748 62822 222760
rect 89622 222748 89628 222760
rect 62816 222720 89628 222748
rect 62816 222708 62822 222720
rect 89622 222708 89628 222720
rect 89680 222708 89686 222760
rect 189534 222708 189540 222760
rect 189592 222748 189598 222760
rect 205174 222748 205180 222760
rect 189592 222720 205180 222748
rect 189592 222708 189598 222720
rect 205174 222708 205180 222720
rect 205232 222708 205238 222760
rect 207382 222708 207388 222760
rect 207440 222748 207446 222760
rect 247126 222748 247132 222760
rect 207440 222720 247132 222748
rect 207440 222708 207446 222720
rect 247126 222708 247132 222720
rect 247184 222708 247190 222760
rect 281442 222708 281448 222760
rect 281500 222748 281506 222760
rect 289906 222748 289912 222760
rect 281500 222720 289912 222748
rect 281500 222708 281506 222720
rect 289906 222708 289912 222720
rect 289964 222708 289970 222760
rect 308858 222708 308864 222760
rect 308916 222748 308922 222760
rect 327074 222748 327080 222760
rect 308916 222720 327080 222748
rect 308916 222708 308922 222720
rect 327074 222708 327080 222720
rect 327132 222708 327138 222760
rect 327902 222708 327908 222760
rect 327960 222748 327966 222760
rect 370866 222748 370872 222760
rect 327960 222720 370872 222748
rect 327960 222708 327966 222720
rect 370866 222708 370872 222720
rect 370924 222708 370930 222760
rect 404354 222708 404360 222760
rect 404412 222748 404418 222760
rect 552198 222748 552204 222760
rect 404412 222720 552204 222748
rect 404412 222708 404418 222720
rect 552198 222708 552204 222720
rect 552256 222708 552262 222760
rect 554746 222748 554774 222788
rect 555050 222748 555056 222760
rect 554746 222720 555056 222748
rect 555050 222708 555056 222720
rect 555108 222708 555114 222760
rect 71222 222640 71228 222692
rect 71280 222680 71286 222692
rect 81342 222680 81348 222692
rect 71280 222652 81348 222680
rect 71280 222640 71286 222652
rect 81342 222640 81348 222652
rect 81400 222640 81406 222692
rect 89714 222640 89720 222692
rect 89772 222680 89778 222692
rect 208394 222680 208400 222692
rect 89772 222652 208400 222680
rect 89772 222640 89778 222652
rect 208394 222640 208400 222652
rect 208452 222640 208458 222692
rect 222562 222640 222568 222692
rect 222620 222680 222626 222692
rect 262582 222680 262588 222692
rect 222620 222652 262588 222680
rect 222620 222640 222626 222652
rect 262582 222640 262588 222652
rect 262640 222640 262646 222692
rect 311434 222640 311440 222692
rect 311492 222680 311498 222692
rect 329650 222680 329656 222692
rect 311492 222652 329656 222680
rect 311492 222640 311498 222652
rect 329650 222640 329656 222652
rect 329708 222640 329714 222692
rect 333790 222640 333796 222692
rect 333848 222680 333854 222692
rect 378410 222680 378416 222692
rect 333848 222652 378416 222680
rect 333848 222640 333854 222652
rect 378410 222640 378416 222652
rect 378468 222640 378474 222692
rect 403986 222640 403992 222692
rect 404044 222680 404050 222692
rect 552106 222680 552112 222692
rect 404044 222652 552112 222680
rect 404044 222640 404050 222652
rect 552106 222640 552112 222652
rect 552164 222640 552170 222692
rect 82170 222572 82176 222624
rect 82228 222612 82234 222624
rect 203794 222612 203800 222624
rect 82228 222584 203800 222612
rect 82228 222572 82234 222584
rect 203794 222572 203800 222584
rect 203852 222572 203858 222624
rect 209130 222572 209136 222624
rect 209188 222612 209194 222624
rect 209188 222584 226334 222612
rect 209188 222572 209194 222584
rect 85482 222504 85488 222556
rect 85540 222544 85546 222556
rect 189534 222544 189540 222556
rect 85540 222516 189540 222544
rect 85540 222504 85546 222516
rect 189534 222504 189540 222516
rect 189592 222504 189598 222556
rect 204438 222544 204444 222556
rect 189644 222516 204444 222544
rect 81250 222436 81256 222488
rect 81308 222476 81314 222488
rect 189644 222476 189672 222516
rect 204438 222504 204444 222516
rect 204496 222504 204502 222556
rect 212350 222504 212356 222556
rect 212408 222544 212414 222556
rect 226306 222544 226334 222584
rect 235810 222572 235816 222624
rect 235868 222612 235874 222624
rect 259822 222612 259828 222624
rect 235868 222584 259828 222612
rect 235868 222572 235874 222584
rect 259822 222572 259828 222584
rect 259880 222572 259886 222624
rect 308490 222572 308496 222624
rect 308548 222612 308554 222624
rect 325694 222612 325700 222624
rect 308548 222584 325700 222612
rect 308548 222572 308554 222584
rect 325694 222572 325700 222584
rect 325752 222572 325758 222624
rect 327994 222572 328000 222624
rect 328052 222612 328058 222624
rect 372614 222612 372620 222624
rect 328052 222584 372620 222612
rect 328052 222572 328058 222584
rect 372614 222572 372620 222584
rect 372672 222572 372678 222624
rect 406286 222572 406292 222624
rect 406344 222612 406350 222624
rect 555160 222612 555188 222856
rect 557902 222844 557908 222856
rect 557960 222884 557966 222896
rect 564066 222884 564072 222896
rect 557960 222856 564072 222884
rect 557960 222844 557966 222856
rect 564066 222844 564072 222856
rect 564124 222844 564130 222896
rect 559098 222776 559104 222828
rect 559156 222816 559162 222828
rect 572806 222816 572812 222828
rect 559156 222788 572812 222816
rect 559156 222776 559162 222788
rect 572806 222776 572812 222788
rect 572864 222776 572870 222828
rect 559116 222748 559144 222776
rect 406344 222584 555188 222612
rect 555252 222720 559144 222748
rect 406344 222572 406350 222584
rect 257062 222544 257068 222556
rect 212408 222516 220952 222544
rect 226306 222516 257068 222544
rect 212408 222504 212414 222516
rect 81308 222448 189672 222476
rect 81308 222436 81314 222448
rect 189718 222436 189724 222488
rect 189776 222476 189782 222488
rect 208762 222476 208768 222488
rect 189776 222448 208768 222476
rect 189776 222436 189782 222448
rect 208762 222436 208768 222448
rect 208820 222436 208826 222488
rect 213362 222436 213368 222488
rect 213420 222476 213426 222488
rect 220814 222476 220820 222488
rect 213420 222448 220820 222476
rect 213420 222436 213426 222448
rect 220814 222436 220820 222448
rect 220872 222436 220878 222488
rect 220924 222476 220952 222516
rect 257062 222504 257068 222516
rect 257120 222504 257126 222556
rect 311526 222504 311532 222556
rect 311584 222544 311590 222556
rect 332962 222544 332968 222556
rect 311584 222516 332968 222544
rect 311584 222504 311590 222516
rect 332962 222504 332968 222516
rect 333020 222504 333026 222556
rect 333882 222504 333888 222556
rect 333940 222544 333946 222556
rect 381814 222544 381820 222556
rect 333940 222516 381820 222544
rect 333940 222504 333946 222516
rect 381814 222504 381820 222516
rect 381872 222504 381878 222556
rect 406470 222504 406476 222556
rect 406528 222544 406534 222556
rect 555252 222544 555280 222720
rect 561674 222708 561680 222760
rect 561732 222748 561738 222760
rect 619634 222748 619640 222760
rect 561732 222720 619640 222748
rect 561732 222708 561738 222720
rect 619634 222708 619640 222720
rect 619692 222708 619698 222760
rect 556062 222640 556068 222692
rect 556120 222680 556126 222692
rect 618714 222680 618720 222692
rect 556120 222652 618720 222680
rect 556120 222640 556126 222652
rect 618714 222640 618720 222652
rect 618772 222640 618778 222692
rect 563974 222612 563980 222624
rect 406528 222516 555280 222544
rect 555344 222584 563980 222612
rect 406528 222504 406534 222516
rect 260098 222476 260104 222488
rect 220924 222448 260104 222476
rect 260098 222436 260104 222448
rect 260156 222436 260162 222488
rect 311342 222436 311348 222488
rect 311400 222476 311406 222488
rect 331306 222476 331312 222488
rect 311400 222448 331312 222476
rect 311400 222436 311406 222448
rect 331306 222436 331312 222448
rect 331364 222436 331370 222488
rect 336090 222436 336096 222488
rect 336148 222476 336154 222488
rect 385126 222476 385132 222488
rect 336148 222448 385132 222476
rect 336148 222436 336154 222448
rect 385126 222436 385132 222448
rect 385184 222436 385190 222488
rect 408770 222436 408776 222488
rect 408828 222476 408834 222488
rect 555344 222476 555372 222584
rect 563974 222572 563980 222584
rect 564032 222572 564038 222624
rect 564066 222572 564072 222624
rect 564124 222612 564130 222624
rect 633618 222612 633624 222624
rect 564124 222584 633624 222612
rect 564124 222572 564130 222584
rect 633618 222572 633624 222584
rect 633676 222572 633682 222624
rect 561582 222504 561588 222556
rect 561640 222544 561646 222556
rect 634078 222544 634084 222556
rect 561640 222516 634084 222544
rect 561640 222504 561646 222516
rect 634078 222504 634084 222516
rect 634136 222504 634142 222556
rect 408828 222448 555372 222476
rect 408828 222436 408834 222448
rect 555418 222436 555424 222488
rect 555476 222476 555482 222488
rect 562870 222476 562876 222488
rect 555476 222448 562876 222476
rect 555476 222436 555482 222448
rect 562870 222436 562876 222448
rect 562928 222436 562934 222488
rect 563974 222436 563980 222488
rect 564032 222476 564038 222488
rect 620094 222476 620100 222488
rect 564032 222448 620100 222476
rect 564032 222436 564038 222448
rect 620094 222436 620100 222448
rect 620152 222436 620158 222488
rect 56042 222368 56048 222420
rect 56100 222408 56106 222420
rect 73062 222408 73068 222420
rect 56100 222380 73068 222408
rect 56100 222368 56106 222380
rect 73062 222368 73068 222380
rect 73120 222368 73126 222420
rect 75362 222368 75368 222420
rect 75420 222408 75426 222420
rect 200942 222408 200948 222420
rect 75420 222380 200948 222408
rect 75420 222368 75426 222380
rect 200942 222368 200948 222380
rect 201000 222368 201006 222420
rect 205818 222368 205824 222420
rect 205876 222408 205882 222420
rect 257338 222408 257344 222420
rect 205876 222380 257344 222408
rect 205876 222368 205882 222380
rect 257338 222368 257344 222380
rect 257396 222368 257402 222420
rect 283190 222368 283196 222420
rect 283248 222408 283254 222420
rect 290090 222408 290096 222420
rect 283248 222380 290096 222408
rect 283248 222368 283254 222380
rect 290090 222368 290096 222380
rect 290148 222368 290154 222420
rect 314102 222368 314108 222420
rect 314160 222408 314166 222420
rect 334710 222408 334716 222420
rect 314160 222380 334716 222408
rect 314160 222368 314166 222380
rect 334710 222368 334716 222380
rect 334768 222368 334774 222420
rect 336458 222368 336464 222420
rect 336516 222408 336522 222420
rect 388530 222408 388536 222420
rect 336516 222380 388536 222408
rect 336516 222368 336522 222380
rect 388530 222368 388536 222380
rect 388588 222368 388594 222420
rect 408126 222368 408132 222420
rect 408184 222408 408190 222420
rect 561766 222408 561772 222420
rect 408184 222380 561772 222408
rect 408184 222368 408190 222380
rect 561766 222368 561772 222380
rect 561824 222368 561830 222420
rect 570230 222408 570236 222420
rect 569880 222380 570236 222408
rect 202414 222300 202420 222352
rect 202472 222340 202478 222352
rect 254210 222340 254216 222352
rect 202472 222312 254216 222340
rect 202472 222300 202478 222312
rect 254210 222300 254216 222312
rect 254268 222300 254274 222352
rect 311618 222300 311624 222352
rect 311676 222340 311682 222352
rect 333974 222340 333980 222352
rect 311676 222312 333980 222340
rect 311676 222300 311682 222312
rect 333974 222300 333980 222312
rect 334032 222300 334038 222352
rect 338850 222300 338856 222352
rect 338908 222340 338914 222352
rect 393590 222340 393596 222352
rect 338908 222312 393596 222340
rect 338908 222300 338914 222312
rect 393590 222300 393596 222312
rect 393648 222300 393654 222352
rect 408218 222300 408224 222352
rect 408276 222340 408282 222352
rect 555418 222340 555424 222352
rect 408276 222312 555424 222340
rect 408276 222300 408282 222312
rect 555418 222300 555424 222312
rect 555476 222300 555482 222352
rect 569880 222340 569908 222380
rect 570230 222368 570236 222380
rect 570288 222368 570294 222420
rect 555528 222312 569908 222340
rect 194042 222232 194048 222284
rect 194100 222272 194106 222284
rect 246942 222272 246948 222284
rect 194100 222244 246948 222272
rect 194100 222232 194106 222244
rect 246942 222232 246948 222244
rect 247000 222232 247006 222284
rect 314286 222232 314292 222284
rect 314344 222272 314350 222284
rect 338022 222272 338028 222284
rect 314344 222244 338028 222272
rect 314344 222232 314350 222244
rect 338022 222232 338028 222244
rect 338080 222232 338086 222284
rect 339218 222232 339224 222284
rect 339276 222272 339282 222284
rect 391934 222272 391940 222284
rect 339276 222244 391940 222272
rect 339276 222232 339282 222244
rect 391934 222232 391940 222244
rect 391992 222232 391998 222284
rect 413830 222232 413836 222284
rect 413888 222272 413894 222284
rect 555528 222272 555556 222312
rect 569954 222300 569960 222352
rect 570012 222340 570018 222352
rect 621014 222340 621020 222352
rect 570012 222312 621020 222340
rect 570012 222300 570018 222312
rect 621014 222300 621020 222312
rect 621072 222300 621078 222352
rect 565998 222272 566004 222284
rect 413888 222244 555556 222272
rect 555620 222244 566004 222272
rect 413888 222232 413894 222244
rect 54386 222164 54392 222216
rect 54444 222204 54450 222216
rect 193306 222204 193312 222216
rect 54444 222176 193312 222204
rect 54444 222164 54450 222176
rect 193306 222164 193312 222176
rect 193364 222164 193370 222216
rect 195698 222164 195704 222216
rect 195756 222204 195762 222216
rect 251450 222204 251456 222216
rect 195756 222176 251456 222204
rect 195756 222164 195762 222176
rect 251450 222164 251456 222176
rect 251508 222164 251514 222216
rect 317046 222164 317052 222216
rect 317104 222204 317110 222216
rect 345014 222204 345020 222216
rect 317104 222176 345020 222204
rect 317104 222164 317110 222176
rect 345014 222164 345020 222176
rect 345072 222164 345078 222216
rect 349062 222164 349068 222216
rect 349120 222204 349126 222216
rect 407022 222204 407028 222216
rect 349120 222176 407028 222204
rect 349120 222164 349126 222176
rect 407022 222164 407028 222176
rect 407080 222164 407086 222216
rect 409690 222164 409696 222216
rect 409748 222204 409754 222216
rect 555620 222204 555648 222244
rect 565998 222232 566004 222244
rect 566056 222272 566062 222284
rect 566056 222244 574094 222272
rect 566056 222232 566062 222244
rect 409748 222176 555648 222204
rect 409748 222164 409754 222176
rect 555694 222164 555700 222216
rect 555752 222204 555758 222216
rect 556154 222204 556160 222216
rect 555752 222176 556160 222204
rect 555752 222164 555758 222176
rect 556154 222164 556160 222176
rect 556212 222204 556218 222216
rect 574066 222204 574094 222244
rect 620554 222204 620560 222216
rect 556212 222176 570092 222204
rect 574066 222176 620560 222204
rect 556212 222164 556218 222176
rect 114922 222096 114928 222148
rect 114980 222136 114986 222148
rect 142154 222136 142160 222148
rect 114980 222108 142160 222136
rect 114980 222096 114986 222108
rect 142154 222096 142160 222108
rect 142212 222096 142218 222148
rect 148594 222096 148600 222148
rect 148652 222136 148658 222148
rect 232314 222136 232320 222148
rect 148652 222108 232320 222136
rect 148652 222096 148658 222108
rect 232314 222096 232320 222108
rect 232372 222096 232378 222148
rect 280614 222096 280620 222148
rect 280672 222136 280678 222148
rect 287238 222136 287244 222148
rect 280672 222108 287244 222136
rect 280672 222096 280678 222108
rect 287238 222096 287244 222108
rect 287296 222096 287302 222148
rect 322658 222096 322664 222148
rect 322716 222136 322722 222148
rect 360746 222136 360752 222148
rect 322716 222108 360752 222136
rect 322716 222096 322722 222108
rect 360746 222096 360752 222108
rect 360804 222096 360810 222148
rect 401410 222096 401416 222148
rect 401468 222136 401474 222148
rect 529014 222136 529020 222148
rect 401468 222108 529020 222136
rect 401468 222096 401474 222108
rect 529014 222096 529020 222108
rect 529072 222096 529078 222148
rect 536282 222096 536288 222148
rect 536340 222136 536346 222148
rect 548334 222136 548340 222148
rect 536340 222108 548340 222136
rect 536340 222096 536346 222108
rect 548334 222096 548340 222108
rect 548392 222096 548398 222148
rect 560754 222096 560760 222148
rect 560812 222136 560818 222148
rect 561582 222136 561588 222148
rect 560812 222108 561588 222136
rect 560812 222096 560818 222108
rect 561582 222096 561588 222108
rect 561640 222096 561646 222148
rect 569126 222096 569132 222148
rect 569184 222136 569190 222148
rect 569954 222136 569960 222148
rect 569184 222108 569960 222136
rect 569184 222096 569190 222108
rect 569954 222096 569960 222108
rect 570012 222096 570018 222148
rect 570064 222136 570092 222176
rect 620554 222164 620560 222176
rect 620612 222164 620618 222216
rect 652846 222164 652852 222216
rect 652904 222204 652910 222216
rect 652904 222176 670694 222204
rect 652904 222164 652910 222176
rect 633158 222136 633164 222148
rect 570064 222108 633164 222136
rect 633158 222096 633164 222108
rect 633216 222096 633222 222148
rect 670666 222136 670694 222176
rect 674558 222164 674564 222216
rect 674616 222204 674622 222216
rect 675754 222204 675760 222216
rect 674616 222176 675760 222204
rect 674616 222164 674622 222176
rect 675754 222164 675760 222176
rect 675812 222164 675818 222216
rect 674650 222136 674656 222148
rect 670666 222108 674656 222136
rect 674650 222096 674656 222108
rect 674708 222136 674714 222148
rect 675570 222136 675576 222148
rect 674708 222108 675576 222136
rect 674708 222096 674714 222108
rect 675570 222096 675576 222108
rect 675628 222096 675634 222148
rect 146938 222028 146944 222080
rect 146996 222068 147002 222080
rect 232590 222068 232596 222080
rect 146996 222040 232596 222068
rect 146996 222028 147002 222040
rect 232590 222028 232596 222040
rect 232648 222028 232654 222080
rect 233510 222028 233516 222080
rect 233568 222068 233574 222080
rect 248782 222068 248788 222080
rect 233568 222040 248788 222068
rect 233568 222028 233574 222040
rect 248782 222028 248788 222040
rect 248840 222028 248846 222080
rect 322566 222028 322572 222080
rect 322624 222068 322630 222080
rect 358262 222068 358268 222080
rect 322624 222040 358268 222068
rect 322624 222028 322630 222040
rect 358262 222028 358268 222040
rect 358320 222028 358326 222080
rect 389082 222028 389088 222080
rect 389140 222068 389146 222080
rect 513374 222068 513380 222080
rect 389140 222040 513380 222068
rect 389140 222028 389146 222040
rect 513374 222028 513380 222040
rect 513432 222028 513438 222080
rect 544930 222028 544936 222080
rect 544988 222068 544994 222080
rect 547506 222068 547512 222080
rect 544988 222040 547512 222068
rect 544988 222028 544994 222040
rect 547506 222028 547512 222040
rect 547564 222028 547570 222080
rect 552106 222028 552112 222080
rect 552164 222068 552170 222080
rect 552842 222068 552848 222080
rect 552164 222040 552848 222068
rect 552164 222028 552170 222040
rect 552842 222028 552848 222040
rect 552900 222068 552906 222080
rect 632698 222068 632704 222080
rect 552900 222040 632704 222068
rect 552900 222028 552906 222040
rect 632698 222028 632704 222040
rect 632756 222028 632762 222080
rect 153654 221960 153660 222012
rect 153712 222000 153718 222012
rect 235442 222000 235448 222012
rect 153712 221972 235448 222000
rect 153712 221960 153718 221972
rect 235442 221960 235448 221972
rect 235500 221960 235506 222012
rect 274726 221960 274732 222012
rect 274784 222000 274790 222012
rect 287606 222000 287612 222012
rect 274784 221972 287612 222000
rect 274784 221960 274790 221972
rect 287606 221960 287612 221972
rect 287664 221960 287670 222012
rect 322750 221960 322756 222012
rect 322808 222000 322814 222012
rect 356514 222000 356520 222012
rect 322808 221972 356520 222000
rect 322808 221960 322814 221972
rect 356514 221960 356520 221972
rect 356572 221960 356578 222012
rect 386322 221960 386328 222012
rect 386380 222000 386386 222012
rect 507946 222000 507952 222012
rect 386380 221972 507952 222000
rect 386380 221960 386386 221972
rect 507946 221960 507952 221972
rect 508004 221960 508010 222012
rect 533154 221960 533160 222012
rect 533212 222000 533218 222012
rect 533798 222000 533804 222012
rect 533212 221972 533804 222000
rect 533212 221960 533218 221972
rect 533798 221960 533804 221972
rect 533856 222000 533862 222012
rect 614574 222000 614580 222012
rect 533856 221972 614580 222000
rect 533856 221960 533862 221972
rect 614574 221960 614580 221972
rect 614632 221960 614638 222012
rect 93026 221892 93032 221944
rect 93084 221932 93090 221944
rect 153102 221932 153108 221944
rect 93084 221904 153108 221932
rect 93084 221892 93090 221904
rect 153102 221892 153108 221904
rect 153160 221892 153166 221944
rect 155310 221892 155316 221944
rect 155368 221932 155374 221944
rect 235166 221932 235172 221944
rect 155368 221904 235172 221932
rect 155368 221892 155374 221904
rect 235166 221892 235172 221904
rect 235224 221892 235230 221944
rect 319990 221892 319996 221944
rect 320048 221932 320054 221944
rect 354030 221932 354036 221944
rect 320048 221904 354036 221932
rect 320048 221892 320054 221904
rect 354030 221892 354036 221904
rect 354088 221892 354094 221944
rect 390554 221892 390560 221944
rect 390612 221932 390618 221944
rect 511350 221932 511356 221944
rect 390612 221904 511356 221932
rect 390612 221892 390618 221904
rect 511350 221892 511356 221904
rect 511408 221892 511414 221944
rect 530946 221892 530952 221944
rect 531004 221932 531010 221944
rect 614022 221932 614028 221944
rect 531004 221904 614028 221932
rect 531004 221892 531010 221904
rect 614022 221892 614028 221904
rect 614080 221892 614086 221944
rect 123386 221824 123392 221876
rect 123444 221864 123450 221876
rect 155954 221864 155960 221876
rect 123444 221836 155960 221864
rect 123444 221824 123450 221836
rect 155954 221824 155960 221836
rect 156012 221824 156018 221876
rect 160370 221824 160376 221876
rect 160428 221864 160434 221876
rect 160428 221836 232452 221864
rect 160428 221824 160434 221836
rect 125042 221756 125048 221808
rect 125100 221796 125106 221808
rect 156046 221796 156052 221808
rect 125100 221768 156052 221796
rect 125100 221756 125106 221768
rect 156046 221756 156052 221768
rect 156104 221756 156110 221808
rect 162026 221756 162032 221808
rect 162084 221796 162090 221808
rect 232222 221796 232228 221808
rect 162084 221768 232228 221796
rect 162084 221756 162090 221768
rect 232222 221756 232228 221768
rect 232280 221756 232286 221808
rect 99834 221688 99840 221740
rect 99892 221728 99898 221740
rect 161474 221728 161480 221740
rect 99892 221700 161480 221728
rect 99892 221688 99898 221700
rect 161474 221688 161480 221700
rect 161532 221688 161538 221740
rect 170490 221688 170496 221740
rect 170548 221728 170554 221740
rect 232424 221728 232452 221836
rect 234338 221824 234344 221876
rect 234396 221864 234402 221876
rect 249702 221864 249708 221876
rect 234396 221836 249708 221864
rect 234396 221824 234402 221836
rect 249702 221824 249708 221836
rect 249760 221824 249766 221876
rect 275554 221824 275560 221876
rect 275612 221864 275618 221876
rect 284846 221864 284852 221876
rect 275612 221836 284852 221864
rect 275612 221824 275618 221836
rect 284846 221824 284852 221836
rect 284904 221824 284910 221876
rect 322842 221824 322848 221876
rect 322900 221864 322906 221876
rect 357342 221864 357348 221876
rect 322900 221836 357348 221864
rect 322900 221824 322906 221836
rect 357342 221824 357348 221836
rect 357400 221824 357406 221876
rect 383562 221824 383568 221876
rect 383620 221864 383626 221876
rect 503530 221864 503536 221876
rect 383620 221836 503536 221864
rect 383620 221824 383626 221836
rect 503530 221824 503536 221836
rect 503588 221824 503594 221876
rect 541434 221824 541440 221876
rect 541492 221864 541498 221876
rect 542354 221864 542360 221876
rect 541492 221836 542360 221864
rect 541492 221824 541498 221836
rect 542354 221824 542360 221836
rect 542412 221824 542418 221876
rect 547506 221824 547512 221876
rect 547564 221864 547570 221876
rect 631778 221864 631784 221876
rect 547564 221836 631784 221864
rect 547564 221824 547570 221836
rect 631778 221824 631784 221836
rect 631836 221824 631842 221876
rect 232498 221756 232504 221808
rect 232556 221796 232562 221808
rect 237650 221796 237656 221808
rect 232556 221768 237656 221796
rect 232556 221756 232562 221768
rect 237650 221756 237656 221768
rect 237708 221756 237714 221808
rect 317138 221756 317144 221808
rect 317196 221796 317202 221808
rect 343910 221796 343916 221808
rect 317196 221768 343916 221796
rect 317196 221756 317202 221768
rect 343910 221756 343916 221768
rect 343968 221756 343974 221808
rect 346394 221756 346400 221808
rect 346452 221796 346458 221808
rect 380066 221796 380072 221808
rect 346452 221768 380072 221796
rect 346452 221756 346458 221768
rect 380066 221756 380072 221768
rect 380124 221756 380130 221808
rect 403066 221756 403072 221808
rect 403124 221796 403130 221808
rect 523954 221796 523960 221808
rect 403124 221768 523960 221796
rect 403124 221756 403130 221768
rect 523954 221756 523960 221768
rect 524012 221756 524018 221808
rect 528554 221756 528560 221808
rect 528612 221796 528618 221808
rect 613562 221796 613568 221808
rect 528612 221768 613568 221796
rect 528612 221756 528618 221768
rect 613562 221756 613568 221768
rect 613620 221756 613626 221808
rect 238294 221728 238300 221740
rect 170548 221700 232360 221728
rect 232424 221700 238300 221728
rect 170548 221688 170554 221700
rect 130102 221620 130108 221672
rect 130160 221660 130166 221672
rect 158622 221660 158628 221672
rect 130160 221632 158628 221660
rect 130160 221620 130166 221632
rect 158622 221620 158628 221632
rect 158680 221620 158686 221672
rect 168742 221620 168748 221672
rect 168800 221660 168806 221672
rect 232222 221660 232228 221672
rect 168800 221632 232228 221660
rect 168800 221620 168806 221632
rect 232222 221620 232228 221632
rect 232280 221620 232286 221672
rect 143442 221552 143448 221604
rect 143500 221592 143506 221604
rect 169662 221592 169668 221604
rect 143500 221564 169668 221592
rect 143500 221552 143506 221564
rect 169662 221552 169668 221564
rect 169720 221552 169726 221604
rect 175458 221552 175464 221604
rect 175516 221592 175522 221604
rect 232130 221592 232136 221604
rect 175516 221564 232136 221592
rect 175516 221552 175522 221564
rect 232130 221552 232136 221564
rect 232188 221552 232194 221604
rect 232332 221592 232360 221700
rect 238294 221688 238300 221700
rect 238352 221688 238358 221740
rect 322474 221688 322480 221740
rect 322532 221728 322538 221740
rect 354858 221728 354864 221740
rect 322532 221700 354864 221728
rect 322532 221688 322538 221700
rect 354858 221688 354864 221700
rect 354916 221688 354922 221740
rect 401318 221688 401324 221740
rect 401376 221728 401382 221740
rect 518894 221728 518900 221740
rect 401376 221700 518900 221728
rect 401376 221688 401382 221700
rect 518894 221688 518900 221700
rect 518952 221688 518958 221740
rect 545022 221688 545028 221740
rect 545080 221728 545086 221740
rect 631318 221728 631324 221740
rect 545080 221700 631324 221728
rect 545080 221688 545086 221700
rect 631318 221688 631324 221700
rect 631376 221688 631382 221740
rect 232406 221620 232412 221672
rect 232464 221660 232470 221672
rect 240502 221660 240508 221672
rect 232464 221632 240508 221660
rect 232464 221620 232470 221632
rect 240502 221620 240508 221632
rect 240560 221620 240566 221672
rect 279786 221620 279792 221672
rect 279844 221660 279850 221672
rect 287422 221660 287428 221672
rect 279844 221632 287428 221660
rect 279844 221620 279850 221632
rect 287422 221620 287428 221632
rect 287480 221620 287486 221672
rect 319806 221620 319812 221672
rect 319864 221660 319870 221672
rect 351454 221660 351460 221672
rect 319864 221632 351460 221660
rect 319864 221620 319870 221632
rect 351454 221620 351460 221632
rect 351512 221620 351518 221672
rect 387794 221620 387800 221672
rect 387852 221660 387858 221672
rect 506290 221660 506296 221672
rect 387852 221632 506296 221660
rect 387852 221620 387858 221632
rect 506290 221620 506296 221632
rect 506348 221620 506354 221672
rect 525886 221620 525892 221672
rect 525944 221660 525950 221672
rect 613102 221660 613108 221672
rect 525944 221632 613108 221660
rect 525944 221620 525950 221632
rect 613102 221620 613108 221632
rect 613160 221620 613166 221672
rect 241606 221592 241612 221604
rect 232332 221564 241612 221592
rect 241606 221552 241612 221564
rect 241664 221552 241670 221604
rect 276474 221552 276480 221604
rect 276532 221592 276538 221604
rect 287054 221592 287060 221604
rect 276532 221564 287060 221592
rect 276532 221552 276538 221564
rect 287054 221552 287060 221564
rect 287112 221552 287118 221604
rect 320082 221552 320088 221604
rect 320140 221592 320146 221604
rect 350626 221592 350632 221604
rect 320140 221564 350632 221592
rect 320140 221552 320146 221564
rect 350626 221552 350632 221564
rect 350684 221552 350690 221604
rect 380802 221552 380808 221604
rect 380860 221592 380866 221604
rect 497366 221592 497372 221604
rect 380860 221564 497372 221592
rect 380860 221552 380866 221564
rect 497366 221552 497372 221564
rect 497424 221592 497430 221604
rect 499482 221592 499488 221604
rect 497424 221564 499488 221592
rect 497424 221552 497430 221564
rect 499482 221552 499488 221564
rect 499540 221552 499546 221604
rect 516106 221564 531820 221592
rect 136818 221484 136824 221536
rect 136876 221524 136882 221536
rect 161566 221524 161572 221536
rect 136876 221496 161572 221524
rect 136876 221484 136882 221496
rect 161566 221484 161572 221496
rect 161624 221484 161630 221536
rect 177206 221484 177212 221536
rect 177264 221524 177270 221536
rect 229278 221524 229284 221536
rect 177264 221496 229284 221524
rect 177264 221484 177270 221496
rect 229278 221484 229284 221496
rect 229336 221484 229342 221536
rect 229554 221484 229560 221536
rect 229612 221524 229618 221536
rect 235994 221524 236000 221536
rect 229612 221496 236000 221524
rect 229612 221484 229618 221496
rect 235994 221484 236000 221496
rect 236052 221484 236058 221536
rect 236914 221484 236920 221536
rect 236972 221524 236978 221536
rect 241514 221524 241520 221536
rect 236972 221496 241520 221524
rect 236972 221484 236978 221496
rect 241514 221484 241520 221496
rect 241572 221484 241578 221536
rect 246114 221484 246120 221536
rect 246172 221524 246178 221536
rect 257982 221524 257988 221536
rect 246172 221496 257988 221524
rect 246172 221484 246178 221496
rect 257982 221484 257988 221496
rect 258040 221484 258046 221536
rect 314378 221484 314384 221536
rect 314436 221524 314442 221536
rect 340598 221524 340604 221536
rect 314436 221496 340604 221524
rect 314436 221484 314442 221496
rect 340598 221484 340604 221496
rect 340656 221484 340662 221536
rect 343726 221484 343732 221536
rect 343784 221524 343790 221536
rect 373350 221524 373356 221536
rect 343784 221496 373356 221524
rect 343784 221484 343790 221496
rect 373350 221484 373356 221496
rect 373408 221484 373414 221536
rect 384942 221484 384948 221536
rect 385000 221524 385006 221536
rect 501230 221524 501236 221536
rect 385000 221496 501236 221524
rect 385000 221484 385006 221496
rect 501230 221484 501236 221496
rect 501288 221484 501294 221536
rect 182082 221416 182088 221468
rect 182140 221456 182146 221468
rect 246022 221456 246028 221468
rect 182140 221428 229324 221456
rect 182140 221416 182146 221428
rect 57698 221348 57704 221400
rect 57756 221388 57762 221400
rect 62022 221388 62028 221400
rect 57756 221360 62028 221388
rect 57756 221348 57762 221360
rect 62022 221348 62028 221360
rect 62080 221348 62086 221400
rect 76282 221348 76288 221400
rect 76340 221388 76346 221400
rect 78582 221388 78588 221400
rect 76340 221360 78588 221388
rect 76340 221348 76346 221360
rect 78582 221348 78588 221360
rect 78640 221348 78646 221400
rect 138474 221348 138480 221400
rect 138532 221388 138538 221400
rect 147582 221388 147588 221400
rect 138532 221360 147588 221388
rect 138532 221348 138538 221360
rect 147582 221348 147588 221360
rect 147640 221348 147646 221400
rect 150342 221388 150348 221400
rect 149026 221360 150348 221388
rect 52730 221280 52736 221332
rect 52788 221320 52794 221332
rect 67542 221320 67548 221332
rect 52788 221292 67548 221320
rect 52788 221280 52794 221292
rect 67542 221280 67548 221292
rect 67600 221280 67606 221332
rect 77938 221280 77944 221332
rect 77996 221320 78002 221332
rect 86862 221320 86868 221332
rect 77996 221292 86868 221320
rect 77996 221280 78002 221292
rect 86862 221280 86868 221292
rect 86920 221280 86926 221332
rect 131758 221280 131764 221332
rect 131816 221320 131822 221332
rect 142062 221320 142068 221332
rect 131816 221292 142068 221320
rect 131816 221280 131822 221292
rect 142062 221280 142068 221292
rect 142120 221280 142126 221332
rect 145190 221280 145196 221332
rect 145248 221320 145254 221332
rect 149026 221320 149054 221360
rect 150342 221348 150348 221360
rect 150400 221348 150406 221400
rect 151722 221348 151728 221400
rect 151780 221388 151786 221400
rect 155862 221388 155868 221400
rect 151780 221360 155868 221388
rect 151780 221348 151786 221360
rect 155862 221348 155868 221360
rect 155920 221348 155926 221400
rect 158714 221348 158720 221400
rect 158772 221388 158778 221400
rect 159818 221388 159824 221400
rect 158772 221360 159824 221388
rect 158772 221348 158778 221360
rect 159818 221348 159824 221360
rect 159876 221348 159882 221400
rect 163682 221348 163688 221400
rect 163740 221388 163746 221400
rect 165338 221388 165344 221400
rect 163740 221360 165344 221388
rect 163740 221348 163746 221360
rect 165338 221348 165344 221360
rect 165396 221348 165402 221400
rect 172146 221348 172152 221400
rect 172204 221388 172210 221400
rect 173802 221388 173808 221400
rect 172204 221360 173808 221388
rect 172204 221348 172210 221360
rect 173802 221348 173808 221360
rect 173860 221348 173866 221400
rect 183922 221348 183928 221400
rect 183980 221388 183986 221400
rect 227530 221388 227536 221400
rect 183980 221360 227536 221388
rect 183980 221348 183986 221360
rect 227530 221348 227536 221360
rect 227588 221348 227594 221400
rect 227622 221348 227628 221400
rect 227680 221388 227686 221400
rect 229002 221388 229008 221400
rect 227680 221360 229008 221388
rect 227680 221348 227686 221360
rect 229002 221348 229008 221360
rect 229060 221348 229066 221400
rect 229296 221388 229324 221428
rect 229480 221428 246028 221456
rect 229480 221388 229508 221428
rect 246022 221416 246028 221428
rect 246080 221416 246086 221468
rect 249518 221416 249524 221468
rect 249576 221456 249582 221468
rect 258166 221456 258172 221468
rect 249576 221428 258172 221456
rect 249576 221416 249582 221428
rect 258166 221416 258172 221428
rect 258224 221416 258230 221468
rect 271414 221416 271420 221468
rect 271472 221456 271478 221468
rect 284662 221456 284668 221468
rect 271472 221428 284668 221456
rect 271472 221416 271478 221428
rect 284662 221416 284668 221428
rect 284720 221416 284726 221468
rect 317322 221416 317328 221468
rect 317380 221456 317386 221468
rect 317380 221428 319668 221456
rect 317380 221416 317386 221428
rect 229296 221360 229508 221388
rect 232130 221348 232136 221400
rect 232188 221388 232194 221400
rect 232188 221360 233648 221388
rect 232188 221348 232194 221360
rect 145248 221292 149054 221320
rect 145248 221280 145254 221292
rect 150250 221280 150256 221332
rect 150308 221320 150314 221332
rect 153194 221320 153200 221332
rect 150308 221292 153200 221320
rect 150308 221280 150314 221292
rect 153194 221280 153200 221292
rect 153252 221280 153258 221332
rect 156966 221280 156972 221332
rect 157024 221320 157030 221332
rect 161382 221320 161388 221332
rect 157024 221292 161388 221320
rect 157024 221280 157030 221292
rect 161382 221280 161388 221292
rect 161440 221280 161446 221332
rect 167086 221280 167092 221332
rect 167144 221320 167150 221332
rect 168098 221320 168104 221332
rect 167144 221292 168104 221320
rect 167144 221280 167150 221292
rect 168098 221280 168104 221292
rect 168156 221280 168162 221332
rect 178862 221280 178868 221332
rect 178920 221320 178926 221332
rect 179322 221320 179328 221332
rect 178920 221292 179328 221320
rect 178920 221280 178926 221292
rect 179322 221280 179328 221292
rect 179380 221280 179386 221332
rect 185578 221280 185584 221332
rect 185636 221320 185642 221332
rect 187602 221320 187608 221332
rect 185636 221292 187608 221320
rect 185636 221280 185642 221292
rect 187602 221280 187608 221292
rect 187660 221280 187666 221332
rect 192294 221280 192300 221332
rect 192352 221320 192358 221332
rect 192938 221320 192944 221332
rect 192352 221292 192944 221320
rect 192352 221280 192358 221292
rect 192938 221280 192944 221292
rect 192996 221280 193002 221332
rect 196526 221280 196532 221332
rect 196584 221320 196590 221332
rect 200850 221320 200856 221332
rect 196584 221292 200856 221320
rect 196584 221280 196590 221292
rect 200850 221280 200856 221292
rect 200908 221280 200914 221332
rect 208026 221280 208032 221332
rect 208084 221320 208090 221332
rect 233510 221320 233516 221332
rect 208084 221292 233516 221320
rect 208084 221280 208090 221292
rect 233510 221280 233516 221292
rect 233568 221280 233574 221332
rect 233620 221320 233648 221360
rect 235258 221348 235264 221400
rect 235316 221388 235322 221400
rect 237282 221388 237288 221400
rect 235316 221360 237288 221388
rect 235316 221348 235322 221360
rect 237282 221348 237288 221360
rect 237340 221348 237346 221400
rect 243262 221388 243268 221400
rect 237392 221360 243268 221388
rect 237392 221320 237420 221360
rect 243262 221348 243268 221360
rect 243320 221348 243326 221400
rect 247034 221348 247040 221400
rect 247092 221388 247098 221400
rect 248322 221388 248328 221400
rect 247092 221360 248328 221388
rect 247092 221348 247098 221360
rect 248322 221348 248328 221360
rect 248380 221348 248386 221400
rect 254578 221348 254584 221400
rect 254636 221388 254642 221400
rect 256510 221388 256516 221400
rect 254636 221360 256516 221388
rect 254636 221348 254642 221360
rect 256510 221348 256516 221360
rect 256568 221348 256574 221400
rect 257062 221348 257068 221400
rect 257120 221388 257126 221400
rect 259178 221388 259184 221400
rect 257120 221360 259184 221388
rect 257120 221348 257126 221360
rect 259178 221348 259184 221360
rect 259236 221348 259242 221400
rect 289722 221348 289728 221400
rect 289780 221388 289786 221400
rect 292942 221388 292948 221400
rect 289780 221360 292948 221388
rect 289780 221348 289786 221360
rect 292942 221348 292948 221360
rect 293000 221348 293006 221400
rect 298094 221348 298100 221400
rect 298152 221388 298158 221400
rect 299382 221388 299388 221400
rect 298152 221360 299388 221388
rect 298152 221348 298158 221360
rect 299382 221348 299388 221360
rect 299440 221348 299446 221400
rect 300946 221348 300952 221400
rect 301004 221388 301010 221400
rect 302694 221388 302700 221400
rect 301004 221360 302700 221388
rect 301004 221348 301010 221360
rect 302694 221348 302700 221360
rect 302752 221348 302758 221400
rect 309778 221348 309784 221400
rect 309836 221388 309842 221400
rect 311158 221388 311164 221400
rect 309836 221360 311164 221388
rect 309836 221348 309842 221360
rect 311158 221348 311164 221360
rect 311216 221348 311222 221400
rect 315022 221348 315028 221400
rect 315080 221388 315086 221400
rect 315482 221388 315488 221400
rect 315080 221360 315488 221388
rect 315080 221348 315086 221360
rect 315482 221348 315488 221360
rect 315540 221348 315546 221400
rect 317782 221348 317788 221400
rect 317840 221388 317846 221400
rect 319530 221388 319536 221400
rect 317840 221360 319536 221388
rect 317840 221348 317846 221360
rect 319530 221348 319536 221360
rect 319588 221348 319594 221400
rect 319640 221388 319668 221428
rect 319898 221416 319904 221468
rect 319956 221456 319962 221468
rect 348142 221456 348148 221468
rect 319956 221428 348148 221456
rect 319956 221416 319962 221428
rect 348142 221416 348148 221428
rect 348200 221416 348206 221468
rect 379422 221416 379428 221468
rect 379480 221456 379486 221468
rect 484394 221456 484400 221468
rect 379480 221428 484400 221456
rect 379480 221416 379486 221428
rect 484394 221416 484400 221428
rect 484452 221416 484458 221468
rect 513374 221416 513380 221468
rect 513432 221456 513438 221468
rect 516106 221456 516134 221564
rect 513432 221428 516134 221456
rect 513432 221416 513438 221428
rect 343082 221388 343088 221400
rect 319640 221360 343088 221388
rect 343082 221348 343088 221360
rect 343140 221348 343146 221400
rect 343634 221348 343640 221400
rect 343692 221388 343698 221400
rect 366634 221388 366640 221400
rect 343692 221360 366640 221388
rect 343692 221348 343698 221360
rect 366634 221348 366640 221360
rect 366692 221348 366698 221400
rect 387610 221348 387616 221400
rect 387668 221388 387674 221400
rect 491294 221388 491300 221400
rect 387668 221360 491300 221388
rect 387668 221348 387674 221360
rect 491294 221348 491300 221360
rect 491352 221348 491358 221400
rect 507946 221348 507952 221400
rect 508004 221388 508010 221400
rect 531792 221388 531820 221564
rect 536742 221552 536748 221604
rect 536800 221592 536806 221604
rect 538030 221592 538036 221604
rect 536800 221564 538036 221592
rect 536800 221552 536806 221564
rect 538030 221552 538036 221564
rect 538088 221592 538094 221604
rect 538088 221564 554360 221592
rect 538088 221552 538094 221564
rect 539502 221484 539508 221536
rect 539560 221524 539566 221536
rect 541618 221524 541624 221536
rect 539560 221496 541624 221524
rect 539560 221484 539566 221496
rect 541618 221484 541624 221496
rect 541676 221484 541682 221536
rect 542262 221484 542268 221536
rect 542320 221524 542326 221536
rect 544102 221524 544108 221536
rect 542320 221496 544108 221524
rect 542320 221484 542326 221496
rect 544102 221484 544108 221496
rect 544160 221484 544166 221536
rect 547782 221484 547788 221536
rect 547840 221524 547846 221536
rect 549254 221524 549260 221536
rect 547840 221496 549260 221524
rect 547840 221484 547846 221496
rect 549254 221484 549260 221496
rect 549312 221484 549318 221536
rect 552290 221484 552296 221536
rect 552348 221524 552354 221536
rect 554222 221524 554228 221536
rect 552348 221496 554228 221524
rect 552348 221484 552354 221496
rect 554222 221484 554228 221496
rect 554280 221484 554286 221536
rect 554332 221524 554360 221564
rect 554406 221552 554412 221604
rect 554464 221592 554470 221604
rect 630858 221592 630864 221604
rect 554464 221564 630864 221592
rect 554464 221552 554470 221564
rect 630858 221552 630864 221564
rect 630916 221552 630922 221604
rect 629938 221524 629944 221536
rect 554332 221496 629944 221524
rect 629938 221484 629944 221496
rect 629996 221484 630002 221536
rect 532970 221416 532976 221468
rect 533028 221456 533034 221468
rect 533982 221456 533988 221468
rect 533028 221428 533988 221456
rect 533028 221416 533034 221428
rect 533982 221416 533988 221428
rect 534040 221456 534046 221468
rect 628926 221456 628932 221468
rect 534040 221428 628932 221456
rect 534040 221416 534046 221428
rect 628926 221416 628932 221428
rect 628984 221416 628990 221468
rect 610802 221388 610808 221400
rect 508004 221360 531636 221388
rect 531792 221360 610808 221388
rect 508004 221348 508010 221360
rect 233620 221292 237420 221320
rect 239398 221280 239404 221332
rect 239456 221320 239462 221332
rect 240042 221320 240048 221332
rect 239456 221292 240048 221320
rect 239456 221280 239462 221292
rect 240042 221280 240048 221292
rect 240100 221280 240106 221332
rect 241974 221280 241980 221332
rect 242032 221320 242038 221332
rect 242802 221320 242808 221332
rect 242032 221292 242808 221320
rect 242032 221280 242038 221292
rect 242802 221280 242808 221292
rect 242860 221280 242866 221332
rect 250346 221280 250352 221332
rect 250404 221320 250410 221332
rect 250990 221320 250996 221332
rect 250404 221292 250996 221320
rect 250404 221280 250410 221292
rect 250990 221280 250996 221292
rect 251048 221280 251054 221332
rect 252922 221280 252928 221332
rect 252980 221320 252986 221332
rect 258074 221320 258080 221332
rect 252980 221292 258080 221320
rect 252980 221280 252986 221292
rect 258074 221280 258080 221292
rect 258132 221280 258138 221332
rect 258810 221280 258816 221332
rect 258868 221320 258874 221332
rect 259362 221320 259368 221332
rect 258868 221292 259368 221320
rect 258868 221280 258874 221292
rect 259362 221280 259368 221292
rect 259420 221280 259426 221332
rect 268838 221280 268844 221332
rect 268896 221320 268902 221332
rect 281718 221320 281724 221332
rect 268896 221292 281724 221320
rect 268896 221280 268902 221292
rect 281718 221280 281724 221292
rect 281776 221280 281782 221332
rect 286502 221280 286508 221332
rect 286560 221320 286566 221332
rect 290366 221320 290372 221332
rect 286560 221292 290372 221320
rect 286560 221280 286566 221292
rect 290366 221280 290372 221292
rect 290424 221280 290430 221332
rect 292390 221280 292396 221332
rect 292448 221320 292454 221332
rect 293218 221320 293224 221332
rect 292448 221292 293224 221320
rect 292448 221280 292454 221292
rect 293218 221280 293224 221292
rect 293276 221280 293282 221332
rect 295794 221280 295800 221332
rect 295852 221320 295858 221332
rect 297634 221320 297640 221332
rect 295852 221292 297640 221320
rect 295852 221280 295858 221292
rect 297634 221280 297640 221292
rect 297692 221280 297698 221332
rect 298278 221280 298284 221332
rect 298336 221320 298342 221332
rect 300210 221320 300216 221332
rect 298336 221292 300216 221320
rect 298336 221280 298342 221292
rect 300210 221280 300216 221292
rect 300268 221280 300274 221332
rect 300854 221280 300860 221332
rect 300912 221320 300918 221332
rect 301866 221320 301872 221332
rect 300912 221292 301872 221320
rect 300912 221280 300918 221292
rect 301866 221280 301872 221292
rect 301924 221280 301930 221332
rect 303706 221280 303712 221332
rect 303764 221320 303770 221332
rect 305270 221320 305276 221332
rect 303764 221292 305276 221320
rect 303764 221280 303770 221292
rect 305270 221280 305276 221292
rect 305328 221280 305334 221332
rect 306742 221280 306748 221332
rect 306800 221320 306806 221332
rect 308582 221320 308588 221332
rect 306800 221292 308588 221320
rect 306800 221280 306806 221292
rect 308582 221280 308588 221292
rect 308640 221280 308646 221332
rect 309410 221280 309416 221332
rect 309468 221320 309474 221332
rect 310238 221320 310244 221332
rect 309468 221292 310244 221320
rect 309468 221280 309474 221292
rect 310238 221280 310244 221292
rect 310296 221280 310302 221332
rect 315298 221280 315304 221332
rect 315356 221320 315362 221332
rect 316126 221320 316132 221332
rect 315356 221292 316132 221320
rect 315356 221280 315362 221292
rect 316126 221280 316132 221292
rect 316184 221280 316190 221332
rect 317598 221280 317604 221332
rect 317656 221320 317662 221332
rect 317966 221320 317972 221332
rect 317656 221292 317972 221320
rect 317656 221280 317662 221292
rect 317966 221280 317972 221292
rect 318024 221280 318030 221332
rect 318076 221292 337056 221320
rect 84654 221212 84660 221264
rect 84712 221252 84718 221264
rect 95142 221252 95148 221264
rect 84712 221224 95148 221252
rect 84712 221212 84718 221224
rect 95142 221212 95148 221224
rect 95200 221212 95206 221264
rect 187234 221212 187240 221264
rect 187292 221252 187298 221264
rect 226610 221252 226616 221264
rect 187292 221224 226616 221252
rect 187292 221212 187298 221224
rect 226610 221212 226616 221224
rect 226668 221212 226674 221264
rect 226702 221212 226708 221264
rect 226760 221252 226766 221264
rect 233234 221252 233240 221264
rect 226760 221224 233240 221252
rect 226760 221212 226766 221224
rect 233234 221212 233240 221224
rect 233292 221212 233298 221264
rect 238570 221212 238576 221264
rect 238628 221252 238634 221264
rect 239950 221252 239956 221264
rect 238628 221224 239956 221252
rect 238628 221212 238634 221224
rect 239950 221212 239956 221224
rect 240008 221212 240014 221264
rect 247862 221212 247868 221264
rect 247920 221252 247926 221264
rect 255222 221252 255228 221264
rect 247920 221224 255228 221252
rect 247920 221212 247926 221224
rect 255222 221212 255228 221224
rect 255280 221212 255286 221264
rect 256234 221212 256240 221264
rect 256292 221252 256298 221264
rect 260834 221252 260840 221264
rect 256292 221224 260840 221252
rect 256292 221212 256298 221224
rect 260834 221212 260840 221224
rect 260892 221212 260898 221264
rect 285674 221212 285680 221264
rect 285732 221252 285738 221264
rect 290458 221252 290464 221264
rect 285732 221224 290464 221252
rect 285732 221212 285738 221224
rect 290458 221212 290464 221224
rect 290516 221212 290522 221264
rect 316954 221212 316960 221264
rect 317012 221252 317018 221264
rect 318076 221252 318104 221292
rect 317012 221224 318104 221252
rect 318168 221224 336964 221252
rect 317012 221212 317018 221224
rect 59170 221144 59176 221196
rect 59228 221184 59234 221196
rect 193674 221184 193680 221196
rect 59228 221156 193680 221184
rect 59228 221144 59234 221156
rect 193674 221144 193680 221156
rect 193732 221144 193738 221196
rect 200758 221144 200764 221196
rect 200816 221184 200822 221196
rect 246942 221184 246948 221196
rect 200816 221156 246948 221184
rect 200816 221144 200822 221156
rect 246942 221144 246948 221156
rect 247000 221144 247006 221196
rect 252002 221144 252008 221196
rect 252060 221184 252066 221196
rect 253750 221184 253756 221196
rect 252060 221156 253756 221184
rect 252060 221144 252066 221156
rect 253750 221144 253756 221156
rect 253808 221144 253814 221196
rect 259362 221144 259368 221196
rect 259420 221184 259426 221196
rect 260742 221184 260748 221196
rect 259420 221156 260748 221184
rect 259420 221144 259426 221156
rect 260742 221144 260748 221156
rect 260800 221144 260806 221196
rect 263778 221144 263784 221196
rect 263836 221184 263842 221196
rect 264698 221184 264704 221196
rect 263836 221156 264704 221184
rect 263836 221144 263842 221156
rect 264698 221144 264704 221156
rect 264756 221144 264762 221196
rect 269666 221144 269672 221196
rect 269724 221184 269730 221196
rect 270402 221184 270408 221196
rect 269724 221156 270408 221184
rect 269724 221144 269730 221156
rect 270402 221144 270408 221156
rect 270460 221144 270466 221196
rect 283926 221144 283932 221196
rect 283984 221184 283990 221196
rect 287882 221184 287888 221196
rect 283984 221156 287888 221184
rect 283984 221144 283990 221156
rect 287882 221144 287888 221156
rect 287940 221144 287946 221196
rect 288250 221144 288256 221196
rect 288308 221184 288314 221196
rect 292850 221184 292856 221196
rect 288308 221156 292856 221184
rect 288308 221144 288314 221156
rect 292850 221144 292856 221156
rect 292908 221144 292914 221196
rect 314470 221144 314476 221196
rect 314528 221184 314534 221196
rect 318168 221184 318196 221224
rect 336734 221184 336740 221196
rect 314528 221156 318196 221184
rect 318260 221156 336740 221184
rect 314528 221144 314534 221156
rect 196342 221116 196348 221128
rect 168346 221088 196348 221116
rect 68646 221008 68652 221060
rect 68704 221048 68710 221060
rect 168346 221048 168374 221088
rect 196342 221076 196348 221088
rect 196400 221076 196406 221128
rect 199930 221076 199936 221128
rect 199988 221116 199994 221128
rect 208118 221116 208124 221128
rect 199988 221088 208124 221116
rect 199988 221076 199994 221088
rect 208118 221076 208124 221088
rect 208176 221076 208182 221128
rect 226702 221116 226708 221128
rect 208228 221088 226708 221116
rect 68704 221020 168374 221048
rect 68704 221008 68710 221020
rect 180518 221008 180524 221060
rect 180576 221048 180582 221060
rect 183462 221048 183468 221060
rect 180576 221020 183468 221048
rect 180576 221008 180582 221020
rect 183462 221008 183468 221020
rect 183520 221008 183526 221060
rect 188982 221008 188988 221060
rect 189040 221048 189046 221060
rect 208026 221048 208032 221060
rect 189040 221020 208032 221048
rect 189040 221008 189046 221020
rect 208026 221008 208032 221020
rect 208084 221008 208090 221060
rect 64506 220940 64512 220992
rect 64564 220980 64570 220992
rect 75822 220980 75828 220992
rect 64564 220952 75828 220980
rect 64564 220940 64570 220952
rect 75822 220940 75828 220952
rect 75880 220940 75886 220992
rect 197354 220940 197360 220992
rect 197412 220980 197418 220992
rect 198642 220980 198648 220992
rect 197412 220952 198648 220980
rect 197412 220940 197418 220952
rect 198642 220940 198648 220952
rect 198700 220940 198706 220992
rect 206646 220940 206652 220992
rect 206704 220980 206710 220992
rect 208118 220980 208124 220992
rect 206704 220952 208124 220980
rect 206704 220940 206710 220952
rect 208118 220940 208124 220952
rect 208176 220940 208182 220992
rect 69474 220872 69480 220924
rect 69532 220912 69538 220924
rect 73154 220912 73160 220924
rect 69532 220884 73160 220912
rect 69532 220872 69538 220884
rect 73154 220872 73160 220884
rect 73212 220872 73218 220924
rect 91370 220872 91376 220924
rect 91428 220912 91434 220924
rect 189718 220912 189724 220924
rect 91428 220884 189724 220912
rect 91428 220872 91434 220884
rect 189718 220872 189724 220884
rect 189776 220872 189782 220924
rect 189810 220872 189816 220924
rect 189868 220912 189874 220924
rect 208228 220912 208256 221088
rect 226702 221076 226708 221088
rect 226760 221076 226766 221128
rect 226794 221076 226800 221128
rect 226852 221116 226858 221128
rect 238754 221116 238760 221128
rect 226852 221088 238760 221116
rect 226852 221076 226858 221088
rect 238754 221076 238760 221088
rect 238812 221076 238818 221128
rect 240042 221076 240048 221128
rect 240100 221116 240106 221128
rect 241422 221116 241428 221128
rect 240100 221088 241428 221116
rect 240100 221076 240106 221088
rect 241422 221076 241428 221088
rect 241480 221076 241486 221128
rect 250990 221076 250996 221128
rect 251048 221116 251054 221128
rect 255406 221116 255412 221128
rect 251048 221088 255412 221116
rect 251048 221076 251054 221088
rect 255406 221076 255412 221088
rect 255464 221076 255470 221128
rect 277302 221076 277308 221128
rect 277360 221116 277366 221128
rect 284478 221116 284484 221128
rect 277360 221088 284484 221116
rect 277360 221076 277366 221088
rect 284478 221076 284484 221088
rect 284536 221076 284542 221128
rect 287330 221076 287336 221128
rect 287388 221116 287394 221128
rect 289998 221116 290004 221128
rect 287388 221088 290004 221116
rect 287388 221076 287394 221088
rect 289998 221076 290004 221088
rect 290056 221076 290062 221128
rect 314562 221076 314568 221128
rect 314620 221116 314626 221128
rect 318260 221116 318288 221156
rect 336734 221144 336740 221156
rect 336792 221144 336798 221196
rect 314620 221088 318288 221116
rect 336936 221116 336964 221224
rect 337028 221184 337056 221292
rect 337102 221280 337108 221332
rect 337160 221320 337166 221332
rect 338850 221320 338856 221332
rect 337160 221292 338856 221320
rect 337160 221280 337166 221292
rect 338850 221280 338856 221292
rect 338908 221280 338914 221332
rect 340782 221280 340788 221332
rect 340840 221320 340846 221332
rect 340840 221292 342254 221320
rect 340840 221280 340846 221292
rect 340874 221212 340880 221264
rect 340932 221252 340938 221264
rect 342226 221252 342254 221292
rect 351086 221280 351092 221332
rect 351144 221320 351150 221332
rect 352374 221320 352380 221332
rect 351144 221292 352380 221320
rect 351144 221280 351150 221292
rect 352374 221280 352380 221292
rect 352432 221280 352438 221332
rect 390370 221280 390376 221332
rect 390428 221320 390434 221332
rect 494514 221320 494520 221332
rect 390428 221292 494520 221320
rect 390428 221280 390434 221292
rect 494514 221280 494520 221292
rect 494572 221280 494578 221332
rect 511902 221280 511908 221332
rect 511960 221320 511966 221332
rect 516410 221320 516416 221332
rect 511960 221292 516416 221320
rect 511960 221280 511966 221292
rect 516410 221280 516416 221292
rect 516468 221280 516474 221332
rect 520182 221280 520188 221332
rect 520240 221320 520246 221332
rect 521654 221320 521660 221332
rect 520240 221292 521660 221320
rect 520240 221280 520246 221292
rect 521654 221280 521660 221292
rect 521712 221280 521718 221332
rect 524414 221280 524420 221332
rect 524472 221320 524478 221332
rect 526438 221320 526444 221332
rect 524472 221292 526444 221320
rect 524472 221280 524478 221292
rect 526438 221280 526444 221292
rect 526496 221280 526502 221332
rect 529934 221280 529940 221332
rect 529992 221320 529998 221332
rect 531498 221320 531504 221332
rect 529992 221292 531504 221320
rect 529992 221280 529998 221292
rect 531498 221280 531504 221292
rect 531556 221280 531562 221332
rect 531608 221320 531636 221360
rect 610802 221348 610808 221360
rect 610860 221348 610866 221400
rect 609882 221320 609888 221332
rect 531608 221292 609888 221320
rect 609882 221280 609888 221292
rect 609940 221280 609946 221332
rect 359918 221252 359924 221264
rect 340932 221224 341564 221252
rect 342226 221224 359924 221252
rect 340932 221212 340938 221224
rect 341426 221184 341432 221196
rect 337028 221156 341432 221184
rect 341426 221144 341432 221156
rect 341484 221144 341490 221196
rect 341536 221184 341564 221224
rect 359918 221212 359924 221224
rect 359976 221212 359982 221264
rect 413922 221212 413928 221264
rect 413980 221252 413986 221264
rect 413980 221224 477494 221252
rect 413980 221212 413986 221224
rect 353294 221184 353300 221196
rect 341536 221156 353300 221184
rect 353294 221144 353300 221156
rect 353352 221144 353358 221196
rect 477466 221184 477494 221224
rect 481542 221212 481548 221264
rect 481600 221252 481606 221264
rect 487798 221252 487804 221264
rect 481600 221224 487804 221252
rect 481600 221212 481606 221224
rect 487798 221212 487804 221224
rect 487856 221212 487862 221264
rect 489822 221212 489828 221264
rect 489880 221252 489886 221264
rect 497826 221252 497832 221264
rect 489880 221224 497832 221252
rect 489880 221212 489886 221224
rect 497826 221212 497832 221224
rect 497884 221212 497890 221264
rect 511074 221212 511080 221264
rect 511132 221252 511138 221264
rect 511994 221252 512000 221264
rect 511132 221224 512000 221252
rect 511132 221212 511138 221224
rect 511994 221212 512000 221224
rect 512052 221252 512058 221264
rect 610342 221252 610348 221264
rect 512052 221224 610348 221252
rect 512052 221212 512058 221224
rect 610342 221212 610348 221224
rect 610400 221212 610406 221264
rect 485222 221184 485228 221196
rect 477466 221156 485228 221184
rect 485222 221144 485228 221156
rect 485280 221144 485286 221196
rect 506106 221144 506112 221196
rect 506164 221184 506170 221196
rect 609422 221184 609428 221196
rect 506164 221156 609428 221184
rect 506164 221144 506170 221156
rect 609422 221144 609428 221156
rect 609480 221144 609486 221196
rect 669682 221144 669688 221196
rect 669740 221184 669746 221196
rect 676030 221184 676036 221196
rect 669740 221156 676036 221184
rect 669740 221144 669746 221156
rect 676030 221144 676036 221156
rect 676088 221144 676094 221196
rect 337194 221116 337200 221128
rect 336936 221088 337200 221116
rect 314620 221076 314626 221088
rect 337194 221076 337200 221088
rect 337252 221076 337258 221128
rect 338114 221076 338120 221128
rect 338172 221116 338178 221128
rect 349798 221116 349804 221128
rect 338172 221088 349804 221116
rect 338172 221076 338178 221088
rect 349798 221076 349804 221088
rect 349856 221076 349862 221128
rect 503530 221076 503536 221128
rect 503588 221116 503594 221128
rect 608962 221116 608968 221128
rect 503588 221088 608968 221116
rect 503588 221076 503594 221088
rect 608962 221076 608968 221088
rect 609020 221076 609026 221128
rect 208394 221008 208400 221060
rect 208452 221048 208458 221060
rect 208452 221020 229784 221048
rect 208452 221008 208458 221020
rect 229756 220980 229784 221020
rect 230198 221008 230204 221060
rect 230256 221048 230262 221060
rect 238938 221048 238944 221060
rect 230256 221020 238944 221048
rect 230256 221008 230262 221020
rect 238938 221008 238944 221020
rect 238996 221008 239002 221060
rect 260466 221008 260472 221060
rect 260524 221048 260530 221060
rect 261938 221048 261944 221060
rect 260524 221020 261944 221048
rect 260524 221008 260530 221020
rect 261938 221008 261944 221020
rect 261996 221008 262002 221060
rect 270402 221008 270408 221060
rect 270460 221048 270466 221060
rect 281994 221048 282000 221060
rect 270460 221020 282000 221048
rect 270460 221008 270466 221020
rect 281994 221008 282000 221020
rect 282052 221008 282058 221060
rect 282362 221008 282368 221060
rect 282420 221048 282426 221060
rect 282420 221020 284294 221048
rect 282420 221008 282426 221020
rect 233142 220980 233148 220992
rect 218026 220952 229692 220980
rect 229756 220952 233148 220980
rect 189868 220884 208256 220912
rect 189868 220872 189874 220884
rect 208302 220872 208308 220924
rect 208360 220912 208366 220924
rect 218026 220912 218054 220952
rect 208360 220884 218054 220912
rect 208360 220872 208366 220884
rect 219250 220872 219256 220924
rect 219308 220912 219314 220924
rect 220630 220912 220636 220924
rect 219308 220884 220636 220912
rect 219308 220872 219314 220884
rect 220630 220872 220636 220884
rect 220688 220872 220694 220924
rect 220814 220872 220820 220924
rect 220872 220912 220878 220924
rect 229554 220912 229560 220924
rect 220872 220884 229560 220912
rect 220872 220872 220878 220884
rect 229554 220872 229560 220884
rect 229612 220872 229618 220924
rect 229664 220912 229692 220952
rect 233142 220940 233148 220952
rect 233200 220940 233206 220992
rect 284266 220980 284294 221020
rect 284846 221008 284852 221060
rect 284904 221048 284910 221060
rect 290274 221048 290280 221060
rect 284904 221020 290280 221048
rect 284904 221008 284910 221020
rect 290274 221008 290280 221020
rect 290332 221008 290338 221060
rect 306282 221008 306288 221060
rect 306340 221048 306346 221060
rect 320358 221048 320364 221060
rect 306340 221020 320364 221048
rect 306340 221008 306346 221020
rect 320358 221008 320364 221020
rect 320416 221008 320422 221060
rect 329742 221008 329748 221060
rect 329800 221048 329806 221060
rect 346486 221048 346492 221060
rect 329800 221020 346492 221048
rect 329800 221008 329806 221020
rect 346486 221008 346492 221020
rect 346544 221008 346550 221060
rect 399294 221008 399300 221060
rect 399352 221048 399358 221060
rect 533982 221048 533988 221060
rect 399352 221020 533988 221048
rect 399352 221008 399358 221020
rect 533982 221008 533988 221020
rect 534040 221008 534046 221060
rect 542170 221008 542176 221060
rect 542228 221048 542234 221060
rect 543090 221048 543096 221060
rect 542228 221020 543096 221048
rect 542228 221008 542234 221020
rect 543090 221008 543096 221020
rect 543148 221048 543154 221060
rect 554406 221048 554412 221060
rect 543148 221020 554412 221048
rect 543148 221008 543154 221020
rect 554406 221008 554412 221020
rect 554464 221008 554470 221060
rect 555050 221008 555056 221060
rect 555108 221048 555114 221060
rect 556798 221048 556804 221060
rect 555108 221020 556804 221048
rect 555108 221008 555114 221020
rect 556798 221008 556804 221020
rect 556856 221008 556862 221060
rect 557534 221008 557540 221060
rect 557592 221048 557598 221060
rect 559282 221048 559288 221060
rect 557592 221020 559288 221048
rect 557592 221008 557598 221020
rect 559282 221008 559288 221020
rect 559340 221008 559346 221060
rect 563146 221008 563152 221060
rect 563204 221048 563210 221060
rect 564342 221048 564348 221060
rect 563204 221020 564348 221048
rect 563204 221008 563210 221020
rect 564342 221008 564348 221020
rect 564400 221008 564406 221060
rect 571702 221008 571708 221060
rect 571760 221048 571766 221060
rect 572714 221048 572720 221060
rect 571760 221020 572720 221048
rect 571760 221008 571766 221020
rect 572714 221008 572720 221020
rect 572772 221008 572778 221060
rect 572806 221008 572812 221060
rect 572864 221048 572870 221060
rect 619174 221048 619180 221060
rect 572864 221020 619180 221048
rect 572864 221008 572870 221020
rect 619174 221008 619180 221020
rect 619232 221008 619238 221060
rect 669590 221008 669596 221060
rect 669648 221048 669654 221060
rect 675846 221048 675852 221060
rect 669648 221020 675852 221048
rect 669648 221008 669654 221020
rect 675846 221008 675852 221020
rect 675904 221008 675910 221060
rect 287790 220980 287796 220992
rect 284266 220952 287796 220980
rect 287790 220940 287796 220952
rect 287848 220940 287854 220992
rect 289078 220940 289084 220992
rect 289136 220980 289142 220992
rect 290182 220980 290188 220992
rect 289136 220952 290188 220980
rect 289136 220940 289142 220952
rect 290182 220940 290188 220952
rect 290240 220940 290246 220992
rect 291562 220940 291568 220992
rect 291620 220980 291626 220992
rect 292758 220980 292764 220992
rect 291620 220952 292764 220980
rect 291620 220940 291626 220952
rect 292758 220940 292764 220952
rect 292816 220940 292822 220992
rect 311802 220940 311808 220992
rect 311860 220980 311866 220992
rect 327902 220980 327908 220992
rect 311860 220952 327908 220980
rect 311860 220940 311866 220952
rect 327902 220940 327908 220952
rect 327960 220940 327966 220992
rect 343266 220940 343272 220992
rect 343324 220980 343330 220992
rect 363230 220980 363236 220992
rect 343324 220952 363236 220980
rect 343324 220940 343330 220952
rect 363230 220940 363236 220952
rect 363288 220940 363294 220992
rect 396810 220940 396816 220992
rect 396868 220980 396874 220992
rect 534902 220980 534908 220992
rect 396868 220952 534908 220980
rect 396868 220940 396874 220952
rect 534902 220940 534908 220952
rect 534960 220940 534966 220992
rect 552198 220940 552204 220992
rect 552256 220980 552262 220992
rect 553670 220980 553676 220992
rect 552256 220952 553676 220980
rect 552256 220940 552262 220952
rect 553670 220940 553676 220952
rect 553728 220980 553734 220992
rect 618254 220980 618260 220992
rect 553728 220952 618260 220980
rect 553728 220940 553734 220952
rect 618254 220940 618260 220952
rect 618312 220940 618318 220992
rect 667106 220940 667112 220992
rect 667164 220980 667170 220992
rect 675938 220980 675944 220992
rect 667164 220952 675944 220980
rect 667164 220940 667170 220952
rect 675938 220940 675944 220952
rect 675996 220940 676002 220992
rect 233418 220912 233424 220924
rect 229664 220884 233424 220912
rect 233418 220872 233424 220884
rect 233476 220872 233482 220924
rect 233510 220872 233516 220924
rect 233568 220912 233574 220924
rect 238662 220912 238668 220924
rect 233568 220884 238668 220912
rect 233568 220872 233574 220884
rect 238662 220872 238668 220884
rect 238720 220872 238726 220924
rect 255406 220872 255412 220924
rect 255464 220912 255470 220924
rect 256602 220912 256608 220924
rect 255464 220884 256608 220912
rect 255464 220872 255470 220884
rect 256602 220872 256608 220884
rect 256660 220872 256666 220924
rect 261294 220872 261300 220924
rect 261352 220912 261358 220924
rect 262030 220912 262036 220924
rect 261352 220884 262036 220912
rect 261352 220872 261358 220884
rect 262030 220872 262036 220884
rect 262088 220872 262094 220924
rect 266354 220872 266360 220924
rect 266412 220912 266418 220924
rect 267458 220912 267464 220924
rect 266412 220884 267464 220912
rect 266412 220872 266418 220884
rect 267458 220872 267464 220884
rect 267516 220872 267522 220924
rect 273898 220872 273904 220924
rect 273956 220912 273962 220924
rect 284386 220912 284392 220924
rect 273956 220884 284392 220912
rect 273956 220872 273962 220884
rect 284386 220872 284392 220884
rect 284444 220872 284450 220924
rect 392210 220872 392216 220924
rect 392268 220912 392274 220924
rect 525058 220912 525064 220924
rect 392268 220884 525064 220912
rect 392268 220872 392274 220884
rect 525058 220872 525064 220884
rect 525116 220872 525122 220924
rect 548334 220872 548340 220924
rect 548392 220912 548398 220924
rect 617334 220912 617340 220924
rect 548392 220884 617340 220912
rect 548392 220872 548398 220884
rect 617334 220872 617340 220884
rect 617392 220872 617398 220924
rect 133414 220804 133420 220856
rect 133472 220844 133478 220856
rect 226886 220844 226892 220856
rect 133472 220816 226892 220844
rect 133472 220804 133478 220816
rect 226886 220804 226892 220816
rect 226944 220804 226950 220856
rect 232682 220804 232688 220856
rect 232740 220844 232746 220856
rect 234522 220844 234528 220856
rect 232740 220816 234528 220844
rect 232740 220804 232746 220816
rect 234522 220804 234528 220816
rect 234580 220804 234586 220856
rect 243630 220804 243636 220856
rect 243688 220844 243694 220856
rect 245562 220844 245568 220856
rect 243688 220816 245568 220844
rect 243688 220804 243694 220816
rect 245562 220804 245568 220816
rect 245620 220804 245626 220856
rect 248690 220804 248696 220856
rect 248748 220844 248754 220856
rect 251082 220844 251088 220856
rect 248748 220816 251088 220844
rect 248748 220804 248754 220816
rect 251082 220804 251088 220816
rect 251140 220804 251146 220856
rect 257890 220804 257896 220856
rect 257948 220844 257954 220856
rect 259270 220844 259276 220856
rect 257948 220816 259276 220844
rect 257948 220804 257954 220816
rect 259270 220804 259276 220816
rect 259328 220804 259334 220856
rect 262950 220804 262956 220856
rect 263008 220844 263014 220856
rect 264882 220844 264888 220856
rect 263008 220816 264888 220844
rect 263008 220804 263014 220816
rect 264882 220804 264888 220816
rect 264940 220804 264946 220856
rect 265526 220804 265532 220856
rect 265584 220844 265590 220856
rect 267642 220844 267648 220856
rect 265584 220816 267648 220844
rect 265584 220804 265590 220816
rect 267642 220804 267648 220816
rect 267700 220804 267706 220856
rect 268010 220804 268016 220856
rect 268068 220844 268074 220856
rect 281810 220844 281816 220856
rect 268068 220816 281816 220844
rect 268068 220804 268074 220816
rect 281810 220804 281816 220816
rect 281868 220804 281874 220856
rect 490190 220804 490196 220856
rect 490248 220844 490254 220856
rect 607122 220844 607128 220856
rect 490248 220816 607128 220844
rect 490248 220804 490254 220816
rect 607122 220804 607128 220816
rect 607180 220804 607186 220856
rect 46014 220328 46020 220380
rect 46072 220368 46078 220380
rect 647142 220368 647148 220380
rect 46072 220340 647148 220368
rect 46072 220328 46078 220340
rect 647142 220328 647148 220340
rect 647200 220328 647206 220380
rect 48498 220260 48504 220312
rect 48556 220300 48562 220312
rect 649902 220300 649908 220312
rect 48556 220272 649908 220300
rect 48556 220260 48562 220272
rect 649902 220260 649908 220272
rect 649960 220260 649966 220312
rect 46290 220192 46296 220244
rect 46348 220232 46354 220244
rect 648522 220232 648528 220244
rect 46348 220204 648528 220232
rect 46348 220192 46354 220204
rect 648522 220192 648528 220204
rect 648580 220192 648586 220244
rect 48590 220124 48596 220176
rect 48648 220164 48654 220176
rect 651282 220164 651288 220176
rect 48648 220136 651288 220164
rect 48648 220124 48654 220136
rect 651282 220124 651288 220136
rect 651340 220124 651346 220176
rect 652662 220124 652668 220176
rect 652720 220164 652726 220176
rect 675570 220164 675576 220176
rect 652720 220136 675576 220164
rect 652720 220124 652726 220136
rect 675570 220124 675576 220136
rect 675628 220164 675634 220176
rect 676030 220164 676036 220176
rect 675628 220136 676036 220164
rect 675628 220124 675634 220136
rect 676030 220124 676036 220136
rect 676088 220124 676094 220176
rect 48682 220056 48688 220108
rect 48740 220096 48746 220108
rect 652754 220096 652760 220108
rect 48740 220068 652760 220096
rect 48740 220056 48746 220068
rect 652754 220056 652760 220068
rect 652812 220056 652818 220108
rect 652846 220056 652852 220108
rect 652904 220096 652910 220108
rect 674834 220096 674840 220108
rect 652904 220068 674840 220096
rect 652904 220056 652910 220068
rect 674834 220056 674840 220068
rect 674892 220096 674898 220108
rect 675938 220096 675944 220108
rect 674892 220068 675944 220096
rect 674892 220056 674898 220068
rect 675938 220056 675944 220068
rect 675996 220056 676002 220108
rect 48866 219988 48872 220040
rect 48924 220028 48930 220040
rect 655514 220028 655520 220040
rect 48924 220000 655520 220028
rect 48924 219988 48930 220000
rect 655514 219988 655520 220000
rect 655572 219988 655578 220040
rect 48774 219920 48780 219972
rect 48832 219960 48838 219972
rect 654134 219960 654140 219972
rect 48832 219932 654140 219960
rect 48832 219920 48838 219932
rect 654134 219920 654140 219932
rect 654192 219920 654198 219972
rect 48958 219852 48964 219904
rect 49016 219892 49022 219904
rect 656894 219892 656900 219904
rect 49016 219864 656900 219892
rect 49016 219852 49022 219864
rect 656894 219852 656900 219864
rect 656952 219852 656958 219904
rect 46658 219784 46664 219836
rect 46716 219824 46722 219836
rect 658274 219824 658280 219836
rect 46716 219796 658280 219824
rect 46716 219784 46722 219796
rect 658274 219784 658280 219796
rect 658332 219784 658338 219836
rect 46750 219716 46756 219768
rect 46808 219756 46814 219768
rect 659746 219756 659752 219768
rect 46808 219728 659752 219756
rect 46808 219716 46814 219728
rect 659746 219716 659752 219728
rect 659804 219716 659810 219768
rect 46198 219648 46204 219700
rect 46256 219688 46262 219700
rect 661126 219688 661132 219700
rect 46256 219660 661132 219688
rect 46256 219648 46262 219660
rect 661126 219648 661132 219660
rect 661184 219648 661190 219700
rect 46106 219580 46112 219632
rect 46164 219620 46170 219632
rect 663426 219620 663432 219632
rect 46164 219592 663432 219620
rect 46164 219580 46170 219592
rect 663426 219580 663432 219592
rect 663484 219580 663490 219632
rect 45830 219512 45836 219564
rect 45888 219552 45894 219564
rect 664346 219552 664352 219564
rect 45888 219524 664352 219552
rect 45888 219512 45894 219524
rect 664346 219512 664352 219524
rect 664404 219512 664410 219564
rect 45922 219444 45928 219496
rect 45980 219484 45986 219496
rect 664806 219484 664812 219496
rect 45980 219456 664812 219484
rect 45980 219444 45986 219456
rect 664806 219444 664812 219456
rect 664864 219444 664870 219496
rect 45738 219376 45744 219428
rect 45796 219416 45802 219428
rect 663886 219416 663892 219428
rect 45796 219388 663892 219416
rect 45796 219376 45802 219388
rect 663886 219376 663892 219388
rect 663944 219376 663950 219428
rect 523402 218356 523408 218408
rect 523460 218396 523466 218408
rect 523770 218396 523776 218408
rect 523460 218368 523776 218396
rect 523460 218356 523466 218368
rect 523770 218356 523776 218368
rect 523828 218396 523834 218408
rect 612642 218396 612648 218408
rect 523828 218368 612648 218396
rect 523828 218356 523834 218368
rect 612642 218356 612648 218368
rect 612700 218356 612706 218408
rect 518986 218288 518992 218340
rect 519044 218328 519050 218340
rect 521194 218328 521200 218340
rect 519044 218300 521200 218328
rect 519044 218288 519050 218300
rect 521194 218288 521200 218300
rect 521252 218328 521258 218340
rect 612182 218328 612188 218340
rect 521252 218300 612188 218328
rect 521252 218288 521258 218300
rect 612182 218288 612188 218300
rect 612240 218288 612246 218340
rect 673914 218288 673920 218340
rect 673972 218328 673978 218340
rect 676030 218328 676036 218340
rect 673972 218300 676036 218328
rect 673972 218288 673978 218300
rect 676030 218288 676036 218300
rect 676088 218288 676094 218340
rect 518066 218220 518072 218272
rect 518124 218260 518130 218272
rect 518618 218260 518624 218272
rect 518124 218232 518624 218260
rect 518124 218220 518130 218232
rect 518618 218220 518624 218232
rect 518676 218260 518682 218272
rect 611722 218260 611728 218272
rect 518676 218232 611728 218260
rect 518676 218220 518682 218232
rect 611722 218220 611728 218232
rect 611780 218220 611786 218272
rect 515490 218152 515496 218204
rect 515548 218192 515554 218204
rect 611262 218192 611268 218204
rect 515548 218164 611268 218192
rect 515548 218152 515554 218164
rect 611262 218152 611268 218164
rect 611320 218152 611326 218204
rect 487154 218084 487160 218136
rect 487212 218124 487218 218136
rect 606662 218124 606668 218136
rect 487212 218096 606668 218124
rect 487212 218084 487218 218096
rect 606662 218084 606668 218096
rect 606720 218084 606726 218136
rect 662782 218084 662788 218136
rect 662840 218124 662846 218136
rect 662966 218124 662972 218136
rect 662840 218096 662972 218124
rect 662840 218084 662846 218096
rect 662966 218084 662972 218096
rect 663024 218084 663030 218136
rect 673454 218084 673460 218136
rect 673512 218124 673518 218136
rect 675938 218124 675944 218136
rect 673512 218096 675944 218124
rect 673512 218084 673518 218096
rect 675938 218084 675944 218096
rect 675996 218084 676002 218136
rect 46934 218016 46940 218068
rect 46992 218056 46998 218068
rect 671154 218056 671160 218068
rect 46992 218028 671160 218056
rect 46992 218016 46998 218028
rect 671154 218016 671160 218028
rect 671212 218016 671218 218068
rect 674374 218016 674380 218068
rect 674432 218056 674438 218068
rect 676030 218056 676036 218068
rect 674432 218028 676036 218056
rect 674432 218016 674438 218028
rect 676030 218016 676036 218028
rect 676088 218016 676094 218068
rect 646958 217948 646964 218000
rect 647016 217988 647022 218000
rect 651466 217988 651472 218000
rect 647016 217960 651472 217988
rect 647016 217948 647022 217960
rect 651466 217948 651472 217960
rect 651524 217948 651530 218000
rect 644106 217880 644112 217932
rect 644164 217920 644170 217932
rect 651558 217920 651564 217932
rect 644164 217892 651564 217920
rect 644164 217880 644170 217892
rect 651558 217880 651564 217892
rect 651616 217880 651622 217932
rect 507854 217608 507860 217660
rect 507912 217648 507918 217660
rect 509924 217648 509930 217660
rect 507912 217620 509930 217648
rect 507912 217608 507918 217620
rect 509924 217608 509930 217620
rect 509982 217608 509988 217660
rect 513834 217608 513840 217660
rect 513892 217648 513898 217660
rect 514984 217648 514990 217660
rect 513892 217620 514990 217648
rect 513892 217608 513898 217620
rect 514984 217608 514990 217620
rect 515042 217608 515048 217660
rect 502702 217472 502708 217524
rect 502760 217512 502766 217524
rect 504864 217512 504870 217524
rect 502760 217484 504870 217512
rect 502760 217472 502766 217484
rect 504864 217472 504870 217484
rect 504922 217472 504928 217524
rect 570552 217472 570558 217524
rect 570610 217512 570616 217524
rect 635918 217512 635924 217524
rect 570610 217484 635924 217512
rect 570610 217472 570616 217484
rect 635918 217472 635924 217484
rect 635976 217472 635982 217524
rect 568298 217404 568304 217456
rect 568356 217444 568362 217456
rect 635458 217444 635464 217456
rect 568356 217416 635464 217444
rect 568356 217404 568362 217416
rect 635458 217404 635464 217416
rect 635516 217404 635522 217456
rect 492582 217336 492588 217388
rect 492640 217376 492646 217388
rect 500310 217376 500316 217388
rect 492640 217348 500316 217376
rect 492640 217336 492646 217348
rect 500310 217336 500316 217348
rect 500368 217336 500374 217388
rect 565722 217336 565728 217388
rect 565780 217376 565786 217388
rect 634998 217376 635004 217388
rect 565780 217348 635004 217376
rect 565780 217336 565786 217348
rect 634998 217336 635004 217348
rect 635056 217336 635062 217388
rect 563054 217268 563060 217320
rect 563112 217308 563118 217320
rect 634538 217308 634544 217320
rect 563112 217280 634544 217308
rect 563112 217268 563118 217280
rect 634538 217268 634544 217280
rect 634596 217268 634602 217320
rect 550634 217200 550640 217252
rect 550692 217240 550698 217252
rect 632238 217240 632244 217252
rect 550692 217212 632244 217240
rect 550692 217200 550698 217212
rect 632238 217200 632244 217212
rect 632296 217200 632302 217252
rect 540514 217132 540520 217184
rect 540572 217172 540578 217184
rect 630398 217172 630404 217184
rect 540572 217144 630404 217172
rect 540572 217132 540578 217144
rect 630398 217132 630404 217144
rect 630456 217132 630462 217184
rect 530302 217064 530308 217116
rect 530360 217104 530366 217116
rect 628466 217104 628472 217116
rect 530360 217076 628472 217104
rect 530360 217064 530366 217076
rect 628466 217064 628472 217076
rect 628524 217064 628530 217116
rect 535362 216996 535368 217048
rect 535420 217036 535426 217048
rect 629478 217036 629484 217048
rect 535420 217008 629484 217036
rect 535420 216996 535426 217008
rect 629478 216996 629484 217008
rect 629536 216996 629542 217048
rect 525426 216928 525432 216980
rect 525484 216968 525490 216980
rect 627546 216968 627552 216980
rect 525484 216940 627552 216968
rect 525484 216928 525490 216940
rect 627546 216928 627552 216940
rect 627604 216928 627610 216980
rect 418522 216860 418528 216912
rect 418580 216900 418586 216912
rect 639690 216900 639696 216912
rect 418580 216872 639696 216900
rect 418580 216860 418586 216872
rect 639690 216860 639696 216872
rect 639748 216860 639754 216912
rect 520366 216792 520372 216844
rect 520424 216832 520430 216844
rect 626626 216832 626632 216844
rect 520424 216804 626632 216832
rect 520424 216792 520430 216804
rect 626626 216792 626632 216804
rect 626684 216792 626690 216844
rect 41506 216724 41512 216776
rect 41564 216764 41570 216776
rect 59354 216764 59360 216776
rect 41564 216736 59360 216764
rect 41564 216724 41570 216736
rect 59354 216724 59360 216736
rect 59412 216724 59418 216776
rect 418430 216724 418436 216776
rect 418488 216764 418494 216776
rect 640150 216764 640156 216776
rect 418488 216736 640156 216764
rect 418488 216724 418494 216736
rect 640150 216724 640156 216736
rect 640208 216724 640214 216776
rect 41414 216656 41420 216708
rect 41472 216696 41478 216708
rect 59446 216696 59452 216708
rect 41472 216668 59452 216696
rect 41472 216656 41478 216668
rect 59446 216656 59452 216668
rect 59504 216656 59510 216708
rect 418062 216656 418068 216708
rect 418120 216696 418126 216708
rect 641070 216696 641076 216708
rect 418120 216668 641076 216696
rect 418120 216656 418126 216668
rect 641070 216656 641076 216668
rect 641128 216656 641134 216708
rect 642726 216656 642732 216708
rect 642784 216696 642790 216708
rect 651374 216696 651380 216708
rect 642784 216668 651380 216696
rect 642784 216656 642790 216668
rect 651374 216656 651380 216668
rect 651432 216656 651438 216708
rect 674006 216656 674012 216708
rect 674064 216696 674070 216708
rect 675754 216696 675760 216708
rect 674064 216668 675760 216696
rect 674064 216656 674070 216668
rect 675754 216656 675760 216668
rect 675812 216656 675818 216708
rect 41598 216588 41604 216640
rect 41656 216628 41662 216640
rect 59262 216628 59268 216640
rect 41656 216600 59268 216628
rect 41656 216588 41662 216600
rect 59262 216588 59268 216600
rect 59320 216588 59326 216640
rect 418154 216588 418160 216640
rect 418212 216628 418218 216640
rect 640610 216628 640616 216640
rect 418212 216600 640616 216628
rect 418212 216588 418218 216600
rect 640610 216588 640616 216600
rect 640668 216588 640674 216640
rect 495986 216520 495992 216572
rect 496044 216560 496050 216572
rect 496044 216532 502656 216560
rect 496044 216520 496050 216532
rect 496998 216452 497004 216504
rect 497056 216492 497062 216504
rect 499298 216492 499304 216504
rect 497056 216464 499304 216492
rect 497056 216452 497062 216464
rect 499298 216452 499304 216464
rect 499356 216492 499362 216504
rect 502518 216492 502524 216504
rect 499356 216464 502524 216492
rect 499356 216452 499362 216464
rect 502518 216452 502524 216464
rect 502576 216452 502582 216504
rect 484210 216384 484216 216436
rect 484268 216384 484274 216436
rect 486694 216384 486700 216436
rect 486752 216424 486758 216436
rect 486752 216396 488534 216424
rect 486752 216384 486758 216396
rect 484228 215948 484256 216384
rect 488506 216016 488534 216396
rect 490098 216384 490104 216436
rect 490156 216424 490162 216436
rect 490156 216396 492444 216424
rect 490156 216384 490162 216396
rect 492416 216084 492444 216396
rect 500218 216384 500224 216436
rect 500276 216384 500282 216436
rect 500310 216384 500316 216436
rect 500368 216424 500374 216436
rect 500368 216396 502564 216424
rect 500368 216384 500374 216396
rect 500236 216152 500264 216384
rect 502536 216220 502564 216396
rect 502628 216288 502656 216532
rect 505002 216520 505008 216572
rect 505060 216560 505066 216572
rect 505060 216532 507900 216560
rect 505060 216520 505066 216532
rect 502702 216384 502708 216436
rect 502760 216424 502766 216436
rect 507872 216424 507900 216532
rect 515122 216520 515128 216572
rect 515180 216560 515186 216572
rect 625706 216560 625712 216572
rect 515180 216532 625712 216560
rect 515180 216520 515186 216532
rect 625706 216520 625712 216532
rect 625764 216520 625770 216572
rect 510246 216452 510252 216504
rect 510304 216492 510310 216504
rect 624786 216492 624792 216504
rect 510304 216464 624792 216492
rect 510304 216452 510310 216464
rect 624786 216452 624792 216464
rect 624844 216452 624850 216504
rect 623866 216424 623872 216436
rect 502760 216396 502840 216424
rect 507872 216396 623872 216424
rect 502760 216384 502766 216396
rect 502812 216356 502840 216396
rect 623866 216384 623872 216396
rect 623924 216384 623930 216436
rect 622946 216356 622952 216368
rect 502812 216328 622952 216356
rect 622946 216316 622952 216328
rect 623004 216316 623010 216368
rect 622486 216288 622492 216300
rect 502628 216260 622492 216288
rect 622486 216248 622492 216260
rect 622544 216248 622550 216300
rect 645578 216248 645584 216300
rect 645636 216288 645642 216300
rect 651650 216288 651656 216300
rect 645636 216260 651656 216288
rect 645636 216248 645642 216260
rect 651650 216248 651656 216260
rect 651708 216248 651714 216300
rect 673822 216248 673828 216300
rect 673880 216288 673886 216300
rect 676030 216288 676036 216300
rect 673880 216260 676036 216288
rect 673880 216248 673886 216260
rect 676030 216248 676036 216260
rect 676088 216248 676094 216300
rect 622026 216220 622032 216232
rect 502536 216192 622032 216220
rect 622026 216180 622032 216192
rect 622084 216180 622090 216232
rect 637850 216152 637856 216164
rect 500236 216124 637856 216152
rect 637850 216112 637856 216124
rect 637908 216112 637914 216164
rect 636378 216084 636384 216096
rect 492416 216056 636384 216084
rect 636378 216044 636384 216056
rect 636436 216044 636442 216096
rect 638310 216016 638316 216028
rect 488506 215988 638316 216016
rect 638310 215976 638316 215988
rect 638368 215976 638374 216028
rect 638770 215948 638776 215960
rect 484228 215920 638776 215948
rect 638770 215908 638776 215920
rect 638828 215908 638834 215960
rect 48222 215840 48228 215892
rect 48280 215880 48286 215892
rect 665726 215880 665732 215892
rect 48280 215852 665732 215880
rect 48280 215840 48286 215852
rect 665726 215840 665732 215852
rect 665784 215840 665790 215892
rect 673546 215840 673552 215892
rect 673604 215880 673610 215892
rect 675938 215880 675944 215892
rect 673604 215852 675944 215880
rect 673604 215840 673610 215852
rect 675938 215840 675944 215852
rect 675996 215840 676002 215892
rect 31846 215772 31852 215824
rect 31904 215812 31910 215824
rect 666186 215812 666192 215824
rect 31904 215784 666192 215812
rect 31904 215772 31910 215784
rect 666186 215772 666192 215784
rect 666244 215772 666250 215824
rect 31662 215704 31668 215756
rect 31720 215744 31726 215756
rect 665266 215744 665272 215756
rect 31720 215716 665272 215744
rect 31720 215704 31726 215716
rect 665266 215704 665272 215716
rect 665324 215704 665330 215756
rect 579706 215636 579712 215688
rect 579764 215676 579770 215688
rect 599762 215676 599768 215688
rect 579764 215648 599768 215676
rect 579764 215636 579770 215648
rect 599762 215636 599768 215648
rect 599820 215636 599826 215688
rect 674098 215432 674104 215484
rect 674156 215472 674162 215484
rect 675846 215472 675852 215484
rect 674156 215444 675852 215472
rect 674156 215432 674162 215444
rect 675846 215432 675852 215444
rect 675904 215432 675910 215484
rect 674190 215364 674196 215416
rect 674248 215404 674254 215416
rect 675938 215404 675944 215416
rect 674248 215376 675944 215404
rect 674248 215364 674254 215376
rect 675938 215364 675944 215376
rect 675996 215364 676002 215416
rect 675202 215296 675208 215348
rect 675260 215336 675266 215348
rect 676030 215336 676036 215348
rect 675260 215308 676036 215336
rect 675260 215296 675266 215308
rect 676030 215296 676036 215308
rect 676088 215296 676094 215348
rect 673638 214616 673644 214668
rect 673696 214656 673702 214668
rect 676030 214656 676036 214668
rect 673696 214628 676036 214656
rect 673696 214616 673702 214628
rect 676030 214616 676036 214628
rect 676088 214616 676094 214668
rect 41506 213868 41512 213920
rect 41564 213908 41570 213920
rect 45554 213908 45560 213920
rect 41564 213880 45560 213908
rect 41564 213868 41570 213880
rect 45554 213868 45560 213880
rect 45612 213868 45618 213920
rect 673730 213800 673736 213852
rect 673788 213840 673794 213852
rect 675938 213840 675944 213852
rect 673788 213812 675944 213840
rect 673788 213800 673794 213812
rect 675938 213800 675944 213812
rect 675996 213800 676002 213852
rect 41506 213664 41512 213716
rect 41564 213704 41570 213716
rect 43438 213704 43444 213716
rect 41564 213676 43444 213704
rect 41564 213664 41570 213676
rect 43438 213664 43444 213676
rect 43496 213664 43502 213716
rect 674650 212848 674656 212900
rect 674708 212888 674714 212900
rect 674708 212860 674788 212888
rect 674708 212848 674714 212860
rect 674760 212696 674788 212860
rect 674742 212644 674748 212696
rect 674800 212644 674806 212696
rect 582282 212576 582288 212628
rect 582340 212616 582346 212628
rect 599946 212616 599952 212628
rect 582340 212588 599952 212616
rect 582340 212576 582346 212588
rect 599946 212576 599952 212588
rect 600004 212576 600010 212628
rect 674650 212576 674656 212628
rect 674708 212616 674714 212628
rect 675938 212616 675944 212628
rect 674708 212588 675944 212616
rect 674708 212576 674714 212588
rect 675938 212576 675944 212588
rect 675996 212576 676002 212628
rect 580258 212508 580264 212560
rect 580316 212548 580322 212560
rect 599854 212548 599860 212560
rect 580316 212520 599860 212548
rect 580316 212508 580322 212520
rect 599854 212508 599860 212520
rect 599912 212508 599918 212560
rect 674466 212508 674472 212560
rect 674524 212548 674530 212560
rect 676030 212548 676036 212560
rect 674524 212520 676036 212548
rect 674524 212508 674530 212520
rect 676030 212508 676036 212520
rect 676088 212508 676094 212560
rect 651282 212440 651288 212492
rect 651340 212480 651346 212492
rect 651374 212480 651380 212492
rect 651340 212452 651380 212480
rect 651340 212440 651346 212452
rect 651374 212440 651380 212452
rect 651432 212440 651438 212492
rect 673178 212440 673184 212492
rect 673236 212480 673242 212492
rect 675386 212480 675392 212492
rect 673236 212452 675392 212480
rect 673236 212440 673242 212452
rect 675386 212440 675392 212452
rect 675444 212440 675450 212492
rect 581638 209856 581644 209908
rect 581696 209896 581702 209908
rect 600038 209896 600044 209908
rect 581696 209868 600044 209896
rect 581696 209856 581702 209868
rect 600038 209856 600044 209868
rect 600096 209856 600102 209908
rect 580534 209788 580540 209840
rect 580592 209828 580598 209840
rect 599118 209828 599124 209840
rect 580592 209800 599124 209828
rect 580592 209788 580598 209800
rect 599118 209788 599124 209800
rect 599176 209788 599182 209840
rect 674282 208360 674288 208412
rect 674340 208400 674346 208412
rect 675570 208400 675576 208412
rect 674340 208372 675576 208400
rect 674340 208360 674346 208372
rect 675570 208360 675576 208372
rect 675628 208360 675634 208412
rect 674834 208292 674840 208344
rect 674892 208332 674898 208344
rect 675202 208332 675208 208344
rect 674892 208304 675208 208332
rect 674892 208292 674898 208304
rect 675202 208292 675208 208304
rect 675260 208292 675266 208344
rect 582282 207068 582288 207120
rect 582340 207108 582346 207120
rect 601142 207108 601148 207120
rect 582340 207080 601148 207108
rect 582340 207068 582346 207080
rect 601142 207068 601148 207080
rect 601200 207068 601206 207120
rect 581454 207000 581460 207052
rect 581512 207040 581518 207052
rect 600958 207040 600964 207052
rect 581512 207012 600964 207040
rect 581512 207000 581518 207012
rect 600958 207000 600964 207012
rect 601016 207000 601022 207052
rect 675662 205980 675668 206032
rect 675720 205980 675726 206032
rect 675754 205980 675760 206032
rect 675812 205980 675818 206032
rect 674374 205504 674380 205556
rect 674432 205544 674438 205556
rect 675294 205544 675300 205556
rect 674432 205516 675300 205544
rect 674432 205504 674438 205516
rect 675294 205504 675300 205516
rect 675352 205504 675358 205556
rect 674374 205368 674380 205420
rect 674432 205408 674438 205420
rect 675680 205408 675708 205980
rect 674432 205380 675708 205408
rect 674432 205368 674438 205380
rect 673914 205164 673920 205216
rect 673972 205204 673978 205216
rect 675294 205204 675300 205216
rect 673972 205176 675300 205204
rect 673972 205164 673978 205176
rect 675294 205164 675300 205176
rect 675352 205164 675358 205216
rect 675772 205012 675800 205980
rect 675754 204960 675760 205012
rect 675812 204960 675818 205012
rect 582282 204280 582288 204332
rect 582340 204320 582346 204332
rect 599946 204320 599952 204332
rect 582340 204292 599952 204320
rect 582340 204280 582346 204292
rect 599946 204280 599952 204292
rect 600004 204280 600010 204332
rect 673822 202716 673828 202768
rect 673880 202756 673886 202768
rect 675478 202756 675484 202768
rect 673880 202728 675484 202756
rect 673880 202716 673886 202728
rect 675478 202716 675484 202728
rect 675536 202716 675542 202768
rect 673638 202580 673644 202632
rect 673696 202620 673702 202632
rect 673822 202620 673828 202632
rect 673696 202592 673828 202620
rect 673696 202580 673702 202592
rect 673822 202580 673828 202592
rect 673880 202580 673886 202632
rect 673546 202308 673552 202360
rect 673604 202348 673610 202360
rect 674374 202348 674380 202360
rect 673604 202320 674380 202348
rect 673604 202308 673610 202320
rect 674374 202308 674380 202320
rect 674432 202308 674438 202360
rect 674834 202036 674840 202088
rect 674892 202076 674898 202088
rect 675386 202076 675392 202088
rect 674892 202048 675392 202076
rect 674892 202036 674898 202048
rect 675386 202036 675392 202048
rect 675444 202036 675450 202088
rect 674098 201900 674104 201952
rect 674156 201940 674162 201952
rect 674834 201940 674840 201952
rect 674156 201912 674840 201940
rect 674156 201900 674162 201912
rect 674834 201900 674840 201912
rect 674892 201900 674898 201952
rect 581822 201560 581828 201612
rect 581880 201600 581886 201612
rect 599026 201600 599032 201612
rect 581880 201572 599032 201600
rect 581880 201560 581886 201572
rect 599026 201560 599032 201572
rect 599084 201560 599090 201612
rect 581086 201492 581092 201544
rect 581144 201532 581150 201544
rect 599946 201532 599952 201544
rect 581144 201504 599952 201532
rect 581144 201492 581150 201504
rect 599946 201492 599952 201504
rect 600004 201492 600010 201544
rect 674190 201492 674196 201544
rect 674248 201532 674254 201544
rect 675386 201532 675392 201544
rect 674248 201504 675392 201532
rect 674248 201492 674254 201504
rect 675386 201492 675392 201504
rect 675444 201492 675450 201544
rect 674466 200880 674472 200932
rect 674524 200920 674530 200932
rect 675386 200920 675392 200932
rect 674524 200892 675392 200920
rect 674524 200880 674530 200892
rect 675386 200880 675392 200892
rect 675444 200880 675450 200932
rect 33042 200200 33048 200252
rect 33100 200240 33106 200252
rect 41874 200240 41880 200252
rect 33100 200212 41880 200240
rect 33100 200200 33106 200212
rect 41874 200200 41880 200212
rect 41932 200200 41938 200252
rect 581086 200064 581092 200116
rect 581144 200104 581150 200116
rect 599946 200104 599952 200116
rect 581144 200076 599952 200104
rect 581144 200064 581150 200076
rect 599946 200064 599952 200076
rect 600004 200064 600010 200116
rect 32950 199996 32956 200048
rect 33008 200036 33014 200048
rect 42518 200036 42524 200048
rect 33008 200008 42524 200036
rect 33008 199996 33014 200008
rect 42518 199996 42524 200008
rect 42576 199996 42582 200048
rect 582282 198704 582288 198756
rect 582340 198744 582346 198756
rect 599118 198744 599124 198756
rect 582340 198716 599124 198744
rect 582340 198704 582346 198716
rect 599118 198704 599124 198716
rect 599176 198704 599182 198756
rect 673638 198364 673644 198416
rect 673696 198404 673702 198416
rect 675386 198404 675392 198416
rect 673696 198376 675392 198404
rect 673696 198364 673702 198376
rect 675386 198364 675392 198376
rect 675444 198364 675450 198416
rect 673730 197548 673736 197600
rect 673788 197588 673794 197600
rect 675478 197588 675484 197600
rect 673788 197560 675484 197588
rect 673788 197548 673794 197560
rect 675478 197548 675484 197560
rect 675536 197548 675542 197600
rect 41874 197412 41880 197464
rect 41932 197412 41938 197464
rect 41892 197192 41920 197412
rect 580810 197344 580816 197396
rect 580868 197384 580874 197396
rect 599302 197384 599308 197396
rect 580868 197356 599308 197384
rect 580868 197344 580874 197356
rect 599302 197344 599308 197356
rect 599360 197344 599366 197396
rect 581270 197276 581276 197328
rect 581328 197316 581334 197328
rect 599946 197316 599952 197328
rect 581328 197288 599952 197316
rect 581328 197276 581334 197288
rect 599946 197276 599952 197288
rect 600004 197276 600010 197328
rect 41874 197140 41880 197192
rect 41932 197140 41938 197192
rect 673822 197004 673828 197056
rect 673880 197044 673886 197056
rect 675386 197044 675392 197056
rect 673880 197016 675392 197044
rect 673880 197004 673886 197016
rect 675386 197004 675392 197016
rect 675444 197004 675450 197056
rect 674650 196528 674656 196580
rect 674708 196568 674714 196580
rect 675386 196568 675392 196580
rect 674708 196540 675392 196568
rect 674708 196528 674714 196540
rect 675386 196528 675392 196540
rect 675444 196528 675450 196580
rect 674466 196392 674472 196444
rect 674524 196432 674530 196444
rect 674650 196432 674656 196444
rect 674524 196404 674656 196432
rect 674524 196392 674530 196404
rect 674650 196392 674656 196404
rect 674708 196392 674714 196444
rect 674834 195304 674840 195356
rect 674892 195344 674898 195356
rect 675386 195344 675392 195356
rect 674892 195316 675392 195344
rect 674892 195304 674898 195316
rect 675386 195304 675392 195316
rect 675444 195304 675450 195356
rect 42150 195236 42156 195288
rect 42208 195276 42214 195288
rect 42518 195276 42524 195288
rect 42208 195248 42524 195276
rect 42208 195236 42214 195248
rect 42518 195236 42524 195248
rect 42576 195236 42582 195288
rect 674374 195168 674380 195220
rect 674432 195208 674438 195220
rect 674834 195208 674840 195220
rect 674432 195180 674840 195208
rect 674432 195168 674438 195180
rect 674834 195168 674840 195180
rect 674892 195168 674898 195220
rect 582190 194624 582196 194676
rect 582248 194664 582254 194676
rect 599118 194664 599124 194676
rect 582248 194636 599124 194664
rect 582248 194624 582254 194636
rect 599118 194624 599124 194636
rect 599176 194624 599182 194676
rect 582282 194556 582288 194608
rect 582340 194596 582346 194608
rect 599946 194596 599952 194608
rect 582340 194568 599952 194596
rect 582340 194556 582346 194568
rect 599946 194556 599952 194568
rect 600004 194556 600010 194608
rect 42058 193468 42064 193520
rect 42116 193508 42122 193520
rect 42886 193508 42892 193520
rect 42116 193480 42892 193508
rect 42116 193468 42122 193480
rect 42886 193468 42892 193480
rect 42944 193468 42950 193520
rect 673454 193468 673460 193520
rect 673512 193508 673518 193520
rect 675386 193508 675392 193520
rect 673512 193480 675392 193508
rect 673512 193468 673518 193480
rect 675386 193468 675392 193480
rect 675444 193468 675450 193520
rect 42150 192176 42156 192228
rect 42208 192216 42214 192228
rect 42794 192216 42800 192228
rect 42208 192188 42800 192216
rect 42208 192176 42214 192188
rect 42794 192176 42800 192188
rect 42852 192176 42858 192228
rect 582282 191836 582288 191888
rect 582340 191876 582346 191888
rect 599854 191876 599860 191888
rect 582340 191848 599860 191876
rect 582340 191836 582346 191848
rect 599854 191836 599860 191848
rect 599912 191836 599918 191888
rect 581270 191768 581276 191820
rect 581328 191808 581334 191820
rect 599946 191808 599952 191820
rect 581328 191780 599952 191808
rect 581328 191768 581334 191780
rect 599946 191768 599952 191780
rect 600004 191768 600010 191820
rect 673546 191632 673552 191684
rect 673604 191672 673610 191684
rect 675386 191672 675392 191684
rect 673604 191644 675392 191672
rect 673604 191632 673610 191644
rect 675386 191632 675392 191644
rect 675444 191632 675450 191684
rect 42058 191428 42064 191480
rect 42116 191468 42122 191480
rect 43070 191468 43076 191480
rect 42116 191440 43076 191468
rect 42116 191428 42122 191440
rect 43070 191428 43076 191440
rect 43128 191428 43134 191480
rect 42150 190952 42156 191004
rect 42208 190992 42214 191004
rect 42978 190992 42984 191004
rect 42208 190964 42984 190992
rect 42208 190952 42214 190964
rect 42978 190952 42984 190964
rect 43036 190952 43042 191004
rect 579706 190408 579712 190460
rect 579764 190448 579770 190460
rect 599854 190448 599860 190460
rect 579764 190420 599860 190448
rect 579764 190408 579770 190420
rect 599854 190408 599860 190420
rect 599912 190408 599918 190460
rect 582190 187620 582196 187672
rect 582248 187660 582254 187672
rect 601602 187660 601608 187672
rect 582248 187632 601608 187660
rect 582248 187620 582254 187632
rect 601602 187620 601608 187632
rect 601660 187620 601666 187672
rect 582282 187552 582288 187604
rect 582340 187592 582346 187604
rect 600958 187592 600964 187604
rect 582340 187564 600964 187592
rect 582340 187552 582346 187564
rect 600958 187552 600964 187564
rect 601016 187552 601022 187604
rect 580258 184832 580264 184884
rect 580316 184872 580322 184884
rect 599946 184872 599952 184884
rect 580316 184844 599952 184872
rect 580316 184832 580322 184844
rect 599946 184832 599952 184844
rect 600004 184832 600010 184884
rect 580902 184764 580908 184816
rect 580960 184804 580966 184816
rect 601510 184804 601516 184816
rect 580960 184776 601516 184804
rect 580960 184764 580966 184776
rect 601510 184764 601516 184776
rect 601568 184764 601574 184816
rect 666738 183880 666744 183932
rect 666796 183920 666802 183932
rect 667106 183920 667112 183932
rect 666796 183892 667112 183920
rect 666796 183880 666802 183892
rect 667106 183880 667112 183892
rect 667164 183880 667170 183932
rect 581822 182112 581828 182164
rect 581880 182152 581886 182164
rect 599854 182152 599860 182164
rect 581880 182124 599860 182152
rect 581880 182112 581886 182124
rect 599854 182112 599860 182124
rect 599912 182112 599918 182164
rect 580534 182044 580540 182096
rect 580592 182084 580598 182096
rect 600038 182084 600044 182096
rect 580592 182056 600044 182084
rect 580592 182044 580598 182056
rect 600038 182044 600044 182056
rect 600096 182044 600102 182096
rect 708506 179500 708512 179512
rect 704384 179472 708512 179500
rect 704384 179376 704412 179472
rect 708506 179460 708512 179472
rect 708564 179460 708570 179512
rect 704458 179392 704464 179444
rect 704516 179432 704522 179444
rect 708414 179432 708420 179444
rect 704516 179404 708420 179432
rect 704516 179392 704522 179404
rect 708414 179392 708420 179404
rect 708472 179392 708478 179444
rect 580718 179324 580724 179376
rect 580776 179364 580782 179376
rect 599946 179364 599952 179376
rect 580776 179336 599952 179364
rect 580776 179324 580782 179336
rect 599946 179324 599952 179336
rect 600004 179324 600010 179376
rect 666922 179324 666928 179376
rect 666980 179364 666986 179376
rect 671430 179364 671436 179376
rect 666980 179336 671436 179364
rect 666980 179324 666986 179336
rect 671430 179324 671436 179336
rect 671488 179324 671494 179376
rect 674742 179324 674748 179376
rect 674800 179364 674806 179376
rect 675846 179364 675852 179376
rect 674800 179336 675852 179364
rect 674800 179324 674806 179336
rect 675846 179324 675852 179336
rect 675904 179324 675910 179376
rect 704366 179324 704372 179376
rect 704424 179324 704430 179376
rect 707494 179364 707500 179376
rect 705488 179336 707500 179364
rect 581086 179256 581092 179308
rect 581144 179296 581150 179308
rect 599762 179296 599768 179308
rect 581144 179268 599768 179296
rect 581144 179256 581150 179268
rect 599762 179256 599768 179268
rect 599820 179256 599826 179308
rect 705286 179188 705292 179240
rect 705344 179228 705350 179240
rect 705488 179228 705516 179336
rect 707494 179324 707500 179336
rect 707552 179324 707558 179376
rect 707034 179296 707040 179308
rect 705764 179268 707040 179296
rect 705764 179240 705792 179268
rect 707034 179256 707040 179268
rect 707092 179256 707098 179308
rect 705344 179200 705516 179228
rect 705344 179188 705350 179200
rect 705746 179188 705752 179240
rect 705804 179188 705810 179240
rect 706206 179188 706212 179240
rect 706264 179228 706270 179240
rect 706666 179228 706672 179240
rect 706264 179200 706672 179228
rect 706264 179188 706270 179200
rect 706666 179188 706672 179200
rect 706724 179188 706730 179240
rect 706298 179120 706304 179172
rect 706356 179160 706362 179172
rect 706574 179160 706580 179172
rect 706356 179132 706580 179160
rect 706356 179120 706362 179132
rect 706574 179120 706580 179132
rect 706632 179120 706638 179172
rect 705838 179052 705844 179104
rect 705896 179092 705902 179104
rect 707034 179092 707040 179104
rect 705896 179064 707040 179092
rect 705896 179052 705902 179064
rect 707034 179052 707040 179064
rect 707092 179052 707098 179104
rect 705378 178984 705384 179036
rect 705436 179024 705442 179036
rect 707494 179024 707500 179036
rect 705436 178996 707500 179024
rect 705436 178984 705442 178996
rect 707494 178984 707500 178996
rect 707552 178984 707558 179036
rect 708046 178984 708052 179036
rect 708104 178984 708110 179036
rect 704918 178916 704924 178968
rect 704976 178956 704982 178968
rect 707954 178956 707960 178968
rect 704976 178928 707960 178956
rect 704976 178916 704982 178928
rect 707954 178916 707960 178928
rect 708012 178916 708018 178968
rect 704826 178848 704832 178900
rect 704884 178888 704890 178900
rect 708064 178888 708092 178984
rect 704884 178860 708092 178888
rect 704884 178848 704890 178860
rect 703998 178780 704004 178832
rect 704056 178820 704062 178832
rect 708874 178820 708880 178832
rect 704056 178792 708880 178820
rect 704056 178780 704062 178792
rect 708874 178780 708880 178792
rect 708932 178780 708938 178832
rect 669406 177080 669412 177132
rect 669464 177120 669470 177132
rect 675938 177120 675944 177132
rect 669464 177092 675944 177120
rect 669464 177080 669470 177092
rect 675938 177080 675944 177092
rect 675996 177080 676002 177132
rect 669130 176944 669136 176996
rect 669188 176984 669194 176996
rect 676030 176984 676036 176996
rect 669188 176956 676036 176984
rect 669188 176944 669194 176956
rect 676030 176944 676036 176956
rect 676088 176944 676094 176996
rect 671430 176876 671436 176928
rect 671488 176916 671494 176928
rect 673270 176916 673276 176928
rect 671488 176888 673276 176916
rect 671488 176876 671494 176888
rect 673270 176876 673276 176888
rect 673328 176916 673334 176928
rect 675938 176916 675944 176928
rect 673328 176888 675944 176916
rect 673328 176876 673334 176888
rect 675938 176876 675944 176888
rect 675996 176876 676002 176928
rect 667014 176808 667020 176860
rect 667072 176848 667078 176860
rect 675754 176848 675760 176860
rect 667072 176820 675760 176848
rect 667072 176808 667078 176820
rect 675754 176808 675760 176820
rect 675812 176808 675818 176860
rect 581086 176672 581092 176724
rect 581144 176712 581150 176724
rect 598934 176712 598940 176724
rect 581144 176684 598940 176712
rect 581144 176672 581150 176684
rect 598934 176672 598940 176684
rect 598992 176672 598998 176724
rect 581454 176604 581460 176656
rect 581512 176644 581518 176656
rect 599854 176644 599860 176656
rect 581512 176616 599860 176644
rect 581512 176604 581518 176616
rect 599854 176604 599860 176616
rect 599912 176604 599918 176656
rect 666830 176604 666836 176656
rect 666888 176644 666894 176656
rect 671890 176644 671896 176656
rect 666888 176616 671896 176644
rect 666888 176604 666894 176616
rect 671890 176604 671896 176616
rect 671948 176604 671954 176656
rect 674834 176604 674840 176656
rect 674892 176644 674898 176656
rect 676030 176644 676036 176656
rect 674892 176616 676036 176644
rect 674892 176604 674898 176616
rect 676030 176604 676036 176616
rect 676088 176604 676094 176656
rect 667106 176536 667112 176588
rect 667164 176576 667170 176588
rect 672166 176576 672172 176588
rect 667164 176548 672172 176576
rect 667164 176536 667170 176548
rect 672166 176536 672172 176548
rect 672224 176536 672230 176588
rect 674558 176332 674564 176384
rect 674616 176372 674622 176384
rect 676030 176372 676036 176384
rect 674616 176344 676036 176372
rect 674616 176332 674622 176344
rect 676030 176332 676036 176344
rect 676088 176332 676094 176384
rect 673362 175992 673368 176044
rect 673420 176032 673426 176044
rect 675938 176032 675944 176044
rect 673420 176004 675944 176032
rect 673420 175992 673426 176004
rect 675938 175992 675944 176004
rect 675996 175992 676002 176044
rect 674650 175516 674656 175568
rect 674708 175556 674714 175568
rect 676030 175556 676036 175568
rect 674708 175528 676036 175556
rect 674708 175516 674714 175528
rect 676030 175516 676036 175528
rect 676088 175516 676094 175568
rect 671890 175244 671896 175296
rect 671948 175284 671954 175296
rect 672258 175284 672264 175296
rect 671948 175256 672264 175284
rect 671948 175244 671954 175256
rect 672258 175244 672264 175256
rect 672316 175284 672322 175296
rect 675938 175284 675944 175296
rect 672316 175256 675944 175284
rect 672316 175244 672322 175256
rect 675938 175244 675944 175256
rect 675996 175244 676002 175296
rect 671890 174428 671896 174480
rect 671948 174468 671954 174480
rect 672166 174468 672172 174480
rect 671948 174440 672172 174468
rect 671948 174428 671954 174440
rect 672166 174428 672172 174440
rect 672224 174468 672230 174480
rect 676030 174468 676036 174480
rect 672224 174440 676036 174468
rect 672224 174428 672230 174440
rect 676030 174428 676036 174440
rect 676088 174428 676094 174480
rect 580810 173884 580816 173936
rect 580868 173924 580874 173936
rect 599946 173924 599952 173936
rect 580868 173896 599952 173924
rect 580868 173884 580874 173896
rect 599946 173884 599952 173896
rect 600004 173884 600010 173936
rect 674098 173884 674104 173936
rect 674156 173924 674162 173936
rect 676030 173924 676036 173936
rect 674156 173896 676036 173924
rect 674156 173884 674162 173896
rect 676030 173884 676036 173896
rect 676088 173884 676094 173936
rect 579706 173816 579712 173868
rect 579764 173856 579770 173868
rect 600038 173856 600044 173868
rect 579764 173828 600044 173856
rect 579764 173816 579770 173828
rect 600038 173816 600044 173828
rect 600096 173816 600102 173868
rect 582282 173748 582288 173800
rect 582340 173788 582346 173800
rect 600130 173788 600136 173800
rect 582340 173760 600136 173788
rect 582340 173748 582346 173760
rect 600130 173748 600136 173760
rect 600188 173748 600194 173800
rect 674834 171640 674840 171692
rect 674892 171680 674898 171692
rect 676030 171680 676036 171692
rect 674892 171652 676036 171680
rect 674892 171640 674898 171652
rect 676030 171640 676036 171652
rect 676088 171640 676094 171692
rect 673454 171300 673460 171352
rect 673512 171340 673518 171352
rect 675938 171340 675944 171352
rect 673512 171312 675944 171340
rect 673512 171300 673518 171312
rect 675938 171300 675944 171312
rect 675996 171300 676002 171352
rect 582190 171164 582196 171216
rect 582248 171204 582254 171216
rect 599946 171204 599952 171216
rect 582248 171176 599952 171204
rect 582248 171164 582254 171176
rect 599946 171164 599952 171176
rect 600004 171164 600010 171216
rect 674558 171164 674564 171216
rect 674616 171204 674622 171216
rect 675938 171204 675944 171216
rect 674616 171176 675944 171204
rect 674616 171164 674622 171176
rect 675938 171164 675944 171176
rect 675996 171164 676002 171216
rect 579890 171096 579896 171148
rect 579948 171136 579954 171148
rect 599854 171136 599860 171148
rect 579948 171108 599860 171136
rect 579948 171096 579954 171108
rect 599854 171096 599860 171108
rect 599912 171096 599918 171148
rect 676030 171136 676036 171148
rect 675220 171108 676036 171136
rect 580902 171028 580908 171080
rect 580960 171068 580966 171080
rect 599670 171068 599676 171080
rect 580960 171040 599676 171068
rect 580960 171028 580966 171040
rect 599670 171028 599676 171040
rect 599728 171028 599734 171080
rect 675220 171012 675248 171108
rect 676030 171096 676036 171108
rect 676088 171096 676094 171148
rect 580074 170960 580080 171012
rect 580132 171000 580138 171012
rect 599762 171000 599768 171012
rect 580132 170972 599768 171000
rect 580132 170960 580138 170972
rect 599762 170960 599768 170972
rect 599820 170960 599826 171012
rect 675202 170960 675208 171012
rect 675260 170960 675266 171012
rect 673546 170008 673552 170060
rect 673604 170048 673610 170060
rect 675938 170048 675944 170060
rect 673604 170020 675944 170048
rect 673604 170008 673610 170020
rect 675938 170008 675944 170020
rect 675996 170008 676002 170060
rect 674650 169600 674656 169652
rect 674708 169640 674714 169652
rect 676030 169640 676036 169652
rect 674708 169612 676036 169640
rect 674708 169600 674714 169612
rect 676030 169600 676036 169612
rect 676088 169600 676094 169652
rect 673730 169192 673736 169244
rect 673788 169232 673794 169244
rect 675938 169232 675944 169244
rect 673788 169204 675944 169232
rect 673788 169192 673794 169204
rect 675938 169192 675944 169204
rect 675996 169192 676002 169244
rect 674006 168716 674012 168768
rect 674064 168756 674070 168768
rect 675938 168756 675944 168768
rect 674064 168728 675944 168756
rect 674064 168716 674070 168728
rect 675938 168716 675944 168728
rect 675996 168716 676002 168768
rect 674742 168648 674748 168700
rect 674800 168688 674806 168700
rect 676030 168688 676036 168700
rect 674800 168660 676036 168688
rect 674800 168648 674806 168660
rect 676030 168648 676036 168660
rect 676088 168648 676094 168700
rect 579706 168512 579712 168564
rect 579764 168552 579770 168564
rect 598934 168552 598940 168564
rect 579764 168524 598940 168552
rect 579764 168512 579770 168524
rect 598934 168512 598940 168524
rect 598992 168512 598998 168564
rect 673638 168512 673644 168564
rect 673696 168552 673702 168564
rect 675846 168552 675852 168564
rect 673696 168524 675852 168552
rect 673696 168512 673702 168524
rect 675846 168512 675852 168524
rect 675904 168512 675910 168564
rect 581914 168444 581920 168496
rect 581972 168484 581978 168496
rect 599946 168484 599952 168496
rect 581972 168456 599952 168484
rect 581972 168444 581978 168456
rect 599946 168444 599952 168456
rect 600004 168444 600010 168496
rect 580258 168376 580264 168428
rect 580316 168416 580322 168428
rect 599486 168416 599492 168428
rect 580316 168388 599492 168416
rect 580316 168376 580322 168388
rect 599486 168376 599492 168388
rect 599544 168376 599550 168428
rect 580166 168308 580172 168360
rect 580224 168348 580230 168360
rect 600222 168348 600228 168360
rect 580224 168320 600228 168348
rect 580224 168308 580230 168320
rect 600222 168308 600228 168320
rect 600280 168308 600286 168360
rect 672350 168240 672356 168292
rect 672408 168280 672414 168292
rect 676030 168280 676036 168292
rect 672408 168252 676036 168280
rect 672408 168240 672414 168252
rect 676030 168240 676036 168252
rect 676088 168240 676094 168292
rect 672166 167832 672172 167884
rect 672224 167872 672230 167884
rect 676030 167872 676036 167884
rect 672224 167844 676036 167872
rect 672224 167832 672230 167844
rect 676030 167832 676036 167844
rect 676088 167832 676094 167884
rect 672074 167424 672080 167476
rect 672132 167464 672138 167476
rect 676030 167464 676036 167476
rect 672132 167436 676036 167464
rect 672132 167424 672138 167436
rect 676030 167424 676036 167436
rect 676088 167424 676094 167476
rect 582282 165724 582288 165776
rect 582340 165764 582346 165776
rect 599854 165764 599860 165776
rect 582340 165736 599860 165764
rect 582340 165724 582346 165736
rect 599854 165724 599860 165736
rect 599912 165724 599918 165776
rect 580074 165656 580080 165708
rect 580132 165696 580138 165708
rect 600038 165696 600044 165708
rect 580132 165668 600044 165696
rect 580132 165656 580138 165668
rect 600038 165656 600044 165668
rect 600096 165656 600102 165708
rect 581546 165588 581552 165640
rect 581604 165628 581610 165640
rect 599946 165628 599952 165640
rect 581604 165600 599952 165628
rect 581604 165588 581610 165600
rect 599946 165588 599952 165600
rect 600004 165588 600010 165640
rect 581822 165520 581828 165572
rect 581880 165560 581886 165572
rect 601418 165560 601424 165572
rect 581880 165532 601424 165560
rect 581880 165520 581886 165532
rect 601418 165520 601424 165532
rect 601476 165520 601482 165572
rect 581638 162936 581644 162988
rect 581696 162976 581702 162988
rect 599854 162976 599860 162988
rect 581696 162948 599860 162976
rect 581696 162936 581702 162948
rect 599854 162936 599860 162948
rect 599912 162936 599918 162988
rect 581086 162868 581092 162920
rect 581144 162908 581150 162920
rect 599946 162908 599952 162920
rect 581144 162880 599952 162908
rect 581144 162868 581150 162880
rect 599946 162868 599952 162880
rect 600004 162868 600010 162920
rect 675754 160964 675760 161016
rect 675812 160964 675818 161016
rect 675772 160812 675800 160964
rect 675754 160760 675760 160812
rect 675812 160760 675818 160812
rect 582006 160216 582012 160268
rect 582064 160256 582070 160268
rect 599946 160256 599952 160268
rect 582064 160228 599952 160256
rect 582064 160216 582070 160228
rect 599946 160216 599952 160228
rect 600004 160216 600010 160268
rect 581730 160148 581736 160200
rect 581788 160188 581794 160200
rect 600038 160188 600044 160200
rect 581788 160160 600044 160188
rect 581788 160148 581794 160160
rect 600038 160148 600044 160160
rect 600096 160148 600102 160200
rect 581178 160080 581184 160132
rect 581236 160120 581242 160132
rect 599854 160120 599860 160132
rect 581236 160092 599860 160120
rect 581236 160080 581242 160092
rect 599854 160080 599860 160092
rect 599912 160080 599918 160132
rect 675202 160012 675208 160064
rect 675260 160052 675266 160064
rect 675386 160052 675392 160064
rect 675260 160024 675392 160052
rect 675260 160012 675266 160024
rect 675386 160012 675392 160024
rect 675444 160012 675450 160064
rect 674098 159332 674104 159384
rect 674156 159372 674162 159384
rect 675478 159372 675484 159384
rect 674156 159344 675484 159372
rect 674156 159332 674162 159344
rect 675478 159332 675484 159344
rect 675536 159332 675542 159384
rect 674834 157700 674840 157752
rect 674892 157740 674898 157752
rect 675478 157740 675484 157752
rect 674892 157712 675484 157740
rect 674892 157700 674898 157712
rect 675478 157700 675484 157712
rect 675536 157700 675542 157752
rect 580902 157496 580908 157548
rect 580960 157536 580966 157548
rect 599946 157536 599952 157548
rect 580960 157508 599952 157536
rect 580960 157496 580966 157508
rect 599946 157496 599952 157508
rect 600004 157496 600010 157548
rect 580994 157428 581000 157480
rect 581052 157468 581058 157480
rect 600038 157468 600044 157480
rect 581052 157440 600044 157468
rect 581052 157428 581058 157440
rect 600038 157428 600044 157440
rect 600096 157428 600102 157480
rect 580718 157360 580724 157412
rect 580776 157400 580782 157412
rect 599854 157400 599860 157412
rect 580776 157372 599860 157400
rect 580776 157360 580782 157372
rect 599854 157360 599860 157372
rect 599912 157360 599918 157412
rect 674558 156884 674564 156936
rect 674616 156924 674622 156936
rect 675386 156924 675392 156936
rect 674616 156896 675392 156924
rect 674616 156884 674622 156896
rect 675386 156884 675392 156896
rect 675444 156884 675450 156936
rect 674650 156476 674656 156528
rect 674708 156516 674714 156528
rect 675386 156516 675392 156528
rect 674708 156488 675392 156516
rect 674708 156476 674714 156488
rect 675386 156476 675392 156488
rect 675444 156476 675450 156528
rect 674742 155864 674748 155916
rect 674800 155904 674806 155916
rect 675478 155904 675484 155916
rect 674800 155876 675484 155904
rect 674800 155864 674806 155876
rect 675478 155864 675484 155876
rect 675536 155864 675542 155916
rect 582098 154640 582104 154692
rect 582156 154680 582162 154692
rect 599946 154680 599952 154692
rect 582156 154652 599952 154680
rect 582156 154640 582162 154652
rect 599946 154640 599952 154652
rect 600004 154640 600010 154692
rect 580626 154572 580632 154624
rect 580684 154612 580690 154624
rect 599854 154612 599860 154624
rect 580684 154584 599860 154612
rect 580684 154572 580690 154584
rect 599854 154572 599860 154584
rect 599912 154572 599918 154624
rect 673454 153348 673460 153400
rect 673512 153388 673518 153400
rect 675386 153388 675392 153400
rect 673512 153360 675392 153388
rect 673512 153348 673518 153360
rect 675386 153348 675392 153360
rect 675444 153348 675450 153400
rect 674006 152736 674012 152788
rect 674064 152776 674070 152788
rect 675386 152776 675392 152788
rect 674064 152748 675392 152776
rect 674064 152736 674070 152748
rect 675386 152736 675392 152748
rect 675444 152736 675450 152788
rect 673730 151988 673736 152040
rect 673788 152028 673794 152040
rect 675386 152028 675392 152040
rect 673788 152000 675392 152028
rect 673788 151988 673794 152000
rect 675386 151988 675392 152000
rect 675444 151988 675450 152040
rect 582190 151920 582196 151972
rect 582248 151960 582254 151972
rect 599854 151960 599860 151972
rect 582248 151932 599860 151960
rect 582248 151920 582254 151932
rect 599854 151920 599860 151932
rect 599912 151920 599918 151972
rect 581914 151852 581920 151904
rect 581972 151892 581978 151904
rect 599946 151892 599952 151904
rect 581972 151864 599952 151892
rect 581972 151852 581978 151864
rect 599946 151852 599952 151864
rect 600004 151852 600010 151904
rect 580810 151784 580816 151836
rect 580868 151824 580874 151836
rect 600038 151824 600044 151836
rect 580868 151796 600044 151824
rect 580868 151784 580874 151796
rect 600038 151784 600044 151796
rect 600096 151784 600102 151836
rect 673638 151376 673644 151428
rect 673696 151416 673702 151428
rect 675386 151416 675392 151428
rect 673696 151388 675392 151416
rect 673696 151376 673702 151388
rect 675386 151376 675392 151388
rect 675444 151376 675450 151428
rect 673546 150356 673552 150408
rect 673604 150396 673610 150408
rect 675386 150396 675392 150408
rect 673604 150368 675392 150396
rect 673604 150356 673610 150368
rect 675386 150356 675392 150368
rect 675444 150356 675450 150408
rect 581822 149200 581828 149252
rect 581880 149240 581886 149252
rect 598934 149240 598940 149252
rect 581880 149212 598940 149240
rect 581880 149200 581886 149212
rect 598934 149200 598940 149212
rect 598992 149200 598998 149252
rect 581454 149132 581460 149184
rect 581512 149172 581518 149184
rect 599854 149172 599860 149184
rect 581512 149144 599860 149172
rect 581512 149132 581518 149144
rect 599854 149132 599860 149144
rect 599912 149132 599918 149184
rect 581638 149064 581644 149116
rect 581696 149104 581702 149116
rect 599946 149104 599952 149116
rect 581696 149076 599952 149104
rect 581696 149064 581702 149076
rect 599946 149064 599952 149076
rect 600004 149064 600010 149116
rect 582282 146344 582288 146396
rect 582340 146384 582346 146396
rect 599854 146384 599860 146396
rect 582340 146356 599860 146384
rect 582340 146344 582346 146356
rect 599854 146344 599860 146356
rect 599912 146344 599918 146396
rect 581270 146276 581276 146328
rect 581328 146316 581334 146328
rect 599946 146316 599952 146328
rect 581328 146288 599952 146316
rect 581328 146276 581334 146288
rect 599946 146276 599952 146288
rect 600004 146276 600010 146328
rect 581730 143692 581736 143744
rect 581788 143732 581794 143744
rect 599946 143732 599952 143744
rect 581788 143704 599952 143732
rect 581788 143692 581794 143704
rect 599946 143692 599952 143704
rect 600004 143692 600010 143744
rect 579706 143624 579712 143676
rect 579764 143664 579770 143676
rect 599578 143664 599584 143676
rect 579764 143636 599584 143664
rect 579764 143624 579770 143636
rect 599578 143624 599584 143636
rect 599636 143624 599642 143676
rect 579798 143556 579804 143608
rect 579856 143596 579862 143608
rect 599670 143596 599676 143608
rect 579856 143568 599676 143596
rect 579856 143556 579862 143568
rect 599670 143556 599676 143568
rect 599728 143556 599734 143608
rect 581546 140904 581552 140956
rect 581604 140944 581610 140956
rect 599854 140944 599860 140956
rect 581604 140916 599860 140944
rect 581604 140904 581610 140916
rect 599854 140904 599860 140916
rect 599912 140904 599918 140956
rect 581362 140836 581368 140888
rect 581420 140876 581426 140888
rect 599946 140876 599952 140888
rect 581420 140848 599952 140876
rect 581420 140836 581426 140848
rect 599946 140836 599952 140848
rect 600004 140836 600010 140888
rect 581178 140768 581184 140820
rect 581236 140808 581242 140820
rect 599302 140808 599308 140820
rect 581236 140780 599308 140808
rect 581236 140768 581242 140780
rect 599302 140768 599308 140780
rect 599360 140768 599366 140820
rect 581086 138116 581092 138168
rect 581144 138156 581150 138168
rect 599946 138156 599952 138168
rect 581144 138128 599952 138156
rect 581144 138116 581150 138128
rect 599946 138116 599952 138128
rect 600004 138116 600010 138168
rect 580994 138048 581000 138100
rect 581052 138088 581058 138100
rect 599854 138088 599860 138100
rect 581052 138060 599860 138088
rect 581052 138048 581058 138060
rect 599854 138048 599860 138060
rect 599912 138048 599918 138100
rect 579890 137980 579896 138032
rect 579948 138020 579954 138032
rect 600038 138020 600044 138032
rect 579948 137992 600044 138020
rect 579948 137980 579954 137992
rect 600038 137980 600044 137992
rect 600096 137980 600102 138032
rect 580074 135328 580080 135380
rect 580132 135368 580138 135380
rect 599854 135368 599860 135380
rect 580132 135340 599860 135368
rect 580132 135328 580138 135340
rect 599854 135328 599860 135340
rect 599912 135328 599918 135380
rect 580166 135260 580172 135312
rect 580224 135300 580230 135312
rect 599946 135300 599952 135312
rect 580224 135272 599952 135300
rect 580224 135260 580230 135272
rect 599946 135260 599952 135272
rect 600004 135260 600010 135312
rect 704366 134308 704372 134360
rect 704424 134348 704430 134360
rect 704424 134320 708552 134348
rect 704424 134308 704430 134320
rect 704458 134240 704464 134292
rect 704516 134280 704522 134292
rect 708414 134280 708420 134292
rect 704516 134252 708420 134280
rect 704516 134240 704522 134252
rect 708414 134240 708420 134252
rect 708472 134240 708478 134292
rect 708524 134224 708552 134320
rect 707494 134212 707500 134224
rect 705304 134184 707500 134212
rect 705304 134088 705332 134184
rect 707494 134172 707500 134184
rect 707552 134172 707558 134224
rect 708506 134172 708512 134224
rect 708564 134172 708570 134224
rect 707034 134144 707040 134156
rect 705764 134116 707040 134144
rect 705764 134088 705792 134116
rect 707034 134104 707040 134116
rect 707092 134104 707098 134156
rect 705286 134036 705292 134088
rect 705344 134036 705350 134088
rect 705746 134036 705752 134088
rect 705804 134036 705810 134088
rect 706206 134036 706212 134088
rect 706264 134076 706270 134088
rect 706574 134076 706580 134088
rect 706264 134048 706580 134076
rect 706264 134036 706270 134048
rect 706574 134036 706580 134048
rect 706632 134036 706638 134088
rect 705838 133968 705844 134020
rect 705896 134008 705902 134020
rect 707034 134008 707040 134020
rect 705896 133980 707040 134008
rect 705896 133968 705902 133980
rect 707034 133968 707040 133980
rect 707092 133968 707098 134020
rect 706298 133900 706304 133952
rect 706356 133940 706362 133952
rect 706574 133940 706580 133952
rect 706356 133912 706580 133940
rect 706356 133900 706362 133912
rect 706574 133900 706580 133912
rect 706632 133900 706638 133952
rect 704826 133832 704832 133884
rect 704884 133832 704890 133884
rect 705378 133832 705384 133884
rect 705436 133872 705442 133884
rect 707494 133872 707500 133884
rect 705436 133844 707500 133872
rect 705436 133832 705442 133844
rect 707494 133832 707500 133844
rect 707552 133832 707558 133884
rect 704844 133736 704872 133832
rect 704918 133764 704924 133816
rect 704976 133804 704982 133816
rect 707954 133804 707960 133816
rect 704976 133776 707960 133804
rect 704976 133764 704982 133776
rect 707954 133764 707960 133776
rect 708012 133764 708018 133816
rect 708046 133736 708052 133748
rect 704844 133708 708052 133736
rect 708046 133696 708052 133708
rect 708104 133696 708110 133748
rect 703998 133628 704004 133680
rect 704056 133668 704062 133680
rect 708874 133668 708880 133680
rect 704056 133640 708880 133668
rect 704056 133628 704062 133640
rect 708874 133628 708880 133640
rect 708932 133628 708938 133680
rect 670050 132880 670056 132932
rect 670108 132920 670114 132932
rect 676214 132920 676220 132932
rect 670108 132892 676220 132920
rect 670108 132880 670114 132892
rect 676214 132880 676220 132892
rect 676272 132880 676278 132932
rect 669498 132744 669504 132796
rect 669556 132784 669562 132796
rect 676122 132784 676128 132796
rect 669556 132756 676128 132784
rect 669556 132744 669562 132756
rect 676122 132744 676128 132756
rect 676180 132744 676186 132796
rect 580902 132608 580908 132660
rect 580960 132648 580966 132660
rect 599302 132648 599308 132660
rect 580960 132620 599308 132648
rect 580960 132608 580966 132620
rect 599302 132608 599308 132620
rect 599360 132608 599366 132660
rect 669314 132608 669320 132660
rect 669372 132648 669378 132660
rect 676030 132648 676036 132660
rect 669372 132620 676036 132648
rect 669372 132608 669378 132620
rect 676030 132608 676036 132620
rect 676088 132608 676094 132660
rect 580258 132540 580264 132592
rect 580316 132580 580322 132592
rect 599946 132580 599952 132592
rect 580316 132552 599952 132580
rect 580316 132540 580322 132552
rect 599946 132540 599952 132552
rect 600004 132540 600010 132592
rect 579982 132472 579988 132524
rect 580040 132512 580046 132524
rect 599854 132512 599860 132524
rect 580040 132484 599860 132512
rect 580040 132472 580046 132484
rect 599854 132472 599860 132484
rect 599912 132472 599918 132524
rect 673270 132268 673276 132320
rect 673328 132308 673334 132320
rect 676214 132308 676220 132320
rect 673328 132280 676220 132308
rect 673328 132268 673334 132280
rect 676214 132268 676220 132280
rect 676272 132268 676278 132320
rect 670786 131656 670792 131708
rect 670844 131696 670850 131708
rect 676030 131696 676036 131708
rect 670844 131668 676036 131696
rect 670844 131656 670850 131668
rect 676030 131656 676036 131668
rect 676088 131656 676094 131708
rect 673362 131452 673368 131504
rect 673420 131492 673426 131504
rect 676214 131492 676220 131504
rect 673420 131464 676220 131492
rect 673420 131452 673426 131464
rect 676214 131452 676220 131464
rect 676272 131452 676278 131504
rect 672442 130840 672448 130892
rect 672500 130880 672506 130892
rect 676030 130880 676036 130892
rect 672500 130852 676036 130880
rect 672500 130840 672506 130852
rect 676030 130840 676036 130852
rect 676088 130840 676094 130892
rect 672258 130636 672264 130688
rect 672316 130676 672322 130688
rect 676214 130676 676220 130688
rect 672316 130648 676220 130676
rect 672316 130636 672322 130648
rect 676214 130636 676220 130648
rect 676272 130636 676278 130688
rect 670878 130024 670884 130076
rect 670936 130064 670942 130076
rect 676030 130064 676036 130076
rect 670936 130036 676036 130064
rect 670936 130024 670942 130036
rect 676030 130024 676036 130036
rect 676088 130024 676094 130076
rect 580534 129888 580540 129940
rect 580592 129928 580598 129940
rect 599854 129928 599860 129940
rect 580592 129900 599860 129928
rect 580592 129888 580598 129900
rect 599854 129888 599860 129900
rect 599912 129888 599918 129940
rect 580350 129820 580356 129872
rect 580408 129860 580414 129872
rect 599946 129860 599952 129872
rect 580408 129832 599952 129860
rect 580408 129820 580414 129832
rect 599946 129820 599952 129832
rect 600004 129820 600010 129872
rect 669222 129820 669228 129872
rect 669280 129860 669286 129872
rect 670786 129860 670792 129872
rect 669280 129832 670792 129860
rect 669280 129820 669286 129832
rect 670786 129820 670792 129832
rect 670844 129820 670850 129872
rect 580442 129752 580448 129804
rect 580500 129792 580506 129804
rect 598934 129792 598940 129804
rect 580500 129764 598940 129792
rect 580500 129752 580506 129764
rect 598934 129752 598940 129764
rect 598992 129752 598998 129804
rect 666738 129752 666744 129804
rect 666796 129792 666802 129804
rect 670878 129792 670884 129804
rect 666796 129764 670884 129792
rect 666796 129752 666802 129764
rect 670878 129752 670884 129764
rect 670936 129752 670942 129804
rect 671890 129684 671896 129736
rect 671948 129724 671954 129736
rect 676030 129724 676036 129736
rect 671948 129696 676036 129724
rect 671948 129684 671954 129696
rect 676030 129684 676036 129696
rect 676088 129684 676094 129736
rect 671982 129412 671988 129464
rect 672040 129452 672046 129464
rect 676214 129452 676220 129464
rect 672040 129424 676220 129452
rect 672040 129412 672046 129424
rect 676214 129412 676220 129424
rect 676272 129412 676278 129464
rect 674466 127712 674472 127764
rect 674524 127752 674530 127764
rect 676030 127752 676036 127764
rect 674524 127724 676036 127752
rect 674524 127712 674530 127724
rect 676030 127712 676036 127724
rect 676088 127712 676094 127764
rect 582190 127032 582196 127084
rect 582248 127072 582254 127084
rect 599946 127072 599952 127084
rect 582248 127044 599952 127072
rect 582248 127032 582254 127044
rect 599946 127032 599952 127044
rect 600004 127032 600010 127084
rect 673638 127032 673644 127084
rect 673696 127072 673702 127084
rect 675938 127072 675944 127084
rect 673696 127044 675944 127072
rect 673696 127032 673702 127044
rect 675938 127032 675944 127044
rect 675996 127032 676002 127084
rect 580718 126964 580724 127016
rect 580776 127004 580782 127016
rect 599854 127004 599860 127016
rect 580776 126976 599860 127004
rect 580776 126964 580782 126976
rect 599854 126964 599860 126976
rect 599912 126964 599918 127016
rect 674558 126964 674564 127016
rect 674616 127004 674622 127016
rect 676030 127004 676036 127016
rect 674616 126976 676036 127004
rect 674616 126964 674622 126976
rect 676030 126964 676036 126976
rect 676088 126964 676094 127016
rect 673454 124856 673460 124908
rect 673512 124896 673518 124908
rect 675846 124896 675852 124908
rect 673512 124868 675852 124896
rect 673512 124856 673518 124868
rect 675846 124856 675852 124868
rect 675904 124856 675910 124908
rect 674742 124448 674748 124500
rect 674800 124488 674806 124500
rect 675938 124488 675944 124500
rect 674800 124460 675944 124488
rect 674800 124448 674806 124460
rect 675938 124448 675944 124460
rect 675996 124448 676002 124500
rect 673546 124380 673552 124432
rect 673604 124420 673610 124432
rect 675846 124420 675852 124432
rect 673604 124392 675852 124420
rect 673604 124380 673610 124392
rect 675846 124380 675852 124392
rect 675904 124380 675910 124432
rect 582006 124312 582012 124364
rect 582064 124352 582070 124364
rect 599946 124352 599952 124364
rect 582064 124324 599952 124352
rect 582064 124312 582070 124324
rect 599946 124312 599952 124324
rect 600004 124312 600010 124364
rect 674650 124312 674656 124364
rect 674708 124352 674714 124364
rect 676122 124352 676128 124364
rect 674708 124324 676128 124352
rect 674708 124312 674714 124324
rect 676122 124312 676128 124324
rect 676180 124312 676186 124364
rect 580810 124244 580816 124296
rect 580868 124284 580874 124296
rect 600038 124284 600044 124296
rect 580868 124256 600044 124284
rect 580868 124244 580874 124256
rect 600038 124244 600044 124256
rect 600096 124244 600102 124296
rect 675110 124244 675116 124296
rect 675168 124284 675174 124296
rect 675938 124284 675944 124296
rect 675168 124256 675944 124284
rect 675168 124244 675174 124256
rect 675938 124244 675944 124256
rect 675996 124244 676002 124296
rect 580626 124176 580632 124228
rect 580684 124216 580690 124228
rect 599854 124216 599860 124228
rect 580684 124188 599860 124216
rect 580684 124176 580690 124188
rect 599854 124176 599860 124188
rect 599912 124176 599918 124228
rect 675202 124176 675208 124228
rect 675260 124216 675266 124228
rect 676030 124216 676036 124228
rect 675260 124188 676036 124216
rect 675260 124176 675266 124188
rect 676030 124176 676036 124188
rect 676088 124176 676094 124228
rect 673822 123224 673828 123276
rect 673880 123264 673886 123276
rect 676030 123264 676036 123276
rect 673880 123236 676036 123264
rect 673880 123224 673886 123236
rect 676030 123224 676036 123236
rect 676088 123224 676094 123276
rect 671430 123088 671436 123140
rect 671488 123128 671494 123140
rect 676030 123128 676036 123140
rect 671488 123100 676036 123128
rect 671488 123088 671494 123100
rect 676030 123088 676036 123100
rect 676088 123088 676094 123140
rect 672902 122680 672908 122732
rect 672960 122720 672966 122732
rect 676030 122720 676036 122732
rect 672960 122692 676036 122720
rect 672960 122680 672966 122692
rect 676030 122680 676036 122692
rect 676088 122680 676094 122732
rect 672258 122272 672264 122324
rect 672316 122312 672322 122324
rect 676030 122312 676036 122324
rect 672316 122284 676036 122312
rect 672316 122272 672322 122284
rect 676030 122272 676036 122284
rect 676088 122272 676094 122324
rect 582282 121592 582288 121644
rect 582340 121632 582346 121644
rect 598934 121632 598940 121644
rect 582340 121604 598940 121632
rect 582340 121592 582346 121604
rect 598934 121592 598940 121604
rect 598992 121592 598998 121644
rect 582098 121524 582104 121576
rect 582156 121564 582162 121576
rect 599854 121564 599860 121576
rect 582156 121536 599860 121564
rect 582156 121524 582162 121536
rect 599854 121524 599860 121536
rect 599912 121524 599918 121576
rect 581914 121456 581920 121508
rect 581972 121496 581978 121508
rect 599946 121496 599952 121508
rect 581972 121468 599952 121496
rect 581972 121456 581978 121468
rect 599946 121456 599952 121468
rect 600004 121456 600010 121508
rect 673730 121456 673736 121508
rect 673788 121496 673794 121508
rect 675938 121496 675944 121508
rect 673788 121468 675944 121496
rect 673788 121456 673794 121468
rect 675938 121456 675944 121468
rect 675996 121456 676002 121508
rect 583662 118804 583668 118856
rect 583720 118844 583726 118856
rect 599854 118844 599860 118856
rect 583720 118816 599860 118844
rect 583720 118804 583726 118816
rect 599854 118804 599860 118816
rect 599912 118804 599918 118856
rect 581638 118736 581644 118788
rect 581696 118776 581702 118788
rect 599946 118776 599952 118788
rect 581696 118748 599952 118776
rect 581696 118736 581702 118748
rect 599946 118736 599952 118748
rect 600004 118736 600010 118788
rect 581822 118668 581828 118720
rect 581880 118708 581886 118720
rect 600038 118708 600044 118720
rect 581880 118680 600044 118708
rect 581880 118668 581886 118680
rect 600038 118668 600044 118680
rect 600096 118668 600102 118720
rect 581730 116016 581736 116068
rect 581788 116056 581794 116068
rect 599854 116056 599860 116068
rect 581788 116028 599860 116056
rect 581788 116016 581794 116028
rect 599854 116016 599860 116028
rect 599912 116016 599918 116068
rect 581270 115948 581276 116000
rect 581328 115988 581334 116000
rect 599946 115988 599952 116000
rect 581328 115960 599952 115988
rect 581328 115948 581334 115960
rect 599946 115948 599952 115960
rect 600004 115948 600010 116000
rect 675754 115744 675760 115796
rect 675812 115744 675818 115796
rect 675772 115592 675800 115744
rect 675754 115540 675760 115592
rect 675812 115540 675818 115592
rect 675202 114996 675208 115048
rect 675260 115036 675266 115048
rect 675386 115036 675392 115048
rect 675260 115008 675392 115036
rect 675260 114996 675266 115008
rect 675386 114996 675392 115008
rect 675444 114996 675450 115048
rect 674466 114180 674472 114232
rect 674524 114220 674530 114232
rect 675386 114220 675392 114232
rect 674524 114192 675392 114220
rect 674524 114180 674530 114192
rect 675386 114180 675392 114192
rect 675444 114180 675450 114232
rect 581362 113228 581368 113280
rect 581420 113268 581426 113280
rect 599946 113268 599952 113280
rect 581420 113240 599952 113268
rect 581420 113228 581426 113240
rect 599946 113228 599952 113240
rect 600004 113228 600010 113280
rect 581546 113160 581552 113212
rect 581604 113200 581610 113212
rect 599854 113200 599860 113212
rect 581604 113172 599860 113200
rect 581604 113160 581610 113172
rect 599854 113160 599860 113172
rect 599912 113160 599918 113212
rect 674558 112344 674564 112396
rect 674616 112384 674622 112396
rect 675386 112384 675392 112396
rect 674616 112356 675392 112384
rect 674616 112344 674622 112356
rect 675386 112344 675392 112356
rect 675444 112344 675450 112396
rect 674742 111868 674748 111920
rect 674800 111908 674806 111920
rect 675386 111908 675392 111920
rect 674800 111880 675392 111908
rect 674800 111868 674806 111880
rect 675386 111868 675392 111880
rect 675444 111868 675450 111920
rect 674650 111120 674656 111172
rect 674708 111160 674714 111172
rect 675386 111160 675392 111172
rect 674708 111132 675392 111160
rect 674708 111120 674714 111132
rect 675386 111120 675392 111132
rect 675444 111120 675450 111172
rect 675110 110644 675116 110696
rect 675168 110684 675174 110696
rect 675386 110684 675392 110696
rect 675168 110656 675392 110684
rect 675168 110644 675174 110656
rect 675386 110644 675392 110656
rect 675444 110644 675450 110696
rect 581454 110508 581460 110560
rect 581512 110548 581518 110560
rect 599946 110548 599952 110560
rect 581512 110520 599952 110548
rect 581512 110508 581518 110520
rect 599946 110508 599952 110520
rect 600004 110508 600010 110560
rect 581178 110440 581184 110492
rect 581236 110480 581242 110492
rect 599762 110480 599768 110492
rect 581236 110452 599768 110480
rect 581236 110440 581242 110452
rect 599762 110440 599768 110452
rect 599820 110440 599826 110492
rect 673638 108196 673644 108248
rect 673696 108236 673702 108248
rect 675478 108236 675484 108248
rect 673696 108208 675484 108236
rect 673696 108196 673702 108208
rect 675478 108196 675484 108208
rect 675536 108196 675542 108248
rect 580994 107652 581000 107704
rect 581052 107692 581058 107704
rect 599946 107692 599952 107704
rect 581052 107664 599952 107692
rect 581052 107652 581058 107664
rect 599946 107652 599952 107664
rect 600004 107652 600010 107704
rect 673822 107516 673828 107568
rect 673880 107556 673886 107568
rect 675386 107556 675392 107568
rect 673880 107528 675392 107556
rect 673880 107516 673886 107528
rect 675386 107516 675392 107528
rect 675444 107516 675450 107568
rect 673546 106972 673552 107024
rect 673604 107012 673610 107024
rect 675386 107012 675392 107024
rect 673604 106984 675392 107012
rect 673604 106972 673610 106984
rect 675386 106972 675392 106984
rect 675444 106972 675450 107024
rect 673730 106360 673736 106412
rect 673788 106400 673794 106412
rect 675386 106400 675392 106412
rect 673788 106372 675392 106400
rect 673788 106360 673794 106372
rect 675386 106360 675392 106372
rect 675444 106360 675450 106412
rect 673454 105136 673460 105188
rect 673512 105176 673518 105188
rect 675478 105176 675484 105188
rect 673512 105148 675484 105176
rect 673512 105136 673518 105148
rect 675478 105136 675484 105148
rect 675536 105136 675542 105188
rect 581086 104864 581092 104916
rect 581144 104904 581150 104916
rect 599946 104904 599952 104916
rect 581144 104876 599952 104904
rect 581144 104864 581150 104876
rect 599946 104864 599952 104876
rect 600004 104864 600010 104916
rect 657722 99764 657728 99816
rect 657780 99804 657786 99816
rect 660896 99804 660902 99816
rect 657780 99776 660902 99804
rect 657780 99764 657786 99776
rect 660896 99764 660902 99776
rect 660954 99764 660960 99816
rect 580902 99356 580908 99408
rect 580960 99396 580966 99408
rect 599946 99396 599952 99408
rect 580960 99368 599952 99396
rect 580960 99356 580966 99368
rect 599946 99356 599952 99368
rect 600004 99356 600010 99408
rect 633066 96568 633072 96620
rect 633124 96608 633130 96620
rect 635274 96608 635280 96620
rect 633124 96580 635280 96608
rect 633124 96568 633130 96580
rect 635274 96568 635280 96580
rect 635332 96568 635338 96620
rect 636286 96568 636292 96620
rect 636344 96608 636350 96620
rect 640978 96608 640984 96620
rect 636344 96580 640984 96608
rect 636344 96568 636350 96580
rect 640978 96568 640984 96580
rect 641036 96568 641042 96620
rect 655974 96568 655980 96620
rect 656032 96608 656038 96620
rect 659562 96608 659568 96620
rect 656032 96580 659568 96608
rect 656032 96568 656038 96580
rect 659562 96568 659568 96580
rect 659620 96568 659626 96620
rect 661862 96568 661868 96620
rect 661920 96608 661926 96620
rect 663058 96608 663064 96620
rect 661920 96580 663064 96608
rect 661920 96568 661926 96580
rect 663058 96568 663064 96580
rect 663116 96568 663122 96620
rect 633802 96500 633808 96552
rect 633860 96540 633866 96552
rect 636378 96540 636384 96552
rect 633860 96512 636384 96540
rect 633860 96500 633866 96512
rect 636378 96500 636384 96512
rect 636436 96500 636442 96552
rect 637022 96500 637028 96552
rect 637080 96540 637086 96552
rect 642358 96540 642364 96552
rect 637080 96512 642364 96540
rect 637080 96500 637086 96512
rect 642358 96500 642364 96512
rect 642416 96500 642422 96552
rect 654686 96500 654692 96552
rect 654744 96540 654750 96552
rect 658274 96540 658280 96552
rect 654744 96512 658280 96540
rect 654744 96500 654750 96512
rect 658274 96500 658280 96512
rect 658332 96500 658338 96552
rect 659102 96500 659108 96552
rect 659160 96540 659166 96552
rect 662506 96540 662512 96552
rect 659160 96512 662512 96540
rect 659160 96500 659166 96512
rect 662506 96500 662512 96512
rect 662564 96500 662570 96552
rect 634446 96432 634452 96484
rect 634504 96472 634510 96484
rect 637574 96472 637580 96484
rect 634504 96444 637580 96472
rect 634504 96432 634510 96444
rect 637574 96432 637580 96444
rect 637632 96432 637638 96484
rect 652018 96432 652024 96484
rect 652076 96472 652082 96484
rect 661954 96472 661960 96484
rect 652076 96444 661960 96472
rect 652076 96432 652082 96444
rect 661954 96432 661960 96444
rect 662012 96432 662018 96484
rect 635734 96364 635740 96416
rect 635792 96404 635798 96416
rect 639874 96404 639880 96416
rect 635792 96376 639880 96404
rect 635792 96364 635798 96376
rect 639874 96364 639880 96376
rect 639932 96364 639938 96416
rect 631134 96024 631140 96076
rect 631192 96064 631198 96076
rect 632100 96064 632106 96076
rect 631192 96036 632106 96064
rect 631192 96024 631198 96036
rect 632100 96024 632106 96036
rect 632158 96024 632164 96076
rect 632422 96024 632428 96076
rect 632480 96064 632486 96076
rect 634400 96064 634406 96076
rect 632480 96036 634406 96064
rect 632480 96024 632486 96036
rect 634400 96024 634406 96036
rect 634458 96024 634464 96076
rect 635090 96024 635096 96076
rect 635148 96064 635154 96076
rect 639000 96064 639006 96076
rect 635148 96036 639006 96064
rect 635148 96024 635154 96036
rect 639000 96024 639006 96036
rect 639058 96024 639064 96076
rect 647510 96024 647516 96076
rect 647568 96064 647574 96076
rect 653214 96064 653220 96076
rect 647568 96036 653220 96064
rect 647568 96024 647574 96036
rect 653214 96024 653220 96036
rect 653272 96024 653278 96076
rect 631778 95888 631784 95940
rect 631836 95928 631842 95940
rect 632974 95928 632980 95940
rect 631836 95900 632980 95928
rect 631836 95888 631842 95900
rect 632974 95888 632980 95900
rect 633032 95888 633038 95940
rect 640058 95888 640064 95940
rect 640116 95928 640122 95940
rect 646038 95928 646044 95940
rect 640116 95900 646044 95928
rect 640116 95888 640122 95900
rect 646038 95888 646044 95900
rect 646096 95888 646102 95940
rect 638862 95820 638868 95872
rect 638920 95860 638926 95872
rect 646222 95860 646228 95872
rect 638920 95832 646228 95860
rect 638920 95820 638926 95832
rect 646222 95820 646228 95832
rect 646280 95820 646286 95872
rect 616782 95752 616788 95804
rect 616840 95792 616846 95804
rect 623222 95792 623228 95804
rect 616840 95764 623228 95792
rect 616840 95752 616846 95764
rect 623222 95752 623228 95764
rect 623280 95752 623286 95804
rect 639598 95752 639604 95804
rect 639656 95792 639662 95804
rect 645946 95792 645952 95804
rect 639656 95764 645952 95792
rect 639656 95752 639662 95764
rect 645946 95752 645952 95764
rect 646004 95752 646010 95804
rect 621198 95684 621204 95736
rect 621256 95724 621262 95736
rect 622026 95724 622032 95736
rect 621256 95696 622032 95724
rect 621256 95684 621262 95696
rect 622026 95684 622032 95696
rect 622084 95684 622090 95736
rect 637482 95684 637488 95736
rect 637540 95724 637546 95736
rect 640518 95724 640524 95736
rect 637540 95696 640524 95724
rect 637540 95684 637546 95696
rect 640518 95684 640524 95696
rect 640576 95684 640582 95736
rect 640886 95684 640892 95736
rect 640944 95724 640950 95736
rect 645854 95724 645860 95736
rect 640944 95696 645860 95724
rect 640944 95684 640950 95696
rect 645854 95684 645860 95696
rect 645912 95684 645918 95736
rect 603534 95616 603540 95668
rect 603592 95656 603598 95668
rect 610434 95656 610440 95668
rect 603592 95628 610440 95656
rect 603592 95616 603598 95628
rect 610434 95616 610440 95628
rect 610492 95616 610498 95668
rect 619358 95616 619364 95668
rect 619416 95656 619422 95668
rect 623406 95656 623412 95668
rect 619416 95628 623412 95656
rect 619416 95616 619422 95628
rect 623406 95616 623412 95628
rect 623464 95616 623470 95668
rect 641622 95616 641628 95668
rect 641680 95656 641686 95668
rect 642818 95656 642824 95668
rect 641680 95628 642824 95656
rect 641680 95616 641686 95628
rect 642818 95616 642824 95628
rect 642876 95616 642882 95668
rect 604454 95548 604460 95600
rect 604512 95588 604518 95600
rect 606386 95588 606392 95600
rect 604512 95560 606392 95588
rect 604512 95548 604518 95560
rect 606386 95548 606392 95560
rect 606444 95548 606450 95600
rect 607490 95548 607496 95600
rect 607548 95588 607554 95600
rect 608962 95588 608968 95600
rect 607548 95560 608968 95588
rect 607548 95548 607554 95560
rect 608962 95548 608968 95560
rect 609020 95548 609026 95600
rect 610250 95548 610256 95600
rect 610308 95588 610314 95600
rect 611538 95588 611544 95600
rect 610308 95560 611544 95588
rect 610308 95548 610314 95560
rect 611538 95548 611544 95560
rect 611596 95548 611602 95600
rect 612826 95548 612832 95600
rect 612884 95588 612890 95600
rect 613562 95588 613568 95600
rect 612884 95560 613568 95588
rect 612884 95548 612890 95560
rect 613562 95548 613568 95560
rect 613620 95548 613626 95600
rect 618254 95548 618260 95600
rect 618312 95588 618318 95600
rect 620094 95588 620100 95600
rect 618312 95560 620100 95588
rect 618312 95548 618318 95560
rect 620094 95548 620100 95560
rect 620152 95548 620158 95600
rect 621474 95548 621480 95600
rect 621532 95588 621538 95600
rect 623314 95588 623320 95600
rect 621532 95560 623320 95588
rect 621532 95548 621538 95560
rect 623314 95548 623320 95560
rect 623372 95548 623378 95600
rect 623774 95548 623780 95600
rect 623832 95588 623838 95600
rect 624602 95588 624608 95600
rect 623832 95560 624608 95588
rect 623832 95548 623838 95560
rect 624602 95548 624608 95560
rect 624660 95548 624666 95600
rect 638310 95548 638316 95600
rect 638368 95548 638374 95600
rect 642266 95548 642272 95600
rect 642324 95588 642330 95600
rect 642910 95588 642916 95600
rect 642324 95560 642916 95588
rect 642324 95548 642330 95560
rect 642910 95548 642916 95560
rect 642968 95548 642974 95600
rect 656986 95548 656992 95600
rect 657044 95588 657050 95600
rect 659194 95588 659200 95600
rect 657044 95560 659200 95588
rect 657044 95548 657050 95560
rect 659194 95548 659200 95560
rect 659252 95548 659258 95600
rect 610158 95480 610164 95532
rect 610216 95520 610222 95532
rect 612182 95520 612188 95532
rect 610216 95492 612188 95520
rect 610216 95480 610222 95492
rect 612182 95480 612188 95492
rect 612240 95480 612246 95532
rect 617426 95480 617432 95532
rect 617484 95520 617490 95532
rect 623130 95520 623136 95532
rect 617484 95492 623136 95520
rect 617484 95480 617490 95492
rect 623130 95480 623136 95492
rect 623188 95480 623194 95532
rect 638328 95520 638356 95548
rect 642726 95520 642732 95532
rect 638328 95492 642732 95520
rect 642726 95480 642732 95492
rect 642784 95480 642790 95532
rect 660574 95480 660580 95532
rect 660632 95520 660638 95532
rect 661402 95520 661408 95532
rect 660632 95492 661408 95520
rect 660632 95480 660638 95492
rect 661402 95480 661408 95492
rect 661460 95480 661466 95532
rect 620002 95412 620008 95464
rect 620060 95452 620066 95464
rect 622302 95452 622308 95464
rect 620060 95424 622308 95452
rect 620060 95412 620066 95424
rect 622302 95412 622308 95424
rect 622360 95412 622366 95464
rect 616138 95344 616144 95396
rect 616196 95384 616202 95396
rect 622486 95384 622492 95396
rect 616196 95356 622492 95384
rect 616196 95344 616202 95356
rect 622486 95344 622492 95356
rect 622544 95344 622550 95396
rect 656618 95344 656624 95396
rect 656676 95384 656682 95396
rect 663150 95384 663156 95396
rect 656676 95356 663156 95384
rect 656676 95344 656682 95356
rect 663150 95344 663156 95356
rect 663208 95344 663214 95396
rect 646774 95276 646780 95328
rect 646832 95316 646838 95328
rect 663334 95316 663340 95328
rect 646832 95288 663340 95316
rect 646832 95276 646838 95288
rect 663334 95276 663340 95288
rect 663392 95276 663398 95328
rect 589182 95208 589188 95260
rect 589240 95248 589246 95260
rect 610894 95248 610900 95260
rect 589240 95220 610900 95248
rect 589240 95208 589246 95220
rect 610894 95208 610900 95220
rect 610952 95208 610958 95260
rect 643554 95208 643560 95260
rect 643612 95248 643618 95260
rect 644842 95248 644848 95260
rect 643612 95220 644848 95248
rect 643612 95208 643618 95220
rect 644842 95208 644848 95220
rect 644900 95208 644906 95260
rect 651466 95208 651472 95260
rect 651524 95248 651530 95260
rect 653398 95248 653404 95260
rect 651524 95220 653404 95248
rect 651524 95208 651530 95220
rect 653398 95208 653404 95220
rect 653456 95208 653462 95260
rect 657078 95208 657084 95260
rect 657136 95248 657142 95260
rect 657906 95248 657912 95260
rect 657136 95220 657912 95248
rect 657136 95208 657142 95220
rect 657906 95208 657912 95220
rect 657964 95208 657970 95260
rect 646130 95140 646136 95192
rect 646188 95180 646194 95192
rect 663426 95180 663432 95192
rect 646188 95152 663432 95180
rect 646188 95140 646194 95152
rect 663426 95140 663432 95152
rect 663484 95140 663490 95192
rect 597462 95072 597468 95124
rect 597520 95112 597526 95124
rect 607674 95112 607680 95124
rect 597520 95084 607680 95112
rect 597520 95072 597526 95084
rect 607674 95072 607680 95084
rect 607732 95072 607738 95124
rect 646682 95072 646688 95124
rect 646740 95112 646746 95124
rect 648154 95112 648160 95124
rect 646740 95084 648160 95112
rect 646740 95072 646746 95084
rect 648154 95072 648160 95084
rect 648212 95072 648218 95124
rect 648890 95072 648896 95124
rect 648948 95112 648954 95124
rect 650730 95112 650736 95124
rect 648948 95084 650736 95112
rect 648948 95072 648954 95084
rect 650730 95072 650736 95084
rect 650788 95072 650794 95124
rect 652662 95072 652668 95124
rect 652720 95112 652726 95124
rect 663794 95112 663800 95124
rect 652720 95084 663800 95112
rect 652720 95072 652726 95084
rect 663794 95072 663800 95084
rect 663852 95072 663858 95124
rect 614850 94936 614856 94988
rect 614908 94976 614914 94988
rect 615402 94976 615408 94988
rect 614908 94948 615408 94976
rect 614908 94936 614914 94948
rect 615402 94936 615408 94948
rect 615460 94936 615466 94988
rect 648706 94800 648712 94852
rect 648764 94840 648770 94852
rect 650086 94840 650092 94852
rect 648764 94812 650092 94840
rect 648764 94800 648770 94812
rect 650086 94800 650092 94812
rect 650144 94800 650150 94852
rect 618714 94732 618720 94784
rect 618772 94772 618778 94784
rect 623314 94772 623320 94784
rect 618772 94744 623320 94772
rect 618772 94732 618778 94744
rect 623314 94732 623320 94744
rect 623372 94732 623378 94784
rect 645946 94732 645952 94784
rect 646004 94772 646010 94784
rect 646222 94772 646228 94784
rect 646004 94744 646228 94772
rect 646004 94732 646010 94744
rect 646222 94732 646228 94744
rect 646280 94732 646286 94784
rect 648798 94664 648804 94716
rect 648856 94704 648862 94716
rect 649442 94704 649448 94716
rect 648856 94676 649448 94704
rect 648856 94664 648862 94676
rect 649442 94664 649448 94676
rect 649500 94664 649506 94716
rect 653306 94664 653312 94716
rect 653364 94704 653370 94716
rect 663702 94704 663708 94716
rect 653364 94676 663708 94704
rect 653364 94664 653370 94676
rect 663702 94664 663708 94676
rect 663760 94664 663766 94716
rect 657262 94596 657268 94648
rect 657320 94636 657326 94648
rect 663518 94636 663524 94648
rect 657320 94608 663524 94636
rect 657320 94596 657326 94608
rect 663518 94596 663524 94608
rect 663576 94596 663582 94648
rect 618070 94528 618076 94580
rect 618128 94568 618134 94580
rect 621934 94568 621940 94580
rect 618128 94540 621940 94568
rect 618128 94528 618134 94540
rect 621934 94528 621940 94540
rect 621992 94528 621998 94580
rect 656894 94528 656900 94580
rect 656952 94568 656958 94580
rect 658550 94568 658556 94580
rect 656952 94540 658556 94568
rect 656952 94528 656958 94540
rect 658550 94528 658556 94540
rect 658608 94528 658614 94580
rect 648062 94460 648068 94512
rect 648120 94500 648126 94512
rect 659838 94500 659844 94512
rect 648120 94472 659844 94500
rect 648120 94460 648126 94472
rect 659838 94460 659844 94472
rect 659896 94460 659902 94512
rect 660390 94460 660396 94512
rect 660448 94460 660454 94512
rect 643462 94188 643468 94240
rect 643520 94228 643526 94240
rect 660408 94228 660436 94460
rect 643520 94200 660436 94228
rect 643520 94188 643526 94200
rect 644198 94052 644204 94104
rect 644256 94092 644262 94104
rect 654042 94092 654048 94104
rect 644256 94064 654048 94092
rect 644256 94052 644262 94064
rect 654042 94052 654048 94064
rect 654100 94052 654106 94104
rect 649350 93984 649356 94036
rect 649408 94024 649414 94036
rect 656894 94024 656900 94036
rect 649408 93996 656900 94024
rect 649408 93984 649414 93996
rect 656894 93984 656900 93996
rect 656952 93984 656958 94036
rect 644750 93848 644756 93900
rect 644808 93888 644814 93900
rect 653490 93888 653496 93900
rect 644808 93860 653496 93888
rect 644808 93848 644814 93860
rect 653490 93848 653496 93860
rect 653548 93848 653554 93900
rect 613010 91672 613016 91724
rect 613068 91712 613074 91724
rect 614942 91712 614948 91724
rect 613068 91684 614948 91712
rect 613068 91672 613074 91684
rect 614942 91672 614948 91684
rect 615000 91672 615006 91724
rect 590654 89632 590660 89684
rect 590712 89672 590718 89684
rect 603534 89672 603540 89684
rect 590712 89644 603540 89672
rect 590712 89632 590718 89644
rect 603534 89632 603540 89644
rect 603592 89632 603598 89684
rect 657078 88816 657084 88868
rect 657136 88856 657142 88868
rect 657998 88856 658004 88868
rect 657136 88828 658004 88856
rect 657136 88816 657142 88828
rect 657998 88816 658004 88828
rect 658056 88816 658062 88868
rect 659470 88816 659476 88868
rect 659528 88856 659534 88868
rect 663610 88856 663616 88868
rect 659528 88828 663616 88856
rect 659528 88816 659534 88828
rect 663610 88816 663616 88828
rect 663668 88816 663674 88868
rect 578142 85552 578148 85604
rect 578200 85592 578206 85604
rect 589182 85592 589188 85604
rect 578200 85564 589188 85592
rect 578200 85552 578206 85564
rect 589182 85552 589188 85564
rect 589240 85552 589246 85604
rect 648890 85484 648896 85536
rect 648948 85524 648954 85536
rect 657170 85524 657176 85536
rect 648948 85496 657176 85524
rect 648948 85484 648954 85496
rect 657170 85484 657176 85496
rect 657228 85484 657234 85536
rect 651466 85416 651472 85468
rect 651524 85456 651530 85468
rect 658826 85456 658832 85468
rect 651524 85428 658832 85456
rect 651524 85416 651530 85428
rect 658826 85416 658832 85428
rect 658884 85416 658890 85468
rect 648798 85348 648804 85400
rect 648856 85388 648862 85400
rect 660666 85388 660672 85400
rect 648856 85360 660672 85388
rect 648856 85348 648862 85360
rect 660666 85348 660672 85360
rect 660724 85348 660730 85400
rect 648706 85280 648712 85332
rect 648764 85320 648770 85332
rect 657722 85320 657728 85332
rect 648764 85292 657728 85320
rect 648764 85280 648770 85292
rect 657722 85280 657728 85292
rect 657780 85280 657786 85332
rect 643554 85212 643560 85264
rect 643612 85252 643618 85264
rect 660114 85252 660120 85264
rect 643612 85224 660120 85252
rect 643612 85212 643618 85224
rect 660114 85212 660120 85224
rect 660172 85212 660178 85264
rect 646682 85144 646688 85196
rect 646740 85184 646746 85196
rect 661402 85184 661408 85196
rect 646740 85156 661408 85184
rect 646740 85144 646746 85156
rect 661402 85144 661408 85156
rect 661460 85144 661466 85196
rect 586422 84600 586428 84652
rect 586480 84640 586486 84652
rect 600314 84640 600320 84652
rect 586480 84612 600320 84640
rect 586480 84600 586486 84612
rect 600314 84600 600320 84612
rect 600372 84600 600378 84652
rect 583846 84532 583852 84584
rect 583904 84572 583910 84584
rect 600498 84572 600504 84584
rect 583904 84544 600504 84572
rect 583904 84532 583910 84544
rect 600498 84532 600504 84544
rect 600556 84532 600562 84584
rect 583754 84464 583760 84516
rect 583812 84504 583818 84516
rect 600682 84504 600688 84516
rect 583812 84476 600688 84504
rect 583812 84464 583818 84476
rect 600682 84464 600688 84476
rect 600740 84464 600746 84516
rect 582282 84396 582288 84448
rect 582340 84436 582346 84448
rect 600222 84436 600228 84448
rect 582340 84408 600228 84436
rect 582340 84396 582346 84408
rect 600222 84396 600228 84408
rect 600280 84396 600286 84448
rect 582006 84328 582012 84380
rect 582064 84368 582070 84380
rect 600406 84368 600412 84380
rect 582064 84340 600412 84368
rect 582064 84328 582070 84340
rect 600406 84328 600412 84340
rect 600464 84328 600470 84380
rect 582190 84260 582196 84312
rect 582248 84300 582254 84312
rect 600590 84300 600596 84312
rect 582248 84272 600596 84300
rect 582248 84260 582254 84272
rect 600590 84260 600596 84272
rect 600648 84260 600654 84312
rect 582098 84192 582104 84244
rect 582156 84232 582162 84244
rect 600774 84232 600780 84244
rect 582156 84204 600780 84232
rect 582156 84192 582162 84204
rect 600774 84192 600780 84204
rect 600832 84192 600838 84244
rect 581914 84124 581920 84176
rect 581972 84164 581978 84176
rect 600866 84164 600872 84176
rect 581972 84136 600872 84164
rect 581972 84124 581978 84136
rect 600866 84124 600872 84136
rect 600924 84124 600930 84176
rect 607214 83784 607220 83836
rect 607272 83824 607278 83836
rect 612918 83824 612924 83836
rect 607272 83796 612924 83824
rect 607272 83784 607278 83796
rect 612918 83784 612924 83796
rect 612976 83784 612982 83836
rect 610158 82940 610164 82952
rect 601804 82912 610164 82940
rect 598934 82764 598940 82816
rect 598992 82804 598998 82816
rect 601804 82804 601832 82912
rect 610158 82900 610164 82912
rect 610216 82900 610222 82952
rect 605742 82832 605748 82884
rect 605800 82872 605806 82884
rect 610342 82872 610348 82884
rect 605800 82844 610348 82872
rect 605800 82832 605806 82844
rect 610342 82832 610348 82844
rect 610400 82832 610406 82884
rect 598992 82776 601832 82804
rect 598992 82764 598998 82776
rect 579614 82628 579620 82680
rect 579672 82668 579678 82680
rect 583662 82668 583668 82680
rect 579672 82640 583668 82668
rect 579672 82628 579678 82640
rect 583662 82628 583668 82640
rect 583720 82628 583726 82680
rect 580810 81472 580816 81524
rect 580868 81512 580874 81524
rect 581086 81512 581092 81524
rect 580868 81484 581092 81512
rect 580868 81472 580874 81484
rect 581086 81472 581092 81484
rect 581144 81472 581150 81524
rect 578234 75760 578240 75812
rect 578292 75800 578298 75812
rect 590654 75800 590660 75812
rect 578292 75772 590660 75800
rect 578292 75760 578298 75772
rect 590654 75760 590660 75772
rect 590712 75760 590718 75812
rect 600314 75352 600320 75404
rect 600372 75392 600378 75404
rect 607214 75392 607220 75404
rect 600372 75364 607220 75392
rect 600372 75352 600378 75364
rect 607214 75352 607220 75364
rect 607272 75352 607278 75404
rect 580994 72156 581000 72208
rect 581052 72196 581058 72208
rect 598842 72196 598848 72208
rect 581052 72168 598848 72196
rect 581052 72156 581058 72168
rect 598842 72156 598848 72168
rect 598900 72156 598906 72208
rect 629294 71952 629300 72004
rect 629352 71992 629358 72004
rect 631502 71992 631508 72004
rect 629352 71964 631508 71992
rect 629352 71952 629358 71964
rect 631502 71952 631508 71964
rect 631560 71952 631566 72004
rect 602614 71748 602620 71800
rect 602672 71788 602678 71800
rect 612826 71788 612832 71800
rect 602672 71760 612832 71788
rect 602672 71748 602678 71760
rect 612826 71748 612832 71760
rect 612884 71748 612890 71800
rect 578326 69028 578332 69080
rect 578384 69068 578390 69080
rect 580994 69068 581000 69080
rect 578384 69040 581000 69068
rect 578384 69028 578390 69040
rect 580994 69028 581000 69040
rect 581052 69028 581058 69080
rect 594702 66240 594708 66292
rect 594760 66280 594766 66292
rect 600314 66280 600320 66292
rect 594760 66252 600320 66280
rect 594760 66240 594766 66252
rect 600314 66240 600320 66252
rect 600372 66240 600378 66292
rect 587894 66172 587900 66224
rect 587952 66212 587958 66224
rect 597462 66212 597468 66224
rect 587952 66184 597468 66212
rect 587952 66172 587958 66184
rect 597462 66172 597468 66184
rect 597520 66172 597526 66224
rect 580718 65968 580724 66020
rect 580776 66008 580782 66020
rect 586422 66008 586428 66020
rect 580776 65980 586428 66008
rect 580776 65968 580782 65980
rect 586422 65968 586428 65980
rect 586480 65968 586486 66020
rect 594334 63724 594340 63776
rect 594392 63764 594398 63776
rect 605742 63764 605748 63776
rect 594392 63736 605748 63764
rect 594392 63724 594398 63736
rect 605742 63724 605748 63736
rect 605800 63724 605806 63776
rect 597554 63520 597560 63572
rect 597612 63560 597618 63572
rect 602614 63560 602620 63572
rect 597612 63532 602620 63560
rect 597612 63520 597618 63532
rect 602614 63520 602620 63532
rect 602672 63520 602678 63572
rect 579614 59848 579620 59900
rect 579672 59888 579678 59900
rect 583754 59888 583760 59900
rect 579672 59860 583760 59888
rect 579672 59848 579678 59860
rect 583754 59848 583760 59860
rect 583812 59848 583818 59900
rect 579798 59032 579804 59084
rect 579856 59072 579862 59084
rect 594334 59072 594340 59084
rect 579856 59044 594340 59072
rect 579856 59032 579862 59044
rect 594334 59032 594340 59044
rect 594392 59032 594398 59084
rect 579614 58624 579620 58676
rect 579672 58664 579678 58676
rect 583846 58664 583852 58676
rect 579672 58636 583852 58664
rect 579672 58624 579678 58636
rect 583846 58624 583852 58636
rect 583904 58624 583910 58676
rect 599118 55496 599124 55548
rect 599176 55536 599182 55548
rect 604454 55536 604460 55548
rect 599176 55508 604460 55536
rect 599176 55496 599182 55508
rect 604454 55496 604460 55508
rect 604512 55496 604518 55548
rect 579798 55264 579804 55276
rect 576872 55236 579804 55264
rect 576762 55156 576768 55208
rect 576820 55196 576826 55208
rect 576872 55196 576900 55236
rect 579798 55224 579804 55236
rect 579856 55224 579862 55276
rect 576820 55168 576900 55196
rect 576820 55156 576826 55168
rect 587894 53700 587900 53712
rect 571352 53672 587900 53700
rect 571352 53644 571380 53672
rect 587894 53660 587900 53672
rect 587952 53660 587958 53712
rect 571334 53592 571340 53644
rect 571392 53592 571398 53644
rect 346854 52368 346860 52420
rect 346912 52408 346918 52420
rect 642910 52408 642916 52420
rect 346912 52380 642916 52408
rect 346912 52368 346918 52380
rect 642910 52368 642916 52380
rect 642968 52368 642974 52420
rect 230382 51416 230388 51468
rect 230440 51456 230446 51468
rect 642818 51456 642824 51468
rect 230440 51428 642824 51456
rect 230440 51416 230446 51428
rect 642818 51416 642824 51428
rect 642876 51416 642882 51468
rect 212442 51348 212448 51400
rect 212500 51388 212506 51400
rect 639322 51388 639328 51400
rect 212500 51360 639328 51388
rect 212500 51348 212506 51360
rect 639322 51348 639328 51360
rect 639380 51348 639386 51400
rect 559466 51008 559472 51060
rect 559524 51048 559530 51060
rect 578234 51048 578240 51060
rect 559524 51020 578240 51048
rect 559524 51008 559530 51020
rect 578234 51008 578240 51020
rect 578292 51008 578298 51060
rect 578326 49756 578332 49768
rect 574066 49728 578332 49756
rect 565814 49648 565820 49700
rect 565872 49688 565878 49700
rect 574066 49688 574094 49728
rect 578326 49716 578332 49728
rect 578384 49716 578390 49768
rect 590654 49716 590660 49768
rect 590712 49756 590718 49768
rect 597554 49756 597560 49768
rect 590712 49728 597560 49756
rect 590712 49716 590718 49728
rect 597554 49716 597560 49728
rect 597612 49716 597618 49768
rect 565872 49660 574094 49688
rect 565872 49648 565878 49660
rect 478138 48492 478144 48544
rect 478196 48532 478202 48544
rect 526162 48532 526168 48544
rect 478196 48504 526168 48532
rect 478196 48492 478202 48504
rect 526162 48492 526168 48504
rect 526220 48492 526226 48544
rect 215202 48424 215208 48476
rect 215260 48464 215266 48476
rect 346486 48464 346492 48476
rect 215260 48436 346492 48464
rect 215260 48424 215266 48436
rect 346486 48424 346492 48436
rect 346544 48424 346550 48476
rect 412634 48424 412640 48476
rect 412692 48464 412698 48476
rect 494054 48464 494060 48476
rect 412692 48436 494060 48464
rect 412692 48424 412698 48436
rect 494054 48424 494060 48436
rect 494112 48424 494118 48476
rect 149974 48356 149980 48408
rect 150032 48396 150038 48408
rect 150250 48396 150256 48408
rect 150032 48368 150256 48396
rect 150032 48356 150038 48368
rect 150250 48356 150256 48368
rect 150308 48396 150314 48408
rect 218054 48396 218060 48408
rect 150308 48368 218060 48396
rect 150308 48356 150314 48368
rect 218054 48356 218060 48368
rect 218112 48356 218118 48408
rect 281442 48356 281448 48408
rect 281500 48396 281506 48408
rect 506382 48396 506388 48408
rect 281500 48368 506388 48396
rect 281500 48356 281506 48368
rect 506382 48356 506388 48368
rect 506440 48356 506446 48408
rect 216122 48288 216128 48340
rect 216180 48328 216186 48340
rect 518526 48328 518532 48340
rect 216180 48300 518532 48328
rect 216180 48288 216186 48300
rect 518526 48288 518532 48300
rect 518584 48288 518590 48340
rect 590746 48288 590752 48340
rect 590804 48328 590810 48340
rect 599118 48328 599124 48340
rect 590804 48300 599124 48328
rect 590804 48288 590810 48300
rect 599118 48288 599124 48300
rect 599176 48288 599182 48340
rect 535454 47200 535460 47252
rect 535512 47240 535518 47252
rect 542998 47240 543004 47252
rect 535512 47212 543004 47240
rect 535512 47200 535518 47212
rect 542998 47200 543004 47212
rect 543056 47200 543062 47252
rect 52086 47064 52092 47116
rect 52144 47104 52150 47116
rect 213822 47104 213828 47116
rect 52144 47076 213828 47104
rect 52144 47064 52150 47076
rect 213822 47064 213828 47076
rect 213880 47104 213886 47116
rect 215202 47104 215208 47116
rect 213880 47076 215208 47104
rect 213880 47064 213886 47076
rect 215202 47064 215208 47076
rect 215260 47064 215266 47116
rect 52270 46996 52276 47048
rect 52328 47036 52334 47048
rect 149974 47036 149980 47048
rect 52328 47008 149980 47036
rect 52328 46996 52334 47008
rect 149974 46996 149980 47008
rect 150032 46996 150038 47048
rect 494054 46860 494060 46912
rect 494112 46900 494118 46912
rect 502242 46900 502248 46912
rect 494112 46872 502248 46900
rect 494112 46860 494118 46872
rect 502242 46860 502248 46872
rect 502300 46860 502306 46912
rect 646314 46860 646320 46912
rect 646372 46900 646378 46912
rect 666554 46900 666560 46912
rect 646372 46872 666560 46900
rect 646372 46860 646378 46872
rect 666554 46860 666560 46872
rect 666612 46860 666618 46912
rect 460658 45772 460664 45824
rect 460716 45812 460722 45824
rect 610250 45812 610256 45824
rect 460716 45784 610256 45812
rect 460716 45772 460722 45784
rect 610250 45772 610256 45784
rect 610308 45772 610314 45824
rect 367094 45704 367100 45756
rect 367152 45744 367158 45756
rect 607306 45744 607312 45756
rect 367152 45716 607312 45744
rect 367152 45704 367158 45716
rect 607306 45704 607312 45716
rect 607364 45704 607370 45756
rect 312814 45636 312820 45688
rect 312872 45676 312878 45688
rect 607582 45676 607588 45688
rect 312872 45648 607588 45676
rect 312872 45636 312878 45648
rect 607582 45636 607588 45648
rect 607640 45636 607646 45688
rect 230842 45568 230848 45620
rect 230900 45608 230906 45620
rect 613010 45608 613016 45620
rect 230900 45580 613016 45608
rect 230900 45568 230906 45580
rect 613010 45568 613016 45580
rect 613068 45568 613074 45620
rect 85114 45500 85120 45552
rect 85172 45540 85178 45552
rect 475654 45540 475660 45552
rect 85172 45512 475660 45540
rect 85172 45500 85178 45512
rect 475654 45500 475660 45512
rect 475712 45500 475718 45552
rect 524046 45500 524052 45552
rect 524104 45540 524110 45552
rect 559466 45540 559472 45552
rect 524104 45512 559472 45540
rect 524104 45500 524110 45512
rect 559466 45500 559472 45512
rect 559524 45500 559530 45552
rect 312814 44180 312820 44192
rect 310440 44152 312820 44180
rect 310440 44124 310468 44152
rect 312814 44140 312820 44152
rect 312872 44140 312878 44192
rect 367094 44180 367100 44192
rect 365180 44152 367100 44180
rect 365180 44124 365208 44152
rect 367094 44140 367100 44152
rect 367152 44140 367158 44192
rect 565814 44140 565820 44192
rect 565872 44180 565878 44192
rect 571334 44180 571340 44192
rect 565872 44152 571340 44180
rect 565872 44140 565878 44152
rect 571334 44140 571340 44152
rect 571392 44140 571398 44192
rect 576762 44180 576768 44192
rect 574066 44152 576768 44180
rect 310422 44072 310428 44124
rect 310480 44072 310486 44124
rect 365162 44072 365168 44124
rect 365220 44072 365226 44124
rect 444558 44072 444564 44124
rect 444616 44112 444622 44124
rect 574066 44112 574094 44152
rect 576762 44140 576768 44152
rect 576820 44140 576826 44192
rect 590654 44180 590660 44192
rect 583680 44152 590660 44180
rect 444616 44084 574094 44112
rect 444616 44072 444622 44084
rect 474458 44004 474464 44056
rect 474516 44044 474522 44056
rect 583680 44044 583708 44152
rect 590654 44140 590660 44152
rect 590712 44140 590718 44192
rect 474516 44016 583708 44044
rect 474516 44004 474522 44016
rect 419718 43936 419724 43988
rect 419776 43976 419782 43988
rect 578142 43976 578148 43988
rect 419776 43948 578148 43976
rect 419776 43936 419782 43948
rect 578142 43936 578148 43948
rect 578200 43936 578206 43988
rect 405550 43868 405556 43920
rect 405608 43908 405614 43920
rect 607490 43908 607496 43920
rect 405608 43880 607496 43908
rect 405608 43868 405614 43880
rect 607490 43868 607496 43880
rect 607548 43868 607554 43920
rect 230566 43800 230572 43852
rect 230624 43840 230630 43852
rect 618254 43840 618260 43852
rect 230624 43812 618260 43840
rect 230624 43800 230630 43812
rect 618254 43800 618260 43812
rect 618312 43800 618318 43852
rect 231026 43732 231032 43784
rect 231084 43772 231090 43784
rect 621474 43772 621480 43784
rect 231084 43744 621480 43772
rect 231084 43732 231090 43744
rect 621474 43732 621480 43744
rect 621532 43732 621538 43784
rect 230934 43664 230940 43716
rect 230992 43704 230998 43716
rect 621198 43704 621204 43716
rect 230992 43676 621204 43704
rect 230992 43664 230998 43676
rect 621198 43664 621204 43676
rect 621256 43664 621262 43716
rect 230750 43596 230756 43648
rect 230808 43636 230814 43648
rect 621566 43636 621572 43648
rect 230808 43608 621572 43636
rect 230808 43596 230814 43608
rect 621566 43596 621572 43608
rect 621624 43596 621630 43648
rect 230658 43528 230664 43580
rect 230716 43568 230722 43580
rect 621290 43568 621296 43580
rect 230716 43540 621296 43568
rect 230716 43528 230722 43540
rect 621290 43528 621296 43540
rect 621348 43528 621354 43580
rect 230474 43460 230480 43512
rect 230532 43500 230538 43512
rect 621382 43500 621388 43512
rect 230532 43472 621388 43500
rect 230532 43460 230538 43472
rect 621382 43460 621388 43472
rect 621440 43460 621446 43512
rect 226242 43392 226248 43444
rect 226300 43432 226306 43444
rect 622486 43432 622492 43444
rect 226300 43404 622492 43432
rect 226300 43392 226306 43404
rect 622486 43392 622492 43404
rect 622544 43392 622550 43444
rect 223482 43324 223488 43376
rect 223540 43364 223546 43376
rect 622302 43364 622308 43376
rect 223540 43336 622308 43364
rect 223540 43324 223546 43336
rect 622302 43324 622308 43336
rect 622360 43324 622366 43376
rect 209682 43256 209688 43308
rect 209740 43296 209746 43308
rect 629294 43296 629300 43308
rect 209740 43268 629300 43296
rect 209740 43256 209746 43268
rect 629294 43256 629300 43268
rect 629352 43256 629358 43308
rect 615402 42916 615408 42968
rect 615460 42956 615466 42968
rect 641162 42956 641168 42968
rect 615460 42928 641168 42956
rect 615460 42916 615466 42928
rect 641162 42916 641168 42928
rect 641220 42916 641226 42968
rect 52178 42848 52184 42900
rect 52236 42888 52242 42900
rect 215294 42888 215300 42900
rect 52236 42860 215300 42888
rect 52236 42848 52242 42860
rect 215294 42848 215300 42860
rect 215352 42848 215358 42900
rect 507854 42236 507860 42288
rect 507912 42276 507918 42288
rect 530670 42276 530676 42288
rect 507912 42248 530676 42276
rect 507912 42236 507918 42248
rect 530670 42236 530676 42248
rect 530728 42236 530734 42288
rect 531038 42236 531044 42288
rect 531096 42276 531102 42288
rect 565722 42276 565728 42288
rect 531096 42248 565728 42276
rect 531096 42236 531102 42248
rect 565722 42236 565728 42248
rect 565780 42236 565786 42288
rect 506382 41896 506388 41948
rect 506440 41936 506446 41948
rect 520366 41936 520372 41948
rect 506440 41908 520372 41936
rect 506440 41896 506446 41908
rect 520366 41896 520372 41908
rect 520424 41896 520430 41948
rect 502242 41828 502248 41880
rect 502300 41868 502306 41880
rect 518526 41868 518532 41880
rect 502300 41840 518532 41868
rect 502300 41828 502306 41840
rect 518526 41828 518532 41840
rect 518584 41828 518590 41880
rect 416682 41760 416688 41812
rect 416740 41800 416746 41812
rect 420730 41800 420736 41812
rect 416740 41772 420736 41800
rect 416740 41760 416746 41772
rect 420730 41760 420736 41772
rect 420788 41760 420794 41812
rect 471698 41760 471704 41812
rect 471756 41800 471762 41812
rect 475562 41800 475568 41812
rect 471756 41772 475568 41800
rect 471756 41760 471762 41772
rect 475562 41760 475568 41772
rect 475620 41760 475626 41812
rect 514018 41760 514024 41812
rect 514076 41800 514082 41812
rect 514846 41800 514852 41812
rect 514076 41772 514852 41800
rect 514076 41760 514082 41772
rect 514846 41760 514852 41772
rect 514904 41760 514910 41812
rect 141786 41488 141792 41540
rect 141844 41528 141850 41540
rect 207014 41528 207020 41540
rect 141844 41500 207020 41528
rect 141844 41488 141850 41500
rect 207014 41488 207020 41500
rect 207072 41528 207078 41540
rect 209682 41528 209688 41540
rect 207072 41500 209688 41528
rect 207072 41488 207078 41500
rect 209682 41488 209688 41500
rect 209740 41488 209746 41540
rect 444558 38672 444564 38684
rect 444300 38644 444564 38672
rect 420730 38564 420736 38616
rect 420788 38604 420794 38616
rect 444300 38604 444328 38644
rect 444558 38632 444564 38644
rect 444616 38632 444622 38684
rect 420788 38576 444328 38604
rect 420788 38564 420794 38576
rect 475562 38564 475568 38616
rect 475620 38604 475626 38616
rect 507854 38604 507860 38616
rect 475620 38576 507860 38604
rect 475620 38564 475626 38576
rect 507854 38564 507860 38576
rect 507912 38564 507918 38616
rect 475654 38496 475660 38548
rect 475712 38536 475718 38548
rect 514018 38536 514024 38548
rect 475712 38508 514024 38536
rect 475712 38496 475718 38508
rect 514018 38496 514024 38508
rect 514076 38496 514082 38548
rect 213178 24760 213184 24812
rect 213236 24800 213242 24812
rect 213822 24800 213828 24812
rect 213236 24772 213828 24800
rect 213236 24760 213242 24772
rect 213822 24760 213828 24772
rect 213880 24760 213886 24812
rect 224586 22992 224592 23044
rect 224644 23032 224650 23044
rect 226242 23032 226248 23044
rect 224644 23004 226248 23032
rect 224644 22992 224650 23004
rect 226242 22992 226248 23004
rect 226300 22992 226306 23044
rect 221734 22516 221740 22568
rect 221792 22556 221798 22568
rect 223482 22556 223488 22568
rect 221792 22528 223488 22556
rect 221792 22516 221798 22528
rect 223482 22516 223488 22528
rect 223540 22516 223546 22568
<< via1 >>
rect 425980 1006000 426032 1006052
rect 458916 1006000 458968 1006052
rect 424324 1005864 424376 1005916
rect 440424 1005864 440476 1005916
rect 423864 1005796 423916 1005848
rect 440240 1005796 440292 1005848
rect 504548 1005660 504600 1005712
rect 519728 1005660 519780 1005712
rect 356060 1005592 356112 1005644
rect 373172 1005592 373224 1005644
rect 505008 1005592 505060 1005644
rect 517428 1005592 517480 1005644
rect 356888 1005524 356940 1005576
rect 378048 1005524 378100 1005576
rect 505376 1005524 505428 1005576
rect 518808 1005524 518860 1005576
rect 502984 1005456 503036 1005508
rect 523040 1005456 523092 1005508
rect 144828 1005388 144880 1005440
rect 160284 1005388 160336 1005440
rect 356520 1005388 356572 1005440
rect 376668 1005388 376720 1005440
rect 425152 1005388 425204 1005440
rect 467932 1005388 467984 1005440
rect 209228 1005320 209280 1005372
rect 227720 1005320 227772 1005372
rect 253296 1005320 253348 1005372
rect 280068 1005320 280120 1005372
rect 361028 1005320 361080 1005372
rect 377956 1005320 378008 1005372
rect 428372 1005320 428424 1005372
rect 453948 1005320 454000 1005372
rect 505836 1005320 505888 1005372
rect 517060 1005320 517112 1005372
rect 92664 1005252 92716 1005304
rect 109316 1005252 109368 1005304
rect 259828 1005252 259880 1005304
rect 280252 1005252 280304 1005304
rect 106464 1005184 106516 1005236
rect 125784 1005184 125836 1005236
rect 260196 1005184 260248 1005236
rect 265072 1005184 265124 1005236
rect 360200 1005184 360252 1005236
rect 380808 1005184 380860 1005236
rect 105636 1005116 105688 1005168
rect 125600 1005116 125652 1005168
rect 195336 1005116 195388 1005168
rect 209596 1005116 209648 1005168
rect 210884 1005116 210936 1005168
rect 227904 1005116 227956 1005168
rect 263048 1005116 263100 1005168
rect 264336 1005116 264388 1005168
rect 427544 1005116 427596 1005168
rect 460848 1005116 460900 1005168
rect 201500 1005048 201552 1005100
rect 202328 1005048 202380 1005100
rect 227628 1005048 227680 1005100
rect 261024 1005048 261076 1005100
rect 265256 1005048 265308 1005100
rect 428832 1005048 428884 1005100
rect 465264 1005048 465316 1005100
rect 502524 1005048 502576 1005100
rect 523224 1005048 523276 1005100
rect 150900 1004980 150952 1005032
rect 175188 1004980 175240 1005032
rect 252836 1004980 252888 1005032
rect 253296 1004980 253348 1005032
rect 260656 1004980 260708 1005032
rect 157800 1004912 157852 1004964
rect 174084 1004912 174136 1004964
rect 208400 1004912 208452 1004964
rect 227812 1004912 227864 1004964
rect 262680 1004912 262732 1004964
rect 264336 1004912 264388 1004964
rect 358176 1004980 358228 1005032
rect 383292 1004980 383344 1005032
rect 426808 1004980 426860 1005032
rect 455604 1004980 455656 1005032
rect 504180 1004980 504232 1005032
rect 519084 1004980 519136 1005032
rect 280160 1004912 280212 1004964
rect 425520 1004912 425572 1004964
rect 455420 1004912 455472 1004964
rect 552756 1004912 552808 1004964
rect 568580 1004912 568632 1004964
rect 108028 1004844 108080 1004896
rect 109684 1004844 109736 1004896
rect 261852 1004844 261904 1004896
rect 266268 1004844 266320 1004896
rect 427176 1004844 427228 1004896
rect 455512 1004844 455564 1004896
rect 114652 1004776 114704 1004828
rect 125692 1004776 125744 1004828
rect 156972 1004776 157024 1004828
rect 173992 1004776 174044 1004828
rect 423496 1004776 423548 1004828
rect 467748 1004776 467800 1004828
rect 553124 1004776 553176 1004828
rect 557448 1004776 557500 1004828
rect 99472 1004708 99524 1004760
rect 92940 1004640 92992 1004692
rect 108856 1004640 108908 1004692
rect 154488 1004708 154540 1004760
rect 125508 1004640 125560 1004692
rect 146024 1004640 146076 1004692
rect 154948 1004640 155000 1004692
rect 159456 1004708 159508 1004760
rect 173900 1004708 173952 1004760
rect 195980 1004708 196032 1004760
rect 206376 1004708 206428 1004760
rect 262220 1004708 262272 1004760
rect 280344 1004708 280396 1004760
rect 358544 1004708 358596 1004760
rect 160652 1004640 160704 1004692
rect 195704 1004640 195756 1004692
rect 205180 1004640 205232 1004692
rect 261484 1004640 261536 1004692
rect 265164 1004640 265216 1004692
rect 315120 1004640 315172 1004692
rect 331220 1004640 331272 1004692
rect 359740 1004640 359792 1004692
rect 369860 1004640 369912 1004692
rect 424692 1004708 424744 1004760
rect 467840 1004708 467892 1004760
rect 501696 1004708 501748 1004760
rect 509148 1004708 509200 1004760
rect 551928 1004708 551980 1004760
rect 558736 1004708 558788 1004760
rect 381728 1004640 381780 1004692
rect 419448 1004640 419500 1004692
rect 422300 1004640 422352 1004692
rect 458916 1004640 458968 1004692
rect 472348 1004640 472400 1004692
rect 496728 1004640 496780 1004692
rect 499304 1004640 499356 1004692
rect 502156 1004640 502208 1004692
rect 509240 1004640 509292 1004692
rect 554320 1004640 554372 1004692
rect 195152 1004572 195204 1004624
rect 205916 1004572 205968 1004624
rect 517428 1004572 517480 1004624
rect 523960 1004572 524012 1004624
rect 561312 1004640 561364 1004692
rect 567476 1004640 567528 1004692
rect 571340 1004572 571392 1004624
rect 557448 1004096 557500 1004148
rect 570144 1004096 570196 1004148
rect 553952 1003892 554004 1003944
rect 571432 1003892 571484 1003944
rect 455420 1003348 455472 1003400
rect 464252 1003348 464304 1003400
rect 455512 1003280 455564 1003332
rect 469128 1003280 469180 1003332
rect 555516 1003280 555568 1003332
rect 574008 1003280 574060 1003332
rect 455604 1003212 455656 1003264
rect 466460 1003212 466512 1003264
rect 554780 1003212 554832 1003264
rect 569960 1003212 570012 1003264
rect 440424 1001988 440476 1002040
rect 440240 1001920 440292 1001972
rect 447140 1001852 447192 1001904
rect 447324 1001852 447376 1001904
rect 466460 1001852 466512 1001904
rect 469772 1001852 469824 1001904
rect 517060 1001852 517112 1001904
rect 519544 1001852 519596 1001904
rect 519728 1001852 519780 1001904
rect 523868 1001852 523920 1001904
rect 558736 1001852 558788 1001904
rect 569868 1001852 569920 1001904
rect 568580 1001784 568632 1001836
rect 572628 1001784 572680 1001836
rect 464252 1001716 464304 1001768
rect 471704 1001716 471756 1001768
rect 376668 1001104 376720 1001156
rect 378324 1001104 378376 1001156
rect 373172 1001036 373224 1001088
rect 381268 1001036 381320 1001088
rect 360568 1000696 360620 1000748
rect 383568 1000696 383620 1000748
rect 361396 1000628 361448 1000680
rect 383384 1000628 383436 1000680
rect 369860 1000560 369912 1000612
rect 383476 1000560 383528 1000612
rect 428004 1000560 428056 1000612
rect 472624 1000560 472676 1000612
rect 358912 1000492 358964 1000544
rect 383568 1000492 383620 1000544
rect 426348 1000492 426400 1000544
rect 472532 1000492 472584 1000544
rect 380900 1000288 380952 1000340
rect 383568 1000288 383620 1000340
rect 503352 999948 503404 1000000
rect 516048 999948 516100 1000000
rect 92572 999880 92624 999932
rect 116032 999880 116084 999932
rect 246764 999880 246816 999932
rect 258632 999880 258684 999932
rect 92480 999812 92532 999864
rect 104348 999812 104400 999864
rect 246580 999812 246632 999864
rect 257344 999812 257396 999864
rect 312176 999812 312228 999864
rect 318892 999812 318944 999864
rect 92296 999744 92348 999796
rect 102784 999744 102836 999796
rect 246672 999744 246724 999796
rect 256976 999744 257028 999796
rect 311440 999744 311492 999796
rect 315948 999744 316000 999796
rect 246948 999676 247000 999728
rect 257804 999676 257856 999728
rect 313832 999676 313884 999728
rect 318708 999676 318760 999728
rect 92388 999608 92440 999660
rect 102324 999608 102376 999660
rect 195244 999608 195296 999660
rect 205548 999608 205600 999660
rect 310152 999608 310204 999660
rect 314936 999608 314988 999660
rect 155776 999540 155828 999592
rect 160284 999540 160336 999592
rect 195612 999540 195664 999592
rect 203524 999540 203576 999592
rect 313004 999540 313056 999592
rect 317604 999540 317656 999592
rect 92756 999472 92808 999524
rect 101956 999472 102008 999524
rect 159088 999472 159140 999524
rect 162860 999472 162912 999524
rect 195428 999472 195480 999524
rect 203892 999472 203944 999524
rect 314660 999472 314712 999524
rect 319076 999472 319128 999524
rect 99288 999404 99340 999456
rect 103152 999404 103204 999456
rect 195520 999404 195572 999456
rect 202328 999404 202380 999456
rect 309784 999404 309836 999456
rect 314844 999404 314896 999456
rect 198372 999336 198424 999388
rect 204720 999336 204772 999388
rect 312636 999336 312688 999388
rect 317420 999336 317472 999388
rect 198464 999268 198516 999320
rect 204352 999268 204404 999320
rect 310980 999268 311032 999320
rect 315028 999268 315080 999320
rect 198648 999200 198700 999252
rect 202696 999200 202748 999252
rect 253848 999200 253900 999252
rect 256516 999200 256568 999252
rect 311808 999200 311860 999252
rect 315120 999200 315172 999252
rect 357348 999200 357400 999252
rect 364892 999200 364944 999252
rect 198556 999132 198608 999184
rect 203064 999132 203116 999184
rect 258540 999132 258592 999184
rect 262220 999132 262272 999184
rect 314292 999132 314344 999184
rect 317512 999132 317564 999184
rect 357716 999132 357768 999184
rect 365076 999132 365128 999184
rect 378048 999132 378100 999184
rect 383200 999132 383252 999184
rect 400036 999132 400088 999184
rect 434628 999812 434680 999864
rect 430856 999744 430908 999796
rect 438124 999744 438176 999796
rect 508688 999744 508740 999796
rect 515220 999744 515272 999796
rect 431684 999676 431736 999728
rect 437940 999676 437992 999728
rect 506204 999676 506256 999728
rect 511908 999676 511960 999728
rect 429200 999608 429252 999660
rect 434720 999608 434772 999660
rect 507032 999608 507084 999660
rect 512092 999608 512144 999660
rect 430028 999540 430080 999592
rect 434812 999540 434864 999592
rect 508228 999540 508280 999592
rect 513472 999540 513524 999592
rect 431224 999472 431276 999524
rect 436192 999472 436244 999524
rect 507860 999472 507912 999524
rect 512276 999472 512328 999524
rect 429660 999404 429712 999456
rect 433432 999404 433484 999456
rect 506572 999404 506624 999456
rect 510896 999404 510948 999456
rect 432512 999336 432564 999388
rect 437388 999336 437440 999388
rect 500500 999336 500552 999388
rect 508780 999336 508832 999388
rect 509056 999336 509108 999388
rect 513656 999336 513708 999388
rect 432880 999268 432932 999320
rect 437572 999268 437624 999320
rect 509516 999268 509568 999320
rect 514852 999268 514904 999320
rect 432052 999200 432104 999252
rect 436100 999200 436152 999252
rect 500868 999200 500920 999252
rect 430396 999132 430448 999184
rect 433340 999132 433392 999184
rect 465264 999132 465316 999184
rect 472440 999132 472492 999184
rect 488908 999132 488960 999184
rect 505652 999132 505704 999184
rect 507400 999200 507452 999252
rect 510712 999200 510764 999252
rect 540336 999200 540388 999252
rect 566556 1000016 566608 1000068
rect 560852 999744 560904 999796
rect 567108 999744 567160 999796
rect 560484 999608 560536 999660
rect 565820 999608 565872 999660
rect 590660 999472 590712 999524
rect 625804 999472 625856 999524
rect 610072 999404 610124 999456
rect 625712 999404 625764 999456
rect 609980 999336 610032 999388
rect 625620 999336 625672 999388
rect 601608 999268 601660 999320
rect 625804 999268 625856 999320
rect 593420 999200 593472 999252
rect 625528 999200 625580 999252
rect 509516 999132 509568 999184
rect 509884 999132 509936 999184
rect 514668 999132 514720 999184
rect 552296 999132 552348 999184
rect 558920 999132 558972 999184
rect 144276 999064 144328 999116
rect 158260 999064 158312 999116
rect 246580 999064 246632 999116
rect 265164 999064 265216 999116
rect 298744 999064 298796 999116
rect 317604 999064 317656 999116
rect 399944 999064 399996 999116
rect 436192 999064 436244 999116
rect 453948 999064 454000 999116
rect 462596 999064 462648 999116
rect 489460 999064 489512 999116
rect 513472 999064 513524 999116
rect 508780 998996 508832 999048
rect 521292 998996 521344 999048
rect 509148 998928 509200 998980
rect 521384 998928 521436 998980
rect 509240 998860 509292 998912
rect 520556 998860 520608 998912
rect 509516 998792 509568 998844
rect 521476 998792 521528 998844
rect 364892 998452 364944 998504
rect 374552 998452 374604 998504
rect 467840 998316 467892 998368
rect 469220 998316 469272 998368
rect 467932 998180 467984 998232
rect 471060 998180 471112 998232
rect 518900 998180 518952 998232
rect 521660 998180 521712 998232
rect 467748 998044 467800 998096
rect 469312 998044 469364 998096
rect 558920 997908 558972 997960
rect 568672 997908 568724 997960
rect 365076 997772 365128 997824
rect 374460 997772 374512 997824
rect 143816 997704 143868 997756
rect 156144 997704 156196 997756
rect 501328 997704 501380 997756
rect 521568 997704 521620 997756
rect 553492 997704 553544 997756
rect 568580 997704 568632 997756
rect 569868 997704 569920 997756
rect 623780 997704 623832 997756
rect 556344 997636 556396 997688
rect 601608 997636 601660 997688
rect 571340 997568 571392 997620
rect 609980 997568 610032 997620
rect 569960 997500 570012 997552
rect 610072 997500 610124 997552
rect 557172 997432 557224 997484
rect 620928 997432 620980 997484
rect 571432 997364 571484 997416
rect 590660 997364 590712 997416
rect 572628 997296 572680 997348
rect 593420 997296 593472 997348
rect 107660 997160 107712 997212
rect 115940 997160 115992 997212
rect 210424 997160 210476 997212
rect 215300 997160 215352 997212
rect 363420 997160 363472 997212
rect 367100 997160 367152 997212
rect 96528 996412 96580 996464
rect 101128 996412 101180 996464
rect 148876 996412 148928 996464
rect 154120 996412 154172 996464
rect 146208 996344 146260 996396
rect 151728 996344 151780 996396
rect 301780 996276 301832 996328
rect 308128 996276 308180 996328
rect 146116 996208 146168 996260
rect 153752 996208 153804 996260
rect 125692 996140 125744 996192
rect 159456 996140 159508 996192
rect 173900 996140 173952 996192
rect 211252 996208 211304 996260
rect 300216 996208 300268 996260
rect 308956 996208 309008 996260
rect 365444 996208 365496 996260
rect 371148 996208 371200 996260
rect 96528 996072 96580 996124
rect 100300 996072 100352 996124
rect 108856 996072 108908 996124
rect 113272 996072 113324 996124
rect 125784 996072 125836 996124
rect 157800 996072 157852 996124
rect 173992 996072 174044 996124
rect 208768 996140 208820 996192
rect 212816 996140 212868 996192
rect 227904 996140 227956 996192
rect 267832 996140 267884 996192
rect 270408 996140 270460 996192
rect 280160 996140 280212 996192
rect 317420 996140 317472 996192
rect 364248 996140 364300 996192
rect 367284 996140 367336 996192
rect 512276 996140 512328 996192
rect 559288 996140 559340 996192
rect 204168 996072 204220 996124
rect 211620 996072 211672 996124
rect 227812 996072 227864 996124
rect 265072 996072 265124 996124
rect 267648 996072 267700 996124
rect 280344 996072 280396 996124
rect 317512 996072 317564 996124
rect 364708 996072 364760 996124
rect 369860 996072 369912 996124
rect 558460 996072 558512 996124
rect 564440 996072 564492 996124
rect 96436 996004 96488 996056
rect 101496 996004 101548 996056
rect 108488 996004 108540 996056
rect 113180 996004 113232 996056
rect 125600 996004 125652 996056
rect 156972 996004 157024 996056
rect 160192 996004 160244 996056
rect 174084 996004 174136 996056
rect 209596 996004 209648 996056
rect 212632 996004 212684 996056
rect 227720 996004 227772 996056
rect 265256 996004 265308 996056
rect 267556 996004 267608 996056
rect 280252 996004 280304 996056
rect 315120 996004 315172 996056
rect 365076 996004 365128 996056
rect 371332 996004 371384 996056
rect 625528 996004 625580 996056
rect 86040 995800 86092 995852
rect 100760 995800 100812 995852
rect 136272 995800 136324 995852
rect 154580 995936 154632 995988
rect 211252 995936 211304 995988
rect 215484 995936 215536 995988
rect 151268 995868 151320 995920
rect 136824 995800 136876 995852
rect 137928 995800 137980 995852
rect 150900 995800 150952 995852
rect 91560 995732 91612 995784
rect 92296 995732 92348 995784
rect 139216 995732 139268 995784
rect 152556 995732 152608 995784
rect 184480 995732 184532 995784
rect 198464 995868 198516 995920
rect 246488 995868 246540 995920
rect 307760 995936 307812 995988
rect 362592 995936 362644 995988
rect 367376 995936 367428 995988
rect 383476 995936 383528 995988
rect 306932 995868 306984 995920
rect 383200 995868 383252 995920
rect 188160 995800 188212 995852
rect 198648 995800 198700 995852
rect 239036 995800 239088 995852
rect 239588 995800 239640 995852
rect 254124 995800 254176 995852
rect 286784 995800 286836 995852
rect 293592 995800 293644 995852
rect 295064 995800 295116 995852
rect 310152 995800 310204 995852
rect 566556 995936 566608 995988
rect 576308 995936 576360 995988
rect 625620 995936 625672 995988
rect 472440 995868 472492 995920
rect 523040 995868 523092 995920
rect 625712 995868 625764 995920
rect 391940 995800 391992 995852
rect 396632 995800 396684 995852
rect 400036 995800 400088 995852
rect 472532 995800 472584 995852
rect 474004 995800 474056 995852
rect 474740 995800 474792 995852
rect 485688 995800 485740 995852
rect 488908 995800 488960 995852
rect 523960 995800 524012 995852
rect 524788 995800 524840 995852
rect 528468 995800 528520 995852
rect 537024 995800 537076 995852
rect 540336 995800 540388 995852
rect 625804 995800 625856 995852
rect 626540 995800 626592 995852
rect 627184 995800 627236 995852
rect 630220 995800 630272 995852
rect 631508 995800 631560 995852
rect 194324 995732 194376 995784
rect 195244 995732 195296 995784
rect 245568 995732 245620 995784
rect 246672 995732 246724 995784
rect 383660 995732 383712 995784
rect 384948 995732 385000 995784
rect 389364 995732 389416 995784
rect 472624 995732 472676 995784
rect 473268 995732 473320 995784
rect 524052 995732 524104 995784
rect 525340 995732 525392 995784
rect 620928 995732 620980 995784
rect 627828 995732 627880 995784
rect 89720 995664 89772 995716
rect 92480 995664 92532 995716
rect 190644 995664 190696 995716
rect 195428 995664 195480 995716
rect 243912 995664 243964 995716
rect 246764 995664 246816 995716
rect 291752 995664 291804 995716
rect 306472 995664 306524 995716
rect 383752 995664 383804 995716
rect 384396 995664 384448 995716
rect 472348 995664 472400 995716
rect 476948 995664 477000 995716
rect 523224 995664 523276 995716
rect 529020 995664 529072 995716
rect 625896 995664 625948 995716
rect 630864 995664 630916 995716
rect 77944 995596 77996 995648
rect 92388 995596 92440 995648
rect 133144 995596 133196 995648
rect 152924 995596 152976 995648
rect 189448 995596 189500 995648
rect 195520 995596 195572 995648
rect 240876 995596 240928 995648
rect 253664 995596 253716 995648
rect 287520 995596 287572 995648
rect 307300 995596 307352 995648
rect 383384 995596 383436 995648
rect 385684 995596 385736 995648
rect 469220 995596 469272 995648
rect 481916 995596 481968 995648
rect 521476 995596 521528 995648
rect 532700 995596 532752 995648
rect 623780 995596 623832 995648
rect 635832 995596 635884 995648
rect 88984 995528 89036 995580
rect 92572 995528 92624 995580
rect 132408 995528 132460 995580
rect 153384 995528 153436 995580
rect 184664 995528 184716 995580
rect 198556 995528 198608 995580
rect 383568 995528 383620 995580
rect 387524 995528 387576 995580
rect 469312 995528 469364 995580
rect 482652 995528 482704 995580
rect 521384 995528 521436 995580
rect 533436 995528 533488 995580
rect 130016 995460 130068 995512
rect 143816 995460 143868 995512
rect 188804 995460 188856 995512
rect 195612 995460 195664 995512
rect 383292 995460 383344 995512
rect 388628 995460 388680 995512
rect 131856 995392 131908 995444
rect 146024 995392 146076 995444
rect 183836 995392 183888 995444
rect 198372 995392 198424 995444
rect 381268 995392 381320 995444
rect 393596 995460 393648 995512
rect 183284 995324 183336 995376
rect 195980 995324 196032 995376
rect 180478 995256 180530 995308
rect 195704 995256 195756 995308
rect 303528 994720 303580 994772
rect 283472 993828 283524 993880
rect 301780 993828 301832 993880
rect 378324 993828 378376 993880
rect 392676 993828 392728 993880
rect 129096 993692 129148 993744
rect 146116 993760 146168 993812
rect 285956 993760 286008 993812
rect 314844 993760 314896 993812
rect 469772 993760 469824 993812
rect 487804 993760 487856 993812
rect 520556 993760 520608 993812
rect 535552 993760 535604 993812
rect 140504 993692 140556 993744
rect 151820 993692 151872 993744
rect 180156 993692 180208 993744
rect 207020 993692 207072 993744
rect 284116 993692 284168 993744
rect 315028 993692 315080 993744
rect 374552 993692 374604 993744
rect 393320 993692 393372 993744
rect 471060 993692 471112 993744
rect 484124 993692 484176 993744
rect 574100 993692 574152 993744
rect 633992 993692 634044 993744
rect 77024 993624 77076 993676
rect 104164 993624 104216 993676
rect 128452 993624 128504 993676
rect 160284 993624 160336 993676
rect 181444 993624 181496 993676
rect 207756 993624 207808 993676
rect 231584 993624 231636 993676
rect 262220 993624 262272 993676
rect 282828 993624 282880 993676
rect 314936 993624 314988 993676
rect 359188 993624 359240 993676
rect 398840 993624 398892 993676
rect 462596 993624 462648 993676
rect 485964 993624 486016 993676
rect 503628 993624 503680 993676
rect 539232 993624 539284 993676
rect 555056 993624 555108 993676
rect 640708 993624 640760 993676
rect 433524 993556 433576 993608
rect 434720 993556 434772 993608
rect 510896 993556 510948 993608
rect 510988 993556 511040 993608
rect 512092 993556 512144 993608
rect 558552 993556 558604 993608
rect 367376 993488 367428 993540
rect 368572 993488 368624 993540
rect 433340 993488 433392 993540
rect 433616 993488 433668 993540
rect 434812 993488 434864 993540
rect 510712 993488 510764 993540
rect 510804 993488 510856 993540
rect 511908 993488 511960 993540
rect 557724 993488 557776 993540
rect 367284 993420 367336 993472
rect 368388 993420 368440 993472
rect 368756 993420 368808 993472
rect 433432 993420 433484 993472
rect 436192 993420 436244 993472
rect 437940 993420 437992 993472
rect 513656 993420 513708 993472
rect 513748 993420 513800 993472
rect 515220 993420 515272 993472
rect 565820 993420 565872 993472
rect 436100 993352 436152 993404
rect 367468 992536 367520 992588
rect 368756 992536 368808 992588
rect 116032 990836 116084 990888
rect 122104 990768 122156 990820
rect 168380 990632 168432 990684
rect 170404 990632 170456 990684
rect 203156 990632 203208 990684
rect 204168 990632 204220 990684
rect 331220 990632 331272 990684
rect 332692 990632 332744 990684
rect 89628 990088 89680 990140
rect 92480 990088 92532 990140
rect 366180 989680 366232 989732
rect 381636 989680 381688 989732
rect 434628 989680 434680 989732
rect 446496 989680 446548 989732
rect 371148 989612 371200 989664
rect 397828 989612 397880 989664
rect 437572 989612 437624 989664
rect 462780 989612 462832 989664
rect 514668 989612 514720 989664
rect 527640 989612 527692 989664
rect 567476 989612 567528 989664
rect 592500 989612 592552 989664
rect 321468 989544 321520 989596
rect 349160 989544 349212 989596
rect 371516 989544 371568 989596
rect 414112 989544 414164 989596
rect 437756 989544 437808 989596
rect 478972 989544 479024 989596
rect 515036 989544 515088 989596
rect 543832 989544 543884 989596
rect 567292 989544 567344 989596
rect 608784 989544 608836 989596
rect 269212 989476 269264 989528
rect 300492 989476 300544 989528
rect 319076 989476 319128 989528
rect 365444 989476 365496 989528
rect 371332 989476 371384 989528
rect 430304 989476 430356 989528
rect 437388 989476 437440 989528
rect 495164 989476 495216 989528
rect 514852 989476 514904 989528
rect 560116 989476 560168 989528
rect 567108 989476 567160 989528
rect 624976 989476 625028 989528
rect 73436 989408 73488 989460
rect 92940 989408 92992 989460
rect 105820 989408 105872 989460
rect 113272 989408 113324 989460
rect 151820 989408 151872 989460
rect 186964 989408 187016 989460
rect 216588 989408 216640 989460
rect 235632 989408 235684 989460
rect 269028 989408 269080 989460
rect 284300 989408 284352 989460
rect 303528 989408 303580 989460
rect 666560 989408 666612 989460
rect 138296 988728 138348 988780
rect 144828 988728 144880 988780
rect 505652 988252 505704 988304
rect 511448 988252 511500 988304
rect 248328 988116 248380 988168
rect 251824 988116 251876 988168
rect 45468 987980 45520 988032
rect 367192 987980 367244 988032
rect 45744 987912 45796 987964
rect 368756 987912 368808 987964
rect 45560 987844 45612 987896
rect 369860 987844 369912 987896
rect 318892 987776 318944 987828
rect 666652 987776 666704 987828
rect 317512 987708 317564 987760
rect 666928 987708 666980 987760
rect 318708 987640 318760 987692
rect 669228 987640 669280 987692
rect 315120 987572 315172 987624
rect 666744 987572 666796 987624
rect 280068 987504 280120 987556
rect 651380 987504 651432 987556
rect 270408 987436 270460 987488
rect 652852 987436 652904 987488
rect 267648 987368 267700 987420
rect 652668 987368 652720 987420
rect 48228 987300 48280 987352
rect 433524 987300 433576 987352
rect 267556 987232 267608 987284
rect 652760 987232 652812 987284
rect 227628 987164 227680 987216
rect 651564 987164 651616 987216
rect 215484 987096 215536 987148
rect 658280 987096 658332 987148
rect 212816 987028 212868 987080
rect 658188 987028 658240 987080
rect 175188 986960 175240 987012
rect 651656 986960 651708 987012
rect 125508 986892 125560 986944
rect 651472 986892 651524 986944
rect 62672 986824 62724 986876
rect 113180 986824 113232 986876
rect 669504 986824 669556 986876
rect 62304 986756 62356 986808
rect 110604 986756 110656 986808
rect 669412 986756 669464 986808
rect 62488 986688 62540 986740
rect 110788 986688 110840 986740
rect 669320 986688 669372 986740
rect 564532 985532 564584 985584
rect 564716 985532 564768 985584
rect 675668 985532 675720 985584
rect 62856 985464 62908 985516
rect 669596 985464 669648 985516
rect 62580 985396 62632 985448
rect 670424 985396 670476 985448
rect 46480 985328 46532 985380
rect 668768 985328 668820 985380
rect 350264 985124 350316 985176
rect 670976 985124 671028 985176
rect 45652 985056 45704 985108
rect 367100 985056 367152 985108
rect 45928 984988 45980 985040
rect 368572 984988 368624 985040
rect 45836 984920 45888 984972
rect 368388 984920 368440 984972
rect 419448 984920 419500 984972
rect 670884 984920 670936 984972
rect 317420 984852 317472 984904
rect 666836 984852 666888 984904
rect 315948 984784 316000 984836
rect 671988 984784 672040 984836
rect 300768 984716 300820 984768
rect 671068 984716 671120 984768
rect 46112 984648 46164 984700
rect 433616 984648 433668 984700
rect 48320 984580 48372 984632
rect 436192 984580 436244 984632
rect 496728 984580 496780 984632
rect 670792 984580 670844 984632
rect 212632 984512 212684 984564
rect 652944 984512 652996 984564
rect 46388 984444 46440 984496
rect 510988 984444 511040 984496
rect 46204 984376 46256 984428
rect 510804 984376 510856 984428
rect 48412 984308 48464 984360
rect 513748 984308 513800 984360
rect 546316 984308 546368 984360
rect 670700 984308 670752 984360
rect 162860 984240 162912 984292
rect 655428 984240 655480 984292
rect 162952 984172 163004 984224
rect 658464 984172 658516 984224
rect 46020 984104 46072 984156
rect 110420 984104 110472 984156
rect 160192 984104 160244 984156
rect 658372 984104 658424 984156
rect 62028 984036 62080 984088
rect 561680 984036 561732 984088
rect 564348 984036 564400 984088
rect 649908 984036 649960 984088
rect 62120 983968 62172 984020
rect 564532 983968 564584 984020
rect 62212 983900 62264 983952
rect 564440 983900 564492 983952
rect 62396 982948 62448 983000
rect 669044 982948 669096 983000
rect 62764 982880 62816 982932
rect 668676 982880 668728 982932
rect 42340 972884 42392 972936
rect 58440 972884 58492 972936
rect 674840 970096 674892 970148
rect 675668 970096 675720 970148
rect 42156 967240 42208 967292
rect 42340 967240 42392 967292
rect 42064 967036 42116 967088
rect 42800 967036 42852 967088
rect 674748 966152 674800 966204
rect 675392 966152 675444 966204
rect 673552 965744 673604 965796
rect 675392 965744 675444 965796
rect 673736 964996 673788 965048
rect 675484 964996 675536 965048
rect 42156 963976 42208 964028
rect 42984 963976 43036 964028
rect 673920 963160 673972 963212
rect 675392 963160 675444 963212
rect 42156 962616 42208 962668
rect 42892 962616 42944 962668
rect 673644 962480 673696 962532
rect 675484 962480 675536 962532
rect 42156 962072 42208 962124
rect 43076 962072 43128 962124
rect 673460 962004 673512 962056
rect 675392 962004 675444 962056
rect 673828 961324 673880 961376
rect 675392 961324 675444 961376
rect 48504 960508 48556 960560
rect 57980 960508 58032 960560
rect 655612 960508 655664 960560
rect 675024 960508 675076 960560
rect 42892 959624 42944 959676
rect 43628 959624 43680 959676
rect 42064 959488 42116 959540
rect 42892 959488 42944 959540
rect 42156 959080 42208 959132
rect 43352 959080 43404 959132
rect 674656 958808 674708 958860
rect 675392 958808 675444 958860
rect 42064 958332 42116 958384
rect 43168 958332 43220 958384
rect 674288 958332 674340 958384
rect 675392 958332 675444 958384
rect 42064 957720 42116 957772
rect 43260 957720 43312 957772
rect 674380 957720 674432 957772
rect 675484 957720 675536 957772
rect 674564 956972 674616 957024
rect 675392 956972 675444 957024
rect 674472 955680 674524 955732
rect 675484 955680 675536 955732
rect 675024 955476 675076 955528
rect 675484 955476 675536 955528
rect 42156 955340 42208 955392
rect 42708 955340 42760 955392
rect 674012 953980 674064 954032
rect 674748 953980 674800 954032
rect 674748 953844 674800 953896
rect 675392 953844 675444 953896
rect 674840 952144 674892 952196
rect 674840 952008 674892 952060
rect 675392 952008 675444 952060
rect 675668 951736 675720 951788
rect 674012 951056 674064 951108
rect 675760 951056 675812 951108
rect 673736 950920 673788 950972
rect 674012 950920 674064 950972
rect 673460 950716 673512 950768
rect 673644 950716 673696 950768
rect 35624 949560 35676 949612
rect 43628 949560 43680 949612
rect 35716 949492 35768 949544
rect 42892 949492 42944 949544
rect 41512 949424 41564 949476
rect 58440 949424 58492 949476
rect 41972 943236 42024 943288
rect 62672 943236 62724 943288
rect 41788 943032 41840 943084
rect 49700 943032 49752 943084
rect 703452 942896 703504 942948
rect 709340 942896 709392 942948
rect 41788 942692 41840 942744
rect 48504 942692 48556 942744
rect 41788 941468 41840 941520
rect 46020 941468 46072 941520
rect 41788 941332 41840 941384
rect 42708 941332 42760 941384
rect 41880 941196 41932 941248
rect 42708 941196 42760 941248
rect 703544 940856 703596 940908
rect 708880 940856 708932 940908
rect 708052 940788 708104 940840
rect 704924 940720 704976 940772
rect 707960 940720 708012 940772
rect 704832 940652 704884 940704
rect 707040 940652 707092 940704
rect 706672 940584 706724 940636
rect 705752 940516 705804 940568
rect 706212 940516 706264 940568
rect 706304 940516 706356 940568
rect 706580 940516 706632 940568
rect 705844 940448 705896 940500
rect 707040 940448 707092 940500
rect 707592 940448 707644 940500
rect 705384 940380 705436 940432
rect 707500 940380 707552 940432
rect 705292 940312 705344 940364
rect 708512 940312 708564 940364
rect 704464 940244 704516 940296
rect 708420 940244 708472 940296
rect 704372 940176 704424 940228
rect 655796 938816 655848 938868
rect 676220 938816 676272 938868
rect 655704 938680 655756 938732
rect 676312 938680 676364 938732
rect 655520 938544 655572 938596
rect 676128 938544 676180 938596
rect 49700 938340 49752 938392
rect 58440 938340 58492 938392
rect 41144 936504 41196 936556
rect 41696 936504 41748 936556
rect 670332 935756 670384 935808
rect 676036 935756 676088 935808
rect 670148 935688 670200 935740
rect 676220 935688 676272 935740
rect 649908 935620 649960 935672
rect 678980 935620 679032 935672
rect 674748 935552 674800 935604
rect 676036 935552 676088 935604
rect 674656 935484 674708 935536
rect 676128 935484 676180 935536
rect 674012 935416 674064 935468
rect 675944 935416 675996 935468
rect 673920 935280 673972 935332
rect 675944 935280 675996 935332
rect 674840 934940 674892 934992
rect 676036 934940 676088 934992
rect 673552 933308 673604 933360
rect 676036 933308 676088 933360
rect 674472 932832 674524 932884
rect 676036 932832 676088 932884
rect 673736 932764 673788 932816
rect 676128 932764 676180 932816
rect 673644 932696 673696 932748
rect 675944 932696 675996 932748
rect 674288 932628 674340 932680
rect 676128 932628 676180 932680
rect 41788 932424 41840 932476
rect 46020 932424 46072 932476
rect 673828 932084 673880 932136
rect 675944 932084 675996 932136
rect 674380 931676 674432 931728
rect 676036 931676 676088 931728
rect 674564 931268 674616 931320
rect 676036 931268 676088 931320
rect 672080 927392 672132 927444
rect 678980 927392 679032 927444
rect 654692 922224 654744 922276
rect 669872 922224 669924 922276
rect 48504 921816 48556 921868
rect 58440 921816 58492 921868
rect 53840 908080 53892 908132
rect 58072 908080 58124 908132
rect 654876 908080 654928 908132
rect 663800 908080 663852 908132
rect 53932 896996 53984 897048
rect 58532 896996 58584 897048
rect 654692 895364 654744 895416
rect 660948 895364 661000 895416
rect 51080 883192 51132 883244
rect 58440 883192 58492 883244
rect 673552 873468 673604 873520
rect 675392 873468 675444 873520
rect 674748 872652 674800 872704
rect 675392 872652 675444 872704
rect 655152 870748 655204 870800
rect 674932 870748 674984 870800
rect 673644 869796 673696 869848
rect 675392 869796 675444 869848
rect 656808 869592 656860 869644
rect 663708 869592 663760 869644
rect 50988 869388 51040 869440
rect 58440 869388 58492 869440
rect 674196 868980 674248 869032
rect 675392 868980 675444 869032
rect 673736 868504 673788 868556
rect 675392 868504 675444 868556
rect 674288 867756 674340 867808
rect 675392 867756 675444 867808
rect 673828 866464 673880 866516
rect 675392 866464 675444 866516
rect 674932 866260 674984 866312
rect 675392 866260 675444 866312
rect 674012 864628 674064 864680
rect 675392 864628 675444 864680
rect 673920 862792 673972 862844
rect 675484 862792 675536 862844
rect 48596 858372 48648 858424
rect 58440 858372 58492 858424
rect 655244 855584 655296 855636
rect 666468 855584 666520 855636
rect 674748 854224 674800 854276
rect 675576 854224 675628 854276
rect 48688 844568 48740 844620
rect 58440 844568 58492 844620
rect 654876 841780 654928 841832
rect 667112 841780 667164 841832
rect 54024 830764 54076 830816
rect 57980 830764 58032 830816
rect 41144 819748 41196 819800
rect 62304 819748 62356 819800
rect 41788 817436 41840 817488
rect 53932 817436 53984 817488
rect 41788 817300 41840 817352
rect 51080 817300 51132 817352
rect 53748 817028 53800 817080
rect 59176 817028 59228 817080
rect 42708 816960 42760 817012
rect 62488 816960 62540 817012
rect 655060 815600 655112 815652
rect 668952 815600 669004 815652
rect 41788 814240 41840 814292
rect 42892 814240 42944 814292
rect 62672 814240 62724 814292
rect 41788 810024 41840 810076
rect 43720 810024 43772 810076
rect 41880 807848 41932 807900
rect 43168 807848 43220 807900
rect 41788 807576 41840 807628
rect 42708 807576 42760 807628
rect 41788 806624 41840 806676
rect 46296 806624 46348 806676
rect 51080 805944 51132 805996
rect 58440 805944 58492 805996
rect 656164 803224 656216 803276
rect 661040 803224 661092 803276
rect 44272 800436 44324 800488
rect 48504 800436 48556 800488
rect 41972 800164 42024 800216
rect 41972 799960 42024 800012
rect 43812 799756 43864 799808
rect 44088 799756 44140 799808
rect 42340 799688 42392 799740
rect 43812 799620 43864 799672
rect 42156 798124 42208 798176
rect 42892 798124 42944 798176
rect 42708 797920 42760 797972
rect 43444 797920 43496 797972
rect 42432 797580 42484 797632
rect 42984 797852 43036 797904
rect 43536 797648 43588 797700
rect 43812 798124 43864 798176
rect 43812 797988 43864 798040
rect 44180 797988 44232 798040
rect 42156 797240 42208 797292
rect 44272 797240 44324 797292
rect 42156 796288 42208 796340
rect 42708 796288 42760 796340
rect 674564 796220 674616 796272
rect 675576 796220 675628 796272
rect 42156 794996 42208 795048
rect 43168 794996 43220 795048
rect 42156 794248 42208 794300
rect 43260 794248 43312 794300
rect 42156 793772 42208 793824
rect 42432 793772 42484 793824
rect 42156 792956 42208 793008
rect 43720 792956 43772 793008
rect 51172 792140 51224 792192
rect 58072 792140 58124 792192
rect 42156 790644 42208 790696
rect 43628 790644 43680 790696
rect 42156 790100 42208 790152
rect 43904 790100 43956 790152
rect 655060 789352 655112 789404
rect 663892 789352 663944 789404
rect 42156 789284 42208 789336
rect 43812 789284 43864 789336
rect 42156 788808 42208 788860
rect 43076 788808 43128 788860
rect 42156 786972 42208 787024
rect 43352 786972 43404 787024
rect 42064 786224 42116 786276
rect 44088 786224 44140 786276
rect 42156 785748 42208 785800
rect 42892 785748 42944 785800
rect 674380 784932 674432 784984
rect 675392 784932 675444 784984
rect 673460 782892 673512 782944
rect 675484 782892 675536 782944
rect 655520 782416 655572 782468
rect 674656 782416 674708 782468
rect 674288 780580 674340 780632
rect 675484 780580 675536 780632
rect 674472 779764 674524 779816
rect 675484 779764 675536 779816
rect 674196 779288 674248 779340
rect 675392 779288 675444 779340
rect 674748 778608 674800 778660
rect 675484 778608 675536 778660
rect 48872 778336 48924 778388
rect 58440 778336 58492 778388
rect 674380 777316 674432 777368
rect 675392 777316 675444 777368
rect 674656 777044 674708 777096
rect 675392 777044 675444 777096
rect 674564 775480 674616 775532
rect 675392 775480 675444 775532
rect 41512 774732 41564 774784
rect 48688 774732 48740 774784
rect 41788 774188 41840 774240
rect 54024 774188 54076 774240
rect 41512 773916 41564 773968
rect 48596 773916 48648 773968
rect 674656 773848 674708 773900
rect 675208 773848 675260 773900
rect 41512 773576 41564 773628
rect 43352 773576 43404 773628
rect 43996 773576 44048 773628
rect 674656 773576 674708 773628
rect 675484 773576 675536 773628
rect 674472 773372 674524 773424
rect 675668 773372 675720 773424
rect 675208 773304 675260 773356
rect 675576 773304 675628 773356
rect 674748 773100 674800 773152
rect 675484 773100 675536 773152
rect 42892 772828 42944 772880
rect 62856 772828 62908 772880
rect 674288 770516 674340 770568
rect 674564 770516 674616 770568
rect 673460 770244 673512 770296
rect 674288 770244 674340 770296
rect 48780 767320 48832 767372
rect 58440 767320 58492 767372
rect 43168 766368 43220 766420
rect 43812 766368 43864 766420
rect 41512 763240 41564 763292
rect 48504 763240 48556 763292
rect 708512 762492 708564 762544
rect 704464 762424 704516 762476
rect 708420 762424 708472 762476
rect 704372 762356 704424 762408
rect 707500 762356 707552 762408
rect 707040 762288 707092 762340
rect 705292 762220 705344 762272
rect 705752 762220 705804 762272
rect 706212 762220 706264 762272
rect 706580 762220 706632 762272
rect 705844 762152 705896 762204
rect 707040 762152 707092 762204
rect 706304 762084 706356 762136
rect 706580 762084 706632 762136
rect 705384 762016 705436 762068
rect 707500 762016 707552 762068
rect 708052 762016 708104 762068
rect 704924 761948 704976 762000
rect 707960 761948 708012 762000
rect 704832 761880 704884 761932
rect 708972 761880 709024 761932
rect 703544 761812 703596 761864
rect 708880 761812 708932 761864
rect 654692 761744 654744 761796
rect 667020 761744 667072 761796
rect 704004 761744 704056 761796
rect 41972 760520 42024 760572
rect 50988 760520 51040 760572
rect 669872 759568 669924 759620
rect 676220 759568 676272 759620
rect 663800 759432 663852 759484
rect 678980 759432 679032 759484
rect 660948 759296 661000 759348
rect 676128 759296 676180 759348
rect 673368 759092 673420 759144
rect 676036 759092 676088 759144
rect 670516 759024 670568 759076
rect 676312 759024 676364 759076
rect 674012 758956 674064 759008
rect 676036 758956 676088 759008
rect 42432 757596 42484 757648
rect 42984 757596 43036 757648
rect 43260 757596 43312 757648
rect 43628 757596 43680 757648
rect 42156 757460 42208 757512
rect 43260 757460 43312 757512
rect 42064 757392 42116 757444
rect 42432 757392 42484 757444
rect 41880 756984 41932 757036
rect 41880 756712 41932 756764
rect 42708 756508 42760 756560
rect 44180 756508 44232 756560
rect 670608 756440 670660 756492
rect 676128 756440 676180 756492
rect 668584 756372 668636 756424
rect 676220 756372 676272 756424
rect 669964 756304 670016 756356
rect 670332 756304 670384 756356
rect 676312 756304 676364 756356
rect 669872 756236 669924 756288
rect 670148 756236 670200 756288
rect 678980 756236 679032 756288
rect 673920 756168 673972 756220
rect 676036 756168 676088 756220
rect 673644 756100 673696 756152
rect 676128 756100 676180 756152
rect 42432 755488 42484 755540
rect 42616 755216 42668 755268
rect 42156 754876 42208 754928
rect 43076 754876 43128 754928
rect 673552 754876 673604 754928
rect 676036 754876 676088 754928
rect 43076 754740 43128 754792
rect 43996 754740 44048 754792
rect 44088 754672 44140 754724
rect 44088 754468 44140 754520
rect 53840 753516 53892 753568
rect 58348 753516 58400 753568
rect 673828 753448 673880 753500
rect 676036 753448 676088 753500
rect 673736 753244 673788 753296
rect 676036 753244 676088 753296
rect 42156 753040 42208 753092
rect 43168 753040 43220 753092
rect 42156 751748 42208 751800
rect 42892 751748 42944 751800
rect 42156 751068 42208 751120
rect 43536 751068 43588 751120
rect 42064 750592 42116 750644
rect 43444 750592 43496 750644
rect 43444 750456 43496 750508
rect 44088 750456 44140 750508
rect 672172 749912 672224 749964
rect 679256 749912 679308 749964
rect 42156 749776 42208 749828
rect 43812 749776 43864 749828
rect 43168 749096 43220 749148
rect 43720 749096 43772 749148
rect 42616 748960 42668 749012
rect 43720 748960 43772 749012
rect 654692 748960 654744 749012
rect 668860 748960 668912 749012
rect 42156 746920 42208 746972
rect 43076 746920 43128 746972
rect 42156 746716 42208 746768
rect 43720 746716 43772 746768
rect 42156 746240 42208 746292
rect 43444 746240 43496 746292
rect 42156 745424 42208 745476
rect 43904 745424 43956 745476
rect 42156 743724 42208 743776
rect 44088 743724 44140 743776
rect 42156 743248 42208 743300
rect 43628 743248 43680 743300
rect 42156 742568 42208 742620
rect 43168 742568 43220 742620
rect 48688 739712 48740 739764
rect 58440 739712 58492 739764
rect 673920 738420 673972 738472
rect 674656 738420 674708 738472
rect 655520 738284 655572 738336
rect 674656 738284 674708 738336
rect 654140 736244 654192 736296
rect 661132 736244 661184 736296
rect 674012 735428 674064 735480
rect 675392 735428 675444 735480
rect 673736 734748 673788 734800
rect 675392 734748 675444 734800
rect 673644 734340 673696 734392
rect 675392 734340 675444 734392
rect 673552 733592 673604 733644
rect 675392 733592 675444 733644
rect 673828 732300 673880 732352
rect 675392 732300 675444 732352
rect 674656 732028 674708 732080
rect 675392 732028 675444 732080
rect 674012 731892 674064 731944
rect 674656 731892 674708 731944
rect 41788 731348 41840 731400
rect 51172 731348 51224 731400
rect 41512 731076 41564 731128
rect 48872 731076 48924 731128
rect 41512 730668 41564 730720
rect 51080 730668 51132 730720
rect 41512 730464 41564 730516
rect 43260 730464 43312 730516
rect 673736 730464 673788 730516
rect 675392 730464 675444 730516
rect 42524 729240 42576 729292
rect 42984 729240 43036 729292
rect 674840 728900 674892 728952
rect 675484 728900 675536 728952
rect 41788 728832 41840 728884
rect 44272 728832 44324 728884
rect 42524 728696 42576 728748
rect 63040 728696 63092 728748
rect 51172 725908 51224 725960
rect 58440 725908 58492 725960
rect 673368 723120 673420 723172
rect 678980 723120 679032 723172
rect 673920 722848 673972 722900
rect 675484 722848 675536 722900
rect 674196 721284 674248 721336
rect 674932 721284 674984 721336
rect 674012 721148 674064 721200
rect 674196 721148 674248 721200
rect 703452 720400 703504 720452
rect 709248 720400 709300 720452
rect 41512 719992 41564 720044
rect 48596 719992 48648 720044
rect 41328 717544 41380 717596
rect 43812 717544 43864 717596
rect 704464 717476 704516 717528
rect 708420 717476 708472 717528
rect 708512 717408 708564 717460
rect 704464 717340 704516 717392
rect 705384 717340 705436 717392
rect 707500 717340 707552 717392
rect 707040 717272 707092 717324
rect 705752 717204 705804 717256
rect 706212 717204 706264 717256
rect 706580 717204 706632 717256
rect 705844 717136 705896 717188
rect 707040 717136 707092 717188
rect 707592 717136 707644 717188
rect 706304 717068 706356 717120
rect 706580 717068 706632 717120
rect 705384 717000 705436 717052
rect 708052 717000 708104 717052
rect 704924 716932 704976 716984
rect 707960 716932 708012 716984
rect 704832 716864 704884 716916
rect 703544 716796 703596 716848
rect 708880 716796 708932 716848
rect 42524 716592 42576 716644
rect 53748 716592 53800 716644
rect 666468 716524 666520 716576
rect 676036 716524 676088 716576
rect 663708 716116 663760 716168
rect 676036 716116 676088 716168
rect 667112 715708 667164 715760
rect 676036 715708 676088 715760
rect 670516 715232 670568 715284
rect 676036 715232 676088 715284
rect 670240 714892 670292 714944
rect 676036 714892 676088 714944
rect 50988 714824 51040 714876
rect 58440 714824 58492 714876
rect 670148 714824 670200 714876
rect 670516 714824 670568 714876
rect 673828 714076 673880 714128
rect 675668 714076 675720 714128
rect 673092 714008 673144 714060
rect 676036 714008 676088 714060
rect 41880 713804 41932 713856
rect 670332 713600 670384 713652
rect 670608 713600 670660 713652
rect 676036 713600 676088 713652
rect 41880 713532 41932 713584
rect 669044 713192 669096 713244
rect 670608 713192 670660 713244
rect 676036 713192 676088 713244
rect 668584 712852 668636 712904
rect 676036 712852 676088 712904
rect 669136 712444 669188 712496
rect 670516 712444 670568 712496
rect 676036 712444 676088 712496
rect 674932 712036 674984 712088
rect 676036 712036 676088 712088
rect 674564 711968 674616 712020
rect 675944 711968 675996 712020
rect 674196 711900 674248 711952
rect 675852 711900 675904 711952
rect 42156 711628 42208 711680
rect 43076 711628 43128 711680
rect 43076 711492 43128 711544
rect 43352 711492 43404 711544
rect 42156 711084 42208 711136
rect 42524 711084 42576 711136
rect 673552 710676 673604 710728
rect 674012 710676 674064 710728
rect 674656 710676 674708 710728
rect 675576 710676 675628 710728
rect 673736 710608 673788 710660
rect 674840 710608 674892 710660
rect 674748 710540 674800 710592
rect 676036 710540 676088 710592
rect 42156 709860 42208 709912
rect 42800 709860 42852 709912
rect 42800 709724 42852 709776
rect 43168 709724 43220 709776
rect 655980 709724 656032 709776
rect 660948 709724 661000 709776
rect 43168 709588 43220 709640
rect 43720 709588 43772 709640
rect 674472 709248 674524 709300
rect 676036 709248 676088 709300
rect 42156 708432 42208 708484
rect 43260 708432 43312 708484
rect 674380 708228 674432 708280
rect 676036 708228 676088 708280
rect 42156 708024 42208 708076
rect 43444 708024 43496 708076
rect 674288 707820 674340 707872
rect 676036 707820 676088 707872
rect 676036 707412 676088 707464
rect 676588 707412 676640 707464
rect 42156 707208 42208 707260
rect 44088 707208 44140 707260
rect 42156 706732 42208 706784
rect 43076 706732 43128 706784
rect 671804 705440 671856 705492
rect 675944 705440 675996 705492
rect 42248 704828 42300 704880
rect 42984 704828 43036 704880
rect 42064 704216 42116 704268
rect 43904 704216 43956 704268
rect 42064 702856 42116 702908
rect 43812 702856 43864 702908
rect 42064 702380 42116 702432
rect 43536 702380 43588 702432
rect 53748 701020 53800 701072
rect 58164 701020 58216 701072
rect 42156 700408 42208 700460
rect 43628 700408 43680 700460
rect 42156 700000 42208 700052
rect 42892 700000 42944 700052
rect 670516 699728 670568 699780
rect 674748 699660 674800 699712
rect 675484 699660 675536 699712
rect 674656 699592 674708 699644
rect 675576 699592 675628 699644
rect 670608 699524 670660 699576
rect 42064 699388 42116 699440
rect 42800 699388 42852 699440
rect 654876 696396 654928 696448
rect 663800 696396 663852 696448
rect 655520 691364 655572 691416
rect 674564 691364 674616 691416
rect 673644 690412 673696 690464
rect 675392 690412 675444 690464
rect 673184 689120 673236 689172
rect 675484 689120 675536 689172
rect 673000 688576 673052 688628
rect 675392 688576 675444 688628
rect 41512 688372 41564 688424
rect 48688 688372 48740 688424
rect 41696 687828 41748 687880
rect 53840 687828 53892 687880
rect 41788 687692 41840 687744
rect 51172 687692 51224 687744
rect 673276 687284 673328 687336
rect 675392 687284 675444 687336
rect 51080 687216 51132 687268
rect 58440 687216 58492 687268
rect 674564 687012 674616 687064
rect 675484 687012 675536 687064
rect 674288 685448 674340 685500
rect 675392 685448 675444 685500
rect 42800 684428 42852 684480
rect 62764 684428 62816 684480
rect 673828 683612 673880 683664
rect 675484 683612 675536 683664
rect 654140 683408 654192 683460
rect 669136 683408 669188 683460
rect 673092 678988 673144 679040
rect 678980 678988 679032 679040
rect 41788 678172 41840 678224
rect 43260 678172 43312 678224
rect 41788 677016 41840 677068
rect 48688 677016 48740 677068
rect 48872 673480 48924 673532
rect 58440 673480 58492 673532
rect 41328 673412 41380 673464
rect 43076 673412 43128 673464
rect 703452 672324 703504 672376
rect 703544 672256 703596 672308
rect 708880 672256 708932 672308
rect 708972 672256 709024 672308
rect 708052 672188 708104 672240
rect 704924 672120 704976 672172
rect 707960 672120 708012 672172
rect 704832 672052 704884 672104
rect 707040 672052 707092 672104
rect 706672 671984 706724 672036
rect 705752 671916 705804 671968
rect 706212 671916 706264 671968
rect 706304 671916 706356 671968
rect 706580 671916 706632 671968
rect 705844 671848 705896 671900
rect 707040 671848 707092 671900
rect 707592 671848 707644 671900
rect 705384 671780 705436 671832
rect 707500 671780 707552 671832
rect 705292 671712 705344 671764
rect 708512 671712 708564 671764
rect 704464 671644 704516 671696
rect 708420 671644 708472 671696
rect 704372 671576 704424 671628
rect 674748 671236 674800 671288
rect 675208 671236 675260 671288
rect 668952 670964 669004 671016
rect 676036 670964 676088 671016
rect 661040 670760 661092 670812
rect 676220 670760 676272 670812
rect 44180 670692 44232 670744
rect 48780 670692 48832 670744
rect 44088 670624 44140 670676
rect 41880 670556 41932 670608
rect 41972 670556 42024 670608
rect 42708 670556 42760 670608
rect 41880 670352 41932 670404
rect 663892 670556 663944 670608
rect 676036 670556 676088 670608
rect 670240 670284 670292 670336
rect 676220 670284 676272 670336
rect 44180 670148 44232 670200
rect 674564 668992 674616 669044
rect 676036 668992 676088 669044
rect 670516 668652 670568 668704
rect 676220 668652 676272 668704
rect 42064 668448 42116 668500
rect 43996 668448 44048 668500
rect 673092 668040 673144 668092
rect 675944 668040 675996 668092
rect 674748 667904 674800 667956
rect 676036 667904 676088 667956
rect 673920 667836 673972 667888
rect 676128 667836 676180 667888
rect 674656 667768 674708 667820
rect 676036 667768 676088 667820
rect 42156 667700 42208 667752
rect 44088 667700 44140 667752
rect 670608 667700 670660 667752
rect 675944 667700 675996 667752
rect 42156 666680 42208 666732
rect 43904 666680 43956 666732
rect 42156 665388 42208 665440
rect 42708 665388 42760 665440
rect 675208 665116 675260 665168
rect 676036 665116 676088 665168
rect 673736 665048 673788 665100
rect 676128 665048 676180 665100
rect 42156 664640 42208 664692
rect 43536 664640 43588 664692
rect 42156 664164 42208 664216
rect 43260 664164 43312 664216
rect 42156 663552 42208 663604
rect 43076 663552 43128 663604
rect 48964 662396 49016 662448
rect 58440 662396 58492 662448
rect 42156 661036 42208 661088
rect 44088 661036 44140 661088
rect 42156 660492 42208 660544
rect 43628 660492 43680 660544
rect 42156 659880 42208 659932
rect 43168 659880 43220 659932
rect 672356 659676 672408 659728
rect 678980 659676 679032 659728
rect 42156 658996 42208 659048
rect 43812 658996 43864 659048
rect 42156 657228 42208 657280
rect 43352 657228 43404 657280
rect 656808 657024 656860 657076
rect 663708 657024 663760 657076
rect 42156 656820 42208 656872
rect 43720 656820 43772 656872
rect 42156 656140 42208 656192
rect 42984 656140 43036 656192
rect 674380 649544 674432 649596
rect 675392 649544 675444 649596
rect 53840 648592 53892 648644
rect 59176 648592 59228 648644
rect 673552 647708 673604 647760
rect 675484 647708 675536 647760
rect 674472 647300 674524 647352
rect 674748 647300 674800 647352
rect 655520 647164 655572 647216
rect 674748 647164 674800 647216
rect 673736 645396 673788 645448
rect 675392 645396 675444 645448
rect 41512 645124 41564 645176
rect 51080 645124 51132 645176
rect 41512 644716 41564 644768
rect 48872 644716 48924 644768
rect 41512 644580 41564 644632
rect 53748 644580 53800 644632
rect 674656 644580 674708 644632
rect 675392 644580 675444 644632
rect 673920 644104 673972 644156
rect 675392 644104 675444 644156
rect 41512 643424 41564 643476
rect 44364 643424 44416 643476
rect 674196 643356 674248 643408
rect 675392 643356 675444 643408
rect 42892 643152 42944 643204
rect 62580 643152 62632 643204
rect 654876 643084 654928 643136
rect 666468 643084 666520 643136
rect 674012 642064 674064 642116
rect 675392 642064 675444 642116
rect 674748 641860 674800 641912
rect 675392 641860 675444 641912
rect 674472 641656 674524 641708
rect 674748 641656 674800 641708
rect 674472 640228 674524 640280
rect 675392 640228 675444 640280
rect 674748 638664 674800 638716
rect 675208 638664 675260 638716
rect 674656 638392 674708 638444
rect 675484 638392 675536 638444
rect 674748 638188 674800 638240
rect 675484 638188 675536 638240
rect 674288 638120 674340 638172
rect 674380 638120 674432 638172
rect 675668 638120 675720 638172
rect 674196 637916 674248 637968
rect 673092 637848 673144 637900
rect 679164 637848 679216 637900
rect 675208 637508 675260 637560
rect 679072 637508 679124 637560
rect 674012 637304 674064 637356
rect 674196 637304 674248 637356
rect 673736 637168 673788 637220
rect 674012 637168 674064 637220
rect 48872 634788 48924 634840
rect 58440 634788 58492 634840
rect 41512 633632 41564 633684
rect 48780 633632 48832 633684
rect 43904 629280 43956 629332
rect 50988 629280 51040 629332
rect 654140 629280 654192 629332
rect 667204 629280 667256 629332
rect 33048 627852 33100 627904
rect 42524 627852 42576 627904
rect 41788 627376 41840 627428
rect 708512 627308 708564 627360
rect 704464 627240 704516 627292
rect 708420 627240 708472 627292
rect 704372 627172 704424 627224
rect 41788 627036 41840 627088
rect 705292 627036 705344 627088
rect 707500 627172 707552 627224
rect 707040 627104 707092 627156
rect 705752 627036 705804 627088
rect 706212 627036 706264 627088
rect 706580 627036 706632 627088
rect 705844 626968 705896 627020
rect 707040 626968 707092 627020
rect 706304 626900 706356 626952
rect 706580 626900 706632 626952
rect 705384 626832 705436 626884
rect 707500 626832 707552 626884
rect 708052 626832 708104 626884
rect 704924 626764 704976 626816
rect 707960 626764 708012 626816
rect 704832 626696 704884 626748
rect 708972 626696 709024 626748
rect 703544 626628 703596 626680
rect 708880 626628 708932 626680
rect 704004 626560 704056 626612
rect 42156 625268 42208 625320
rect 43536 625268 43588 625320
rect 42156 624656 42208 624708
rect 43904 624656 43956 624708
rect 670608 624248 670660 624300
rect 674564 624248 674616 624300
rect 676036 624248 676088 624300
rect 668860 624112 668912 624164
rect 678980 624112 679032 624164
rect 667020 623976 667072 624028
rect 676128 623976 676180 624028
rect 673368 623908 673420 623960
rect 676036 623908 676088 623960
rect 661132 623840 661184 623892
rect 676312 623840 676364 623892
rect 51080 623772 51132 623824
rect 58440 623772 58492 623824
rect 670240 623772 670292 623824
rect 670424 623772 670476 623824
rect 676220 623772 676272 623824
rect 674288 623704 674340 623756
rect 676036 623704 676088 623756
rect 42156 623432 42208 623484
rect 42892 623432 42944 623484
rect 42064 622140 42116 622192
rect 42524 622140 42576 622192
rect 42156 621460 42208 621512
rect 43352 621460 43404 621512
rect 670516 621052 670568 621104
rect 676220 621052 676272 621104
rect 42064 620984 42116 621036
rect 43260 620984 43312 621036
rect 670424 620984 670476 621036
rect 678980 620984 679032 621036
rect 673828 620916 673880 620968
rect 676036 620916 676088 620968
rect 673644 620848 673696 620900
rect 676128 620848 676180 620900
rect 42064 620168 42116 620220
rect 43444 620168 43496 620220
rect 42248 619012 42300 619064
rect 43168 619012 43220 619064
rect 673276 618196 673328 618248
rect 676036 618196 676088 618248
rect 673184 617924 673236 617976
rect 676220 617924 676272 617976
rect 42156 617856 42208 617908
rect 43628 617856 43680 617908
rect 42064 617108 42116 617160
rect 43812 617108 43864 617160
rect 673000 616700 673052 616752
rect 676220 616700 676272 616752
rect 42156 616632 42208 616684
rect 43720 616632 43772 616684
rect 672448 614728 672500 614780
rect 679256 614728 679308 614780
rect 42156 614184 42208 614236
rect 43076 614184 43128 614236
rect 42156 613640 42208 613692
rect 42984 613640 43036 613692
rect 42156 612960 42208 613012
rect 42800 612960 42852 613012
rect 50988 609968 51040 610020
rect 58440 609968 58492 610020
rect 674380 608744 674432 608796
rect 675668 608744 675720 608796
rect 654600 603032 654652 603084
rect 674564 603032 674616 603084
rect 654324 602148 654376 602200
rect 661040 602148 661092 602200
rect 41512 601876 41564 601928
rect 48872 601876 48924 601928
rect 41512 601468 41564 601520
rect 51080 601468 51132 601520
rect 674288 600380 674340 600432
rect 675484 600380 675536 600432
rect 41512 599836 41564 599888
rect 44456 599836 44508 599888
rect 674748 599564 674800 599616
rect 675484 599564 675536 599616
rect 673736 599088 673788 599140
rect 675392 599088 675444 599140
rect 41512 598952 41564 599004
rect 43352 598952 43404 599004
rect 673644 598408 673696 598460
rect 675484 598408 675536 598460
rect 673828 597116 673880 597168
rect 675392 597116 675444 597168
rect 674564 596844 674616 596896
rect 675392 596844 675444 596896
rect 674472 596776 674524 596828
rect 674472 596572 674524 596624
rect 53748 596164 53800 596216
rect 59176 596164 59228 596216
rect 674380 595280 674432 595332
rect 675392 595280 675444 595332
rect 675208 593648 675260 593700
rect 675484 593648 675536 593700
rect 674564 593036 674616 593088
rect 675576 593036 675628 593088
rect 43444 592560 43496 592612
rect 43996 592560 44048 592612
rect 43260 592424 43312 592476
rect 43444 592424 43496 592476
rect 656808 590656 656860 590708
rect 669044 590656 669096 590708
rect 673368 587868 673420 587920
rect 678980 587868 679032 587920
rect 41328 585148 41380 585200
rect 44088 585148 44140 585200
rect 44180 585148 44232 585200
rect 48964 585148 49016 585200
rect 41880 584196 41932 584248
rect 703452 584128 703504 584180
rect 709340 584128 709392 584180
rect 41880 583924 41932 583976
rect 674380 583924 674432 583976
rect 674564 583924 674616 583976
rect 674656 583924 674708 583976
rect 675392 583924 675444 583976
rect 43168 583856 43220 583908
rect 43444 583856 43496 583908
rect 673828 583856 673880 583908
rect 673644 583720 673696 583772
rect 673828 583720 673880 583772
rect 674748 583720 674800 583772
rect 675484 583720 675536 583772
rect 42432 583652 42484 583704
rect 43260 583652 43312 583704
rect 674380 583652 674432 583704
rect 674564 583652 674616 583704
rect 675208 583652 675260 583704
rect 48964 582360 49016 582412
rect 58440 582360 58492 582412
rect 42156 582088 42208 582140
rect 42892 582088 42944 582140
rect 704004 582088 704056 582140
rect 708880 582088 708932 582140
rect 708052 582020 708104 582072
rect 704924 581952 704976 582004
rect 707960 581952 708012 582004
rect 704832 581884 704884 581936
rect 707040 581884 707092 581936
rect 706672 581816 706724 581868
rect 705752 581748 705804 581800
rect 706212 581748 706264 581800
rect 706304 581748 706356 581800
rect 706580 581748 706632 581800
rect 705844 581680 705896 581732
rect 707040 581680 707092 581732
rect 707592 581680 707644 581732
rect 705384 581612 705436 581664
rect 707500 581612 707552 581664
rect 705292 581544 705344 581596
rect 708512 581544 708564 581596
rect 704464 581476 704516 581528
rect 708420 581476 708472 581528
rect 704372 581408 704424 581460
rect 42156 581272 42208 581324
rect 44180 581272 44232 581324
rect 42156 580252 42208 580304
rect 42800 580252 42852 580304
rect 670240 580184 670292 580236
rect 676036 580184 676088 580236
rect 669136 580048 669188 580100
rect 676220 580048 676272 580100
rect 663800 579912 663852 579964
rect 676128 579912 676180 579964
rect 660948 579776 661000 579828
rect 676312 579776 676364 579828
rect 672540 579232 672592 579284
rect 673276 579232 673328 579284
rect 676220 579232 676272 579284
rect 42156 578960 42208 579012
rect 42708 578960 42760 579012
rect 42156 578416 42208 578468
rect 43628 578416 43680 578468
rect 673092 578416 673144 578468
rect 676220 578416 676272 578468
rect 42156 577804 42208 577856
rect 43168 577804 43220 577856
rect 672724 577600 672776 577652
rect 673184 577600 673236 577652
rect 676220 577600 676272 577652
rect 670516 577124 670568 577176
rect 676220 577124 676272 577176
rect 42156 576920 42208 576972
rect 43996 576920 44048 576972
rect 673368 576920 673420 576972
rect 676036 576920 676088 576972
rect 654508 576852 654560 576904
rect 663892 576852 663944 576904
rect 674472 576784 674524 576836
rect 676036 576784 676088 576836
rect 674012 576036 674064 576088
rect 676036 576036 676088 576088
rect 42156 574676 42208 574728
rect 43720 574676 43772 574728
rect 42156 574064 42208 574116
rect 42984 574064 43036 574116
rect 674196 573588 674248 573640
rect 676036 573588 676088 573640
rect 42156 573452 42208 573504
rect 44088 573452 44140 573504
rect 42064 572840 42116 572892
rect 43904 572840 43956 572892
rect 673920 572772 673972 572824
rect 676036 572772 676088 572824
rect 673552 572364 673604 572416
rect 676036 572364 676088 572416
rect 42064 570868 42116 570920
rect 43812 570868 43864 570920
rect 42156 570392 42208 570444
rect 43444 570392 43496 570444
rect 42064 569576 42116 569628
rect 43536 569576 43588 569628
rect 672540 568556 672592 568608
rect 678980 568556 679032 568608
rect 673552 559512 673604 559564
rect 675484 559512 675536 559564
rect 41512 558764 41564 558816
rect 48964 558764 49016 558816
rect 41512 558288 41564 558340
rect 53748 558288 53800 558340
rect 41788 558220 41840 558272
rect 58440 558220 58492 558272
rect 49056 557540 49108 557592
rect 57980 557540 58032 557592
rect 654324 556112 654376 556164
rect 675300 556112 675352 556164
rect 674196 555228 674248 555280
rect 675392 555228 675444 555280
rect 673460 554548 673512 554600
rect 675392 554548 675444 554600
rect 673920 553732 673972 553784
rect 675392 553732 675444 553784
rect 673644 553188 673696 553240
rect 675392 553188 675444 553240
rect 674012 551896 674064 551948
rect 675392 551896 675444 551948
rect 655060 550196 655112 550248
rect 669136 550196 669188 550248
rect 674472 548836 674524 548888
rect 675300 548836 675352 548888
rect 674656 548224 674708 548276
rect 675300 548224 675352 548276
rect 41420 547272 41472 547324
rect 48964 547272 49016 547324
rect 673092 546252 673144 546304
rect 679072 546252 679124 546304
rect 53840 543736 53892 543788
rect 59176 543736 59228 543788
rect 41604 543124 41656 543176
rect 43260 543124 43312 543176
rect 41512 542444 41564 542496
rect 42800 542444 42852 542496
rect 41788 541016 41840 541068
rect 43904 541016 43956 541068
rect 50988 541016 51040 541068
rect 41788 540744 41840 540796
rect 42064 538908 42116 538960
rect 42708 538908 42760 538960
rect 42156 538092 42208 538144
rect 43904 538092 43956 538144
rect 703452 537140 703504 537192
rect 42064 537072 42116 537124
rect 42892 537072 42944 537124
rect 703544 537072 703596 537124
rect 708880 537072 708932 537124
rect 708972 537072 709024 537124
rect 708052 537004 708104 537056
rect 704924 536936 704976 536988
rect 707960 536936 708012 536988
rect 42984 536868 43036 536920
rect 43352 536868 43404 536920
rect 704832 536868 704884 536920
rect 707040 536868 707092 536920
rect 706672 536800 706724 536852
rect 43352 536732 43404 536784
rect 43536 536732 43588 536784
rect 705752 536732 705804 536784
rect 706212 536732 706264 536784
rect 706304 536732 706356 536784
rect 706580 536732 706632 536784
rect 705844 536664 705896 536716
rect 707040 536664 707092 536716
rect 707592 536664 707644 536716
rect 705384 536596 705436 536648
rect 707500 536596 707552 536648
rect 705292 536528 705344 536580
rect 708512 536528 708564 536580
rect 704464 536460 704516 536512
rect 708420 536460 708472 536512
rect 654692 536392 654744 536444
rect 667112 536392 667164 536444
rect 704372 536392 704424 536444
rect 42156 535780 42208 535832
rect 42800 535780 42852 535832
rect 666468 535712 666520 535764
rect 676220 535712 676272 535764
rect 663708 535576 663760 535628
rect 676036 535576 676088 535628
rect 42064 535032 42116 535084
rect 43444 535032 43496 535084
rect 673276 534896 673328 534948
rect 676036 534896 676088 534948
rect 42156 534556 42208 534608
rect 43260 534556 43312 534608
rect 42156 533740 42208 533792
rect 43168 533740 43220 533792
rect 673184 533264 673236 533316
rect 676036 533264 676088 533316
rect 667204 532856 667256 532908
rect 678980 532856 679032 532908
rect 670056 532788 670108 532840
rect 675852 532788 675904 532840
rect 676128 532788 676180 532840
rect 674748 532652 674800 532704
rect 676036 532652 676088 532704
rect 672816 532584 672868 532636
rect 673368 532584 673420 532636
rect 676220 532584 676272 532636
rect 42156 531428 42208 531480
rect 43812 531428 43864 531480
rect 674288 531088 674340 531140
rect 676036 531088 676088 531140
rect 42156 530680 42208 530732
rect 43720 530680 43772 530732
rect 42156 530272 42208 530324
rect 43076 530272 43128 530324
rect 674564 529864 674616 529916
rect 676036 529864 676088 529916
rect 42156 529592 42208 529644
rect 42892 529592 42944 529644
rect 674380 529456 674432 529508
rect 676036 529456 676088 529508
rect 673736 527824 673788 527876
rect 676036 527824 676088 527876
rect 42064 527212 42116 527264
rect 43352 527212 43404 527264
rect 42156 527144 42208 527196
rect 43628 527144 43680 527196
rect 673828 527076 673880 527128
rect 676036 527076 676088 527128
rect 42156 526600 42208 526652
rect 42984 526600 43036 526652
rect 672632 524424 672684 524476
rect 678980 524424 679032 524476
rect 677508 524356 677560 524408
rect 679072 524356 679124 524408
rect 654140 522452 654192 522504
rect 661224 522452 661276 522504
rect 51264 518916 51316 518968
rect 58440 518916 58492 518968
rect 654784 510620 654836 510672
rect 667020 510620 667072 510672
rect 50988 505112 51040 505164
rect 58440 505112 58492 505164
rect 656808 497632 656860 497684
rect 663800 497632 663852 497684
rect 704372 493076 704424 493128
rect 704464 493008 704516 493060
rect 708420 493008 708472 493060
rect 705384 492940 705436 492992
rect 707040 492872 707092 492924
rect 705752 492804 705804 492856
rect 706212 492804 706264 492856
rect 706580 492804 706632 492856
rect 708512 492940 708564 492992
rect 707592 492804 707644 492856
rect 705844 492736 705896 492788
rect 707040 492736 707092 492788
rect 706304 492668 706356 492720
rect 706580 492668 706632 492720
rect 705384 492600 705436 492652
rect 707500 492600 707552 492652
rect 704832 492532 704884 492584
rect 707960 492532 708012 492584
rect 703912 492464 703964 492516
rect 708880 492464 708932 492516
rect 704924 492396 704976 492448
rect 707960 492396 708012 492448
rect 703544 492328 703596 492380
rect 708880 492328 708932 492380
rect 669044 491648 669096 491700
rect 676036 491648 676088 491700
rect 663892 491512 663944 491564
rect 676036 491512 676088 491564
rect 661040 491376 661092 491428
rect 675944 491376 675996 491428
rect 49148 491308 49200 491360
rect 57980 491308 58032 491360
rect 676220 491240 676272 491292
rect 677508 491240 677560 491292
rect 676128 490152 676180 490204
rect 676036 489948 676088 490000
rect 669596 488520 669648 488572
rect 675576 488520 675628 488572
rect 675944 488520 675996 488572
rect 669688 488044 669740 488096
rect 675208 488044 675260 488096
rect 674472 487840 674524 487892
rect 676036 487840 676088 487892
rect 673552 487432 673604 487484
rect 675944 487432 675996 487484
rect 674196 487092 674248 487144
rect 676036 487092 676088 487144
rect 674656 485732 674708 485784
rect 676036 485732 676088 485784
rect 674012 485460 674064 485512
rect 676036 485460 676088 485512
rect 673920 483828 673972 483880
rect 676036 483828 676088 483880
rect 655060 483284 655112 483336
rect 670056 483284 670108 483336
rect 673644 482944 673696 482996
rect 676036 482944 676088 482996
rect 673460 482876 673512 482928
rect 675944 482876 675996 482928
rect 672724 481040 672776 481092
rect 676036 481108 676088 481160
rect 51172 480224 51224 480276
rect 58440 480224 58492 480276
rect 675576 478864 675628 478916
rect 676128 478864 676180 478916
rect 654876 470500 654928 470552
rect 663708 470500 663760 470552
rect 54024 466420 54076 466472
rect 58624 466420 58676 466472
rect 654140 457308 654192 457360
rect 661040 457308 661092 457360
rect 53748 452616 53800 452668
rect 59176 452616 59228 452668
rect 656808 444456 656860 444508
rect 663892 444456 663944 444508
rect 51080 438880 51132 438932
rect 58440 438880 58492 438932
rect 43996 430652 44048 430704
rect 62396 430652 62448 430704
rect 41788 430584 41840 430636
rect 59268 430584 59320 430636
rect 654876 430584 654928 430636
rect 666468 430584 666520 430636
rect 53932 427864 53984 427916
rect 57980 427864 58032 427916
rect 41788 427796 41840 427848
rect 44088 427796 44140 427848
rect 62948 427796 63000 427848
rect 655060 417460 655112 417512
rect 660948 417460 661000 417512
rect 41788 416304 41840 416356
rect 43076 416304 43128 416356
rect 49240 413992 49292 414044
rect 58440 413992 58492 414044
rect 41880 413380 41932 413432
rect 41880 413108 41932 413160
rect 42800 411340 42852 411392
rect 42156 411272 42208 411324
rect 42156 410660 42208 410712
rect 49056 410660 49108 410712
rect 42156 409368 42208 409420
rect 42984 409368 43036 409420
rect 42064 408144 42116 408196
rect 42524 408144 42576 408196
rect 42156 407464 42208 407516
rect 43352 407464 43404 407516
rect 42064 406988 42116 407040
rect 43076 406988 43128 407040
rect 42156 406172 42208 406224
rect 43444 406172 43496 406224
rect 703544 404880 703596 404932
rect 704004 404880 704056 404932
rect 708880 404880 708932 404932
rect 708972 404880 709024 404932
rect 708052 404812 708104 404864
rect 704924 404744 704976 404796
rect 707960 404744 708012 404796
rect 704832 404676 704884 404728
rect 705752 404540 705804 404592
rect 707040 404676 707092 404728
rect 706672 404608 706724 404660
rect 706212 404540 706264 404592
rect 706304 404540 706356 404592
rect 706580 404540 706632 404592
rect 705844 404472 705896 404524
rect 707040 404472 707092 404524
rect 707592 404472 707644 404524
rect 705384 404404 705436 404456
rect 707500 404404 707552 404456
rect 705292 404336 705344 404388
rect 708512 404336 708564 404388
rect 704464 404268 704516 404320
rect 708420 404268 708472 404320
rect 704372 404200 704424 404252
rect 654876 403996 654928 404048
rect 661132 403996 661184 404048
rect 42156 403860 42208 403912
rect 43996 403860 44048 403912
rect 669136 403384 669188 403436
rect 675944 403384 675996 403436
rect 42156 403316 42208 403368
rect 43628 403316 43680 403368
rect 667112 403248 667164 403300
rect 676220 403248 676272 403300
rect 661224 403112 661276 403164
rect 675944 403112 675996 403164
rect 42156 402500 42208 402552
rect 43812 402500 43864 402552
rect 42156 402024 42208 402076
rect 43168 402024 43220 402076
rect 674656 401208 674708 401260
rect 676128 401208 676180 401260
rect 49056 400188 49108 400240
rect 58440 400188 58492 400240
rect 42156 399984 42208 400036
rect 43260 399984 43312 400036
rect 42156 399440 42208 399492
rect 43812 399440 43864 399492
rect 674380 399440 674432 399492
rect 676036 399440 676088 399492
rect 42156 398964 42208 399016
rect 42892 398964 42944 399016
rect 674472 398216 674524 398268
rect 676036 398216 676088 398268
rect 673736 397604 673788 397656
rect 675944 397604 675996 397656
rect 674288 397536 674340 397588
rect 676128 397536 676180 397588
rect 674932 397468 674984 397520
rect 676036 397468 676088 397520
rect 673460 396584 673512 396636
rect 676036 396584 676088 396636
rect 673552 395360 673604 395412
rect 675944 395360 675996 395412
rect 675116 394952 675168 395004
rect 676036 394952 676088 395004
rect 673644 394816 673696 394868
rect 675944 394816 675996 394868
rect 675024 394748 675076 394800
rect 676128 394748 676180 394800
rect 675208 394680 675260 394732
rect 676036 394680 676088 394732
rect 673828 394136 673880 394188
rect 676036 394136 676088 394188
rect 672908 392028 672960 392080
rect 678980 392028 679032 392080
rect 674012 391960 674064 392012
rect 676036 391960 676088 392012
rect 674748 390532 674800 390584
rect 675760 390532 675812 390584
rect 674564 390464 674616 390516
rect 675668 390464 675720 390516
rect 654140 389784 654192 389836
rect 669596 389784 669648 389836
rect 53840 389172 53892 389224
rect 57980 389172 58032 389224
rect 41512 387948 41564 388000
rect 51172 387948 51224 388000
rect 41788 387404 41840 387456
rect 54024 387404 54076 387456
rect 41512 387132 41564 387184
rect 49148 387132 49200 387184
rect 42800 386384 42852 386436
rect 63132 386384 63184 386436
rect 675760 386384 675812 386436
rect 675760 386112 675812 386164
rect 674472 384956 674524 385008
rect 675300 384956 675352 385008
rect 675208 384072 675260 384124
rect 675300 383868 675352 383920
rect 674932 383120 674984 383172
rect 675392 383120 675444 383172
rect 675116 382440 675168 382492
rect 675392 382440 675444 382492
rect 674380 382304 674432 382356
rect 675116 382304 675168 382356
rect 675024 381896 675076 381948
rect 675392 381896 675444 381948
rect 673736 379448 673788 379500
rect 675300 379448 675352 379500
rect 656808 378156 656860 378208
rect 669688 378156 669740 378208
rect 673644 378156 673696 378208
rect 675300 378156 675352 378208
rect 673828 377952 673880 378004
rect 675484 377952 675536 378004
rect 674012 376932 674064 376984
rect 675484 376932 675536 376984
rect 673552 376864 673604 376916
rect 675300 376864 675352 376916
rect 41420 376456 41472 376508
rect 46756 376456 46808 376508
rect 49148 375368 49200 375420
rect 58440 375368 58492 375420
rect 675116 374076 675168 374128
rect 675300 374076 675352 374128
rect 674288 373872 674340 373924
rect 675392 373872 675444 373924
rect 675300 372852 675352 372904
rect 675300 372648 675352 372700
rect 673460 372036 673512 372088
rect 675392 372036 675444 372088
rect 42800 371764 42852 371816
rect 43352 371764 43404 371816
rect 41512 371424 41564 371476
rect 42800 371424 42852 371476
rect 674748 370744 674800 370796
rect 675760 370744 675812 370796
rect 674564 370676 674616 370728
rect 675668 370676 675720 370728
rect 42156 369928 42208 369980
rect 42340 369928 42392 369980
rect 42156 368092 42208 368144
rect 42708 368092 42760 368144
rect 42156 366800 42208 366852
rect 50988 366800 51040 366852
rect 42156 366256 42208 366308
rect 43076 366256 43128 366308
rect 42156 364964 42208 365016
rect 42800 364964 42852 365016
rect 42156 364420 42208 364472
rect 43260 364420 43312 364472
rect 656808 364352 656860 364404
rect 667112 364352 667164 364404
rect 42156 363808 42208 363860
rect 43168 363808 43220 363860
rect 42156 363128 42208 363180
rect 43352 363128 43404 363180
rect 43168 362788 43220 362840
rect 43628 362788 43680 362840
rect 703452 361700 703504 361752
rect 709340 361700 709392 361752
rect 51172 361564 51224 361616
rect 58440 361564 58492 361616
rect 42064 360680 42116 360732
rect 43076 360680 43128 360732
rect 42156 359932 42208 359984
rect 43812 359932 43864 359984
rect 708512 359660 708564 359712
rect 704464 359592 704516 359644
rect 708420 359592 708472 359644
rect 704372 359524 704424 359576
rect 42156 359456 42208 359508
rect 43628 359456 43680 359508
rect 707500 359524 707552 359576
rect 707040 359456 707092 359508
rect 705292 359388 705344 359440
rect 705752 359388 705804 359440
rect 706212 359388 706264 359440
rect 706580 359388 706632 359440
rect 705844 359320 705896 359372
rect 707040 359320 707092 359372
rect 706304 359252 706356 359304
rect 706580 359252 706632 359304
rect 705384 359184 705436 359236
rect 707500 359184 707552 359236
rect 708052 359184 708104 359236
rect 704924 359116 704976 359168
rect 707960 359116 708012 359168
rect 704832 359048 704884 359100
rect 703820 358844 703872 358896
rect 708880 358844 708932 358896
rect 42064 358776 42116 358828
rect 42892 358776 42944 358828
rect 673276 357008 673328 357060
rect 675576 357008 675628 357060
rect 42064 356940 42116 356992
rect 42984 356940 43036 356992
rect 670056 356464 670108 356516
rect 676036 356464 676088 356516
rect 667020 356328 667072 356380
rect 675944 356328 675996 356380
rect 42156 356260 42208 356312
rect 43168 356260 43220 356312
rect 663800 356192 663852 356244
rect 675852 356192 675904 356244
rect 673368 356124 673420 356176
rect 676036 356124 676088 356176
rect 669504 356056 669556 356108
rect 673000 356056 673052 356108
rect 673276 356056 673328 356108
rect 673184 355376 673236 355428
rect 676036 355376 676088 355428
rect 673276 354560 673328 354612
rect 676036 354560 676088 354612
rect 669412 353472 669464 353524
rect 673092 353472 673144 353524
rect 673276 353472 673328 353524
rect 673552 353472 673604 353524
rect 676036 353472 676088 353524
rect 669320 353336 669372 353388
rect 673184 353336 673236 353388
rect 674012 353268 674064 353320
rect 676036 353268 676088 353320
rect 674564 351432 674616 351484
rect 676036 351432 676088 351484
rect 673460 351024 673512 351076
rect 675944 351024 675996 351076
rect 674656 350616 674708 350668
rect 675944 350616 675996 350668
rect 654876 350548 654928 350600
rect 669412 350548 669464 350600
rect 674748 350548 674800 350600
rect 676036 350548 676088 350600
rect 673736 349800 673788 349852
rect 676036 349800 676088 349852
rect 673828 347896 673880 347948
rect 675852 347896 675904 347948
rect 673920 347828 673972 347880
rect 675944 347828 675996 347880
rect 50988 347760 51040 347812
rect 58440 347760 58492 347812
rect 674840 347760 674892 347812
rect 676036 347760 676088 347812
rect 44364 344972 44416 345024
rect 48412 344972 48464 345024
rect 41512 344224 41564 344276
rect 53932 344224 53984 344276
rect 41788 344156 41840 344208
rect 49240 344156 49292 344208
rect 41512 344088 41564 344140
rect 43536 344088 43588 344140
rect 41604 343884 41656 343936
rect 51080 343884 51132 343936
rect 41788 343340 41840 343392
rect 44364 343340 44416 343392
rect 673000 342388 673052 342440
rect 675760 342388 675812 342440
rect 674012 340960 674064 341012
rect 675484 340960 675536 341012
rect 673552 339736 673604 339788
rect 675484 339736 675536 339788
rect 674564 337900 674616 337952
rect 675484 337900 675536 337952
rect 674748 337016 674800 337068
rect 675392 337016 675444 337068
rect 654324 336812 654376 336864
rect 667020 336812 667072 336864
rect 48412 336744 48464 336796
rect 58440 336744 58492 336796
rect 674656 336540 674708 336592
rect 675392 336540 675444 336592
rect 674840 336064 674892 336116
rect 675484 336064 675536 336116
rect 673460 333548 673512 333600
rect 675392 333548 675444 333600
rect 41512 333208 41564 333260
rect 46204 333208 46256 333260
rect 673920 332936 673972 332988
rect 675392 332936 675444 332988
rect 673736 332188 673788 332240
rect 675392 332188 675444 332240
rect 673828 331576 673880 331628
rect 675392 331576 675444 331628
rect 33048 330080 33100 330132
rect 41880 330080 41932 330132
rect 32956 329944 33008 329996
rect 42892 329944 42944 329996
rect 32680 329876 32732 329928
rect 42800 329876 42852 329928
rect 32864 329808 32916 329860
rect 43352 329808 43404 329860
rect 41880 326952 41932 327004
rect 41880 326748 41932 326800
rect 42064 324912 42116 324964
rect 42800 324912 42852 324964
rect 42800 324776 42852 324828
rect 43076 324776 43128 324828
rect 654324 323892 654376 323944
rect 669136 323892 669188 323944
rect 53932 323484 53984 323536
rect 58164 323484 58216 323536
rect 42156 323280 42208 323332
rect 42616 323280 42668 323332
rect 42064 323076 42116 323128
rect 42892 323076 42944 323128
rect 42156 321784 42208 321836
rect 43168 321784 43220 321836
rect 42156 321036 42208 321088
rect 43352 321036 43404 321088
rect 42156 320560 42208 320612
rect 42984 320560 43036 320612
rect 42616 320084 42668 320136
rect 53748 320084 53800 320136
rect 42156 317432 42208 317484
rect 42800 317432 42852 317484
rect 704004 314712 704056 314764
rect 708880 314712 708932 314764
rect 658464 314576 658516 314628
rect 671160 314576 671212 314628
rect 708512 314644 708564 314696
rect 704464 314576 704516 314628
rect 708420 314576 708472 314628
rect 704372 314508 704424 314560
rect 707500 314508 707552 314560
rect 707040 314440 707092 314492
rect 705292 314372 705344 314424
rect 705752 314372 705804 314424
rect 706212 314372 706264 314424
rect 706580 314372 706632 314424
rect 705844 314304 705896 314356
rect 707040 314304 707092 314356
rect 706304 314236 706356 314288
rect 706580 314236 706632 314288
rect 705384 314168 705436 314220
rect 707500 314168 707552 314220
rect 708052 314168 708104 314220
rect 704924 314100 704976 314152
rect 707960 314100 708012 314152
rect 704832 314032 704884 314084
rect 703544 313964 703596 314016
rect 708880 313964 708932 314016
rect 663708 313284 663760 313336
rect 676036 313284 676088 313336
rect 663892 312876 663944 312928
rect 676036 312876 676088 312928
rect 673184 312468 673236 312520
rect 676036 312468 676088 312520
rect 671160 312060 671212 312112
rect 672264 312060 672316 312112
rect 676036 312060 676088 312112
rect 661040 311992 661092 312044
rect 676220 311992 676272 312044
rect 658372 311788 658424 311840
rect 671160 311788 671212 311840
rect 654140 311652 654192 311704
rect 669320 311652 669372 311704
rect 673368 311652 673420 311704
rect 676036 311652 676088 311704
rect 674748 310972 674800 311024
rect 676036 310972 676088 311024
rect 673276 310836 673328 310888
rect 676036 310836 676088 310888
rect 655428 310428 655480 310480
rect 671896 310428 671948 310480
rect 676036 310428 676088 310480
rect 673092 310020 673144 310072
rect 676036 310020 676088 310072
rect 671160 309612 671212 309664
rect 673184 309612 673236 309664
rect 676036 309612 676088 309664
rect 674196 309136 674248 309188
rect 676036 309136 676088 309188
rect 673552 308048 673604 308100
rect 676036 308048 676088 308100
rect 674472 306824 674524 306876
rect 676036 306824 676088 306876
rect 673460 306484 673512 306536
rect 675944 306484 675996 306536
rect 673920 306416 673972 306468
rect 676128 306416 676180 306468
rect 676036 306348 676088 306400
rect 675116 306212 675168 306264
rect 673736 305056 673788 305108
rect 676128 305056 676180 305108
rect 674656 304784 674708 304836
rect 676036 304784 676088 304836
rect 673828 304240 673880 304292
rect 676128 304240 676180 304292
rect 673644 303764 673696 303816
rect 675944 303764 675996 303816
rect 674012 303696 674064 303748
rect 676128 303696 676180 303748
rect 674564 303628 674616 303680
rect 676036 303628 676088 303680
rect 41512 301588 41564 301640
rect 49148 301588 49200 301640
rect 41788 300908 41840 300960
rect 51172 300908 51224 300960
rect 673092 300840 673144 300892
rect 679072 300840 679124 300892
rect 656808 298392 656860 298444
rect 669504 298392 669556 298444
rect 675760 296148 675812 296200
rect 675760 295944 675812 295996
rect 675208 295060 675260 295112
rect 675392 295060 675444 295112
rect 674196 294516 674248 294568
rect 675392 294516 675444 294568
rect 674472 292884 674524 292936
rect 675392 292884 675444 292936
rect 674656 291524 674708 291576
rect 675392 291524 675444 291576
rect 674564 291048 674616 291100
rect 675392 291048 675444 291100
rect 673920 288532 673972 288584
rect 675392 288532 675444 288584
rect 674012 287920 674064 287972
rect 675392 287920 675444 287972
rect 673828 287172 673880 287224
rect 675484 287172 675536 287224
rect 35808 286968 35860 287020
rect 42708 286968 42760 287020
rect 673644 286560 673696 286612
rect 675392 286560 675444 286612
rect 32864 285744 32916 285796
rect 42800 285744 42852 285796
rect 32956 285676 33008 285728
rect 43260 285676 43312 285728
rect 32680 285608 32732 285660
rect 41880 285608 41932 285660
rect 673736 285540 673788 285592
rect 675484 285540 675536 285592
rect 655704 284724 655756 284776
rect 670056 284724 670108 284776
rect 41880 283772 41932 283824
rect 673552 283704 673604 283756
rect 675484 283704 675536 283756
rect 41880 283568 41932 283620
rect 673460 281868 673512 281920
rect 675392 281868 675444 281920
rect 42156 281732 42208 281784
rect 42708 281732 42760 281784
rect 42156 281052 42208 281104
rect 49056 281052 49108 281104
rect 42156 279828 42208 279880
rect 42984 279828 43036 279880
rect 42064 278604 42116 278656
rect 43352 278604 43404 278656
rect 46480 278536 46532 278588
rect 670608 278536 670660 278588
rect 46572 278468 46624 278520
rect 670424 278468 670476 278520
rect 62580 278400 62632 278452
rect 670516 278400 670568 278452
rect 62028 278332 62080 278384
rect 669872 278332 669924 278384
rect 62396 278264 62448 278316
rect 670148 278264 670200 278316
rect 62764 278196 62816 278248
rect 670332 278196 670384 278248
rect 62948 278128 63000 278180
rect 668584 278128 668636 278180
rect 63316 278060 63368 278112
rect 669964 278060 670016 278112
rect 42156 277992 42208 278044
rect 43168 277992 43220 278044
rect 63132 277992 63184 278044
rect 669780 277992 669832 278044
rect 42156 277380 42208 277432
rect 43628 277380 43680 277432
rect 42064 276700 42116 276752
rect 42800 276700 42852 276752
rect 345112 275952 345164 276004
rect 471336 275952 471388 276004
rect 343732 275884 343784 275936
rect 467840 275884 467892 275936
rect 349068 275816 349120 275868
rect 482008 275816 482060 275868
rect 350172 275748 350224 275800
rect 485504 275748 485556 275800
rect 354404 275680 354456 275732
rect 496176 275680 496228 275732
rect 355784 275612 355836 275664
rect 499764 275612 499816 275664
rect 358452 275544 358504 275596
rect 506848 275544 506900 275596
rect 361120 275476 361172 275528
rect 513932 275476 513984 275528
rect 364064 275408 364116 275460
rect 521016 275408 521068 275460
rect 366456 275340 366508 275392
rect 528100 275340 528152 275392
rect 369124 275272 369176 275324
rect 535184 275272 535236 275324
rect 371792 275204 371844 275256
rect 542268 275204 542320 275256
rect 374920 275136 374972 275188
rect 550548 275136 550600 275188
rect 377588 275068 377640 275120
rect 557632 275068 557684 275120
rect 380256 275000 380308 275052
rect 564716 275000 564768 275052
rect 382924 274932 382976 274984
rect 571800 274932 571852 274984
rect 385592 274864 385644 274916
rect 578884 274864 578936 274916
rect 318892 274796 318944 274848
rect 401600 274796 401652 274848
rect 403900 274796 403952 274848
rect 320180 274728 320232 274780
rect 405188 274728 405240 274780
rect 406568 274728 406620 274780
rect 420920 274796 420972 274848
rect 620284 274796 620336 274848
rect 321008 274660 321060 274712
rect 407488 274660 407540 274712
rect 409236 274660 409288 274712
rect 627368 274728 627420 274780
rect 322756 274592 322808 274644
rect 411076 274592 411128 274644
rect 634452 274660 634504 274712
rect 641628 274592 641680 274644
rect 342536 274524 342588 274576
rect 464252 274524 464304 274576
rect 341064 274456 341116 274508
rect 460664 274456 460716 274508
rect 337108 274388 337160 274440
rect 450084 274388 450136 274440
rect 336096 274320 336148 274372
rect 446496 274320 446548 274372
rect 42156 274252 42208 274304
rect 43076 274252 43128 274304
rect 333152 274252 333204 274304
rect 439412 274252 439464 274304
rect 334348 274184 334400 274236
rect 443000 274184 443052 274236
rect 332140 274116 332192 274168
rect 437020 274116 437072 274168
rect 351828 274048 351880 274100
rect 432328 274048 432380 274100
rect 331680 273980 331732 274032
rect 435916 273980 435968 274032
rect 327724 273912 327776 273964
rect 425244 273912 425296 273964
rect 329012 273844 329064 273896
rect 428832 273844 428884 273896
rect 326804 273776 326856 273828
rect 422852 273776 422904 273828
rect 42064 273708 42116 273760
rect 42892 273708 42944 273760
rect 325424 273708 325476 273760
rect 418160 273708 418212 273760
rect 326344 273640 326396 273692
rect 323676 273572 323728 273624
rect 330392 273504 330444 273556
rect 351828 273504 351880 273556
rect 421656 273572 421708 273624
rect 414572 273504 414624 273556
rect 401140 273436 401192 273488
rect 420920 273436 420972 273488
rect 155684 273096 155736 273148
rect 226156 273164 226208 273216
rect 263232 273164 263284 273216
rect 266728 273164 266780 273216
rect 292028 273164 292080 273216
rect 329472 273164 329524 273216
rect 339500 273164 339552 273216
rect 344836 273164 344888 273216
rect 354864 273164 354916 273216
rect 177856 273096 177908 273148
rect 227076 273096 227128 273148
rect 264428 273096 264480 273148
rect 267188 273096 267240 273148
rect 292580 273096 292632 273148
rect 331864 273096 331916 273148
rect 355324 273096 355376 273148
rect 362960 273164 363012 273216
rect 491484 273164 491536 273216
rect 148600 273028 148652 273080
rect 223488 273028 223540 273080
rect 243176 273028 243228 273080
rect 259184 273028 259236 273080
rect 260932 273028 260984 273080
rect 265808 273028 265860 273080
rect 293868 273028 293920 273080
rect 335360 273028 335412 273080
rect 358820 273028 358872 273080
rect 497372 273096 497424 273148
rect 149796 272960 149848 273012
rect 224408 272960 224460 273012
rect 241980 272960 242032 273012
rect 258724 272960 258776 273012
rect 293408 272960 293460 273012
rect 334164 272960 334216 273012
rect 344008 272960 344060 273012
rect 362592 272960 362644 273012
rect 498568 273028 498620 273080
rect 498844 273028 498896 273080
rect 617984 273028 618036 273080
rect 504456 272960 504508 273012
rect 42156 272892 42208 272944
rect 43260 272892 43312 272944
rect 150992 272892 151044 272944
rect 223948 272892 224000 272944
rect 239588 272892 239640 272944
rect 257804 272892 257856 272944
rect 304908 272892 304960 272944
rect 346032 272892 346084 272944
rect 357992 272892 358044 272944
rect 505652 272892 505704 272944
rect 143908 272824 143960 272876
rect 221280 272824 221332 272876
rect 236092 272824 236144 272876
rect 256424 272824 256476 272876
rect 307852 272824 307904 272876
rect 348424 272824 348476 272876
rect 360660 272824 360712 272876
rect 512736 272824 512788 272876
rect 145012 272756 145064 272808
rect 222200 272756 222252 272808
rect 234896 272756 234948 272808
rect 256056 272756 256108 272808
rect 300768 272756 300820 272808
rect 353116 272756 353168 272808
rect 360568 272756 360620 272808
rect 511540 272756 511592 272808
rect 511632 272756 511684 272808
rect 610808 272756 610860 272808
rect 146208 272688 146260 272740
rect 223028 272688 223080 272740
rect 232504 272688 232556 272740
rect 255136 272688 255188 272740
rect 294880 272688 294932 272740
rect 338948 272688 339000 272740
rect 344744 272688 344796 272740
rect 470140 272688 470192 272740
rect 471980 272688 472032 272740
rect 625068 272688 625120 272740
rect 139124 272620 139176 272672
rect 220360 272620 220412 272672
rect 237288 272620 237340 272672
rect 257160 272620 257212 272672
rect 301412 272620 301464 272672
rect 355508 272620 355560 272672
rect 363144 272620 363196 272672
rect 518624 272620 518676 272672
rect 137928 272552 137980 272604
rect 219164 272552 219216 272604
rect 233700 272552 233752 272604
rect 255596 272552 255648 272604
rect 300676 272552 300728 272604
rect 351920 272552 351972 272604
rect 353116 272552 353168 272604
rect 362960 272552 363012 272604
rect 368204 272552 368256 272604
rect 532792 272552 532844 272604
rect 136824 272484 136876 272536
rect 218612 272484 218664 272536
rect 230204 272484 230256 272536
rect 254216 272484 254268 272536
rect 296076 272484 296128 272536
rect 341340 272484 341392 272536
rect 342076 272484 342128 272536
rect 463056 272484 463108 272536
rect 465908 272484 465960 272536
rect 632152 272484 632204 272536
rect 132040 272416 132092 272468
rect 217692 272416 217744 272468
rect 301872 272416 301924 272468
rect 356704 272416 356756 272468
rect 373172 272416 373224 272468
rect 545856 272416 545908 272468
rect 124956 272348 125008 272400
rect 215024 272348 215076 272400
rect 303344 272348 303396 272400
rect 360200 272348 360252 272400
rect 376668 272348 376720 272400
rect 555240 272348 555292 272400
rect 129648 272280 129700 272332
rect 215668 272280 215720 272332
rect 294788 272280 294840 272332
rect 337752 272280 337804 272332
rect 339316 272280 339368 272332
rect 455972 272280 456024 272332
rect 459468 272280 459520 272332
rect 639236 272280 639288 272332
rect 117872 272212 117924 272264
rect 206652 272212 206704 272264
rect 302792 272212 302844 272264
rect 359004 272212 359056 272264
rect 382004 272212 382056 272264
rect 569500 272212 569552 272264
rect 93032 272144 93084 272196
rect 184940 272144 184992 272196
rect 188804 272144 188856 272196
rect 234620 272144 234672 272196
rect 238484 272144 238536 272196
rect 257252 272144 257304 272196
rect 306288 272144 306340 272196
rect 367284 272144 367336 272196
rect 384672 272144 384724 272196
rect 576584 272144 576636 272196
rect 104900 272076 104952 272128
rect 202788 272076 202840 272128
rect 205364 272076 205416 272128
rect 240140 272076 240192 272128
rect 308956 272076 309008 272128
rect 374368 272076 374420 272128
rect 387340 272076 387392 272128
rect 583668 272076 583720 272128
rect 89536 272008 89588 272060
rect 178040 272008 178092 272060
rect 178132 272008 178184 272060
rect 197268 272008 197320 272060
rect 199476 272008 199528 272060
rect 242624 272008 242676 272060
rect 284208 272008 284260 272060
rect 309416 272008 309468 272060
rect 311624 272008 311676 272060
rect 381544 272008 381596 272060
rect 394608 272008 394660 272060
rect 590752 272008 590804 272060
rect 75276 271940 75328 271992
rect 195428 271940 195480 271992
rect 201776 271940 201828 271992
rect 243544 271940 243596 271992
rect 285404 271940 285456 271992
rect 312912 271940 312964 271992
rect 314292 271940 314344 271992
rect 388628 271940 388680 271992
rect 395436 271940 395488 271992
rect 604920 271940 604972 271992
rect 66996 271872 67048 271924
rect 192484 271872 192536 271924
rect 65892 271804 65944 271856
rect 192116 271804 192168 271856
rect 120264 271736 120316 271788
rect 156788 271736 156840 271788
rect 156880 271736 156932 271788
rect 177856 271736 177908 271788
rect 177948 271736 178000 271788
rect 194508 271736 194560 271788
rect 130844 271668 130896 271720
rect 197176 271804 197228 271856
rect 198280 271804 198332 271856
rect 242256 271872 242308 271924
rect 244372 271872 244424 271924
rect 259552 271872 259604 271924
rect 290280 271872 290332 271924
rect 325976 271872 326028 271924
rect 326712 271872 326764 271924
rect 402796 271872 402848 271924
rect 402888 271872 402940 271924
rect 619088 271872 619140 271924
rect 194692 271668 194744 271720
rect 240876 271804 240928 271856
rect 245568 271804 245620 271856
rect 260012 271804 260064 271856
rect 289360 271804 289412 271856
rect 323584 271804 323636 271856
rect 325608 271804 325660 271856
rect 409880 271804 409932 271856
rect 411996 271804 412048 271856
rect 633348 271804 633400 271856
rect 240784 271736 240836 271788
rect 258264 271736 258316 271788
rect 262128 271736 262180 271788
rect 266268 271736 266320 271788
rect 292488 271736 292540 271788
rect 330668 271736 330720 271788
rect 349988 271736 350040 271788
rect 484308 271736 484360 271788
rect 208492 271668 208544 271720
rect 226340 271668 226392 271720
rect 229008 271668 229060 271720
rect 253756 271668 253808 271720
rect 290740 271668 290792 271720
rect 327080 271668 327132 271720
rect 336740 271668 336792 271720
rect 343640 271668 343692 271720
rect 350908 271668 350960 271720
rect 486700 271668 486752 271720
rect 165160 271600 165212 271652
rect 229284 271600 229336 271652
rect 231400 271600 231452 271652
rect 254676 271600 254728 271652
rect 289820 271600 289872 271652
rect 324780 271600 324832 271652
rect 348240 271600 348292 271652
rect 479616 271600 479668 271652
rect 163964 271532 164016 271584
rect 229744 271532 229796 271584
rect 249064 271532 249116 271584
rect 261392 271532 261444 271584
rect 291200 271532 291252 271584
rect 328276 271532 328328 271584
rect 347596 271532 347648 271584
rect 477224 271532 477276 271584
rect 158076 271464 158128 271516
rect 177948 271464 178000 271516
rect 178132 271464 178184 271516
rect 228824 271464 228876 271516
rect 252652 271464 252704 271516
rect 262864 271464 262916 271516
rect 288992 271464 289044 271516
rect 322388 271464 322440 271516
rect 342812 271464 342864 271516
rect 465448 271464 465500 271516
rect 171048 271396 171100 271448
rect 232412 271396 232464 271448
rect 258540 271396 258592 271448
rect 264888 271396 264940 271448
rect 288532 271396 288584 271448
rect 321192 271396 321244 271448
rect 354772 271396 354824 271448
rect 472532 271396 472584 271448
rect 172244 271328 172296 271380
rect 162768 271260 162820 271312
rect 178132 271260 178184 271312
rect 180064 271328 180116 271380
rect 231492 271328 231544 271380
rect 256148 271328 256200 271380
rect 264060 271328 264112 271380
rect 286600 271328 286652 271380
rect 315304 271328 315356 271380
rect 340236 271328 340288 271380
rect 458364 271328 458416 271380
rect 231768 271260 231820 271312
rect 255044 271260 255096 271312
rect 263600 271260 263652 271312
rect 287612 271260 287664 271312
rect 318800 271260 318852 271312
rect 337476 271260 337528 271312
rect 451280 271260 451332 271312
rect 178040 271192 178092 271244
rect 189264 271192 189316 271244
rect 197268 271192 197320 271244
rect 232688 271192 232740 271244
rect 251456 271192 251508 271244
rect 262220 271192 262272 271244
rect 266820 271192 266872 271244
rect 268016 271192 268068 271244
rect 287152 271192 287204 271244
rect 317696 271192 317748 271244
rect 329748 271192 329800 271244
rect 340144 271192 340196 271244
rect 179328 271124 179380 271176
rect 234528 271124 234580 271176
rect 247868 271124 247920 271176
rect 260932 271124 260984 271176
rect 286692 271124 286744 271176
rect 316500 271124 316552 271176
rect 336648 271124 336700 271176
rect 448888 271192 448940 271244
rect 169852 271056 169904 271108
rect 180064 271056 180116 271108
rect 182916 271056 182968 271108
rect 232964 271056 233016 271108
rect 253848 271056 253900 271108
rect 263140 271056 263192 271108
rect 288164 271056 288216 271108
rect 319996 271056 320048 271108
rect 334808 271056 334860 271108
rect 415308 271124 415360 271176
rect 420920 271124 420972 271176
rect 441804 271124 441856 271176
rect 176936 270988 176988 271040
rect 227628 270988 227680 271040
rect 246764 270988 246816 271040
rect 260472 270988 260524 271040
rect 285864 270988 285916 271040
rect 314108 270988 314160 271040
rect 333980 270988 334032 271040
rect 420736 271056 420788 271108
rect 185216 270920 185268 270972
rect 234712 270920 234764 270972
rect 250260 270920 250312 270972
rect 261852 270920 261904 270972
rect 331312 270920 331364 270972
rect 186412 270852 186464 270904
rect 233424 270852 233476 270904
rect 329932 270852 329984 270904
rect 175832 270784 175884 270836
rect 179328 270784 179380 270836
rect 190000 270784 190052 270836
rect 231860 270784 231912 270836
rect 259736 270784 259788 270836
rect 265440 270784 265492 270836
rect 327264 270784 327316 270836
rect 340788 270784 340840 270836
rect 187608 270716 187660 270768
rect 230756 270716 230808 270768
rect 326436 270716 326488 270768
rect 395712 270716 395764 270768
rect 191196 270648 191248 270700
rect 192300 270512 192352 270564
rect 198648 270512 198700 270564
rect 229100 270648 229152 270700
rect 257344 270648 257396 270700
rect 264520 270648 264572 270700
rect 331128 270648 331180 270700
rect 377956 270648 378008 270700
rect 227812 270580 227864 270632
rect 253388 270580 253440 270632
rect 324596 270580 324648 270632
rect 340788 270580 340840 270632
rect 351736 270580 351788 270632
rect 394516 270580 394568 270632
rect 415308 270988 415360 271040
rect 444196 271056 444248 271108
rect 434720 270852 434772 270904
rect 431132 270784 431184 270836
rect 424048 270648 424100 270700
rect 416964 270580 417016 270632
rect 226616 270512 226668 270564
rect 252928 270512 252980 270564
rect 357440 270512 357492 270564
rect 385040 270512 385092 270564
rect 411812 270512 411864 270564
rect 413100 270512 413152 270564
rect 152188 270444 152240 270496
rect 208032 270444 208084 270496
rect 147404 270376 147456 270428
rect 208124 270376 208176 270428
rect 141516 270308 141568 270360
rect 220820 270444 220872 270496
rect 225420 270444 225472 270496
rect 252468 270444 252520 270496
rect 265624 270444 265676 270496
rect 267556 270444 267608 270496
rect 269856 270444 269908 270496
rect 271512 270444 271564 270496
rect 272064 270444 272116 270496
rect 277492 270444 277544 270496
rect 304080 270444 304132 270496
rect 344008 270444 344060 270496
rect 346860 270444 346912 270496
rect 476120 270444 476172 270496
rect 140320 270240 140372 270292
rect 219992 270376 220044 270428
rect 221924 270376 221976 270428
rect 251088 270376 251140 270428
rect 270316 270376 270368 270428
rect 272708 270376 272760 270428
rect 273720 270376 273772 270428
rect 280988 270376 281040 270428
rect 294328 270376 294380 270428
rect 336556 270376 336608 270428
rect 348608 270376 348660 270428
rect 480812 270376 480864 270428
rect 219072 270308 219124 270360
rect 224224 270308 224276 270360
rect 252008 270308 252060 270360
rect 271144 270308 271196 270360
rect 275100 270308 275152 270360
rect 277400 270308 277452 270360
rect 291660 270308 291712 270360
rect 296996 270308 297048 270360
rect 336740 270308 336792 270360
rect 349528 270308 349580 270360
rect 483204 270308 483256 270360
rect 133236 270172 133288 270224
rect 202512 270172 202564 270224
rect 202604 270172 202656 270224
rect 214656 270172 214708 270224
rect 135628 270104 135680 270156
rect 219532 270240 219584 270292
rect 250260 270240 250312 270292
rect 274272 270240 274324 270292
rect 283380 270240 283432 270292
rect 283472 270240 283524 270292
rect 290464 270240 290516 270292
rect 297456 270240 297508 270292
rect 339500 270240 339552 270292
rect 351276 270240 351328 270292
rect 487896 270240 487948 270292
rect 217140 270172 217192 270224
rect 249340 270172 249392 270224
rect 277860 270172 277912 270224
rect 292856 270172 292908 270224
rect 296536 270172 296588 270224
rect 342444 270172 342496 270224
rect 352196 270172 352248 270224
rect 490288 270172 490340 270224
rect 134432 270036 134484 270088
rect 218152 270104 218204 270156
rect 223120 270104 223172 270156
rect 251548 270104 251600 270156
rect 278596 270104 278648 270156
rect 295156 270104 295208 270156
rect 298284 270104 298336 270156
rect 347228 270104 347280 270156
rect 353576 270104 353628 270156
rect 493784 270104 493836 270156
rect 220728 270036 220780 270088
rect 250720 270036 250772 270088
rect 278320 270036 278372 270088
rect 294052 270036 294104 270088
rect 299204 270036 299256 270088
rect 349620 270036 349672 270088
rect 356244 270036 356296 270088
rect 500868 270036 500920 270088
rect 126152 269968 126204 270020
rect 202604 269968 202656 270020
rect 119068 269900 119120 269952
rect 211896 269968 211948 270020
rect 215944 269968 215996 270020
rect 248880 269968 248932 270020
rect 279148 269968 279200 270020
rect 296352 269968 296404 270020
rect 345480 269968 345532 270020
rect 354772 269968 354824 270020
rect 364708 269968 364760 270020
rect 114284 269832 114336 269884
rect 211068 269900 211120 269952
rect 214840 269900 214892 269952
rect 248420 269900 248472 269952
rect 279608 269900 279660 269952
rect 297548 269900 297600 269952
rect 305460 269900 305512 269952
rect 366088 269900 366140 269952
rect 367376 269900 367428 269952
rect 382464 269968 382516 270020
rect 515128 269968 515180 270020
rect 110788 269764 110840 269816
rect 209688 269832 209740 269884
rect 210056 269832 210108 269884
rect 246672 269832 246724 269884
rect 274732 269832 274784 269884
rect 284576 269832 284628 269884
rect 306748 269832 306800 269884
rect 369676 269832 369728 269884
rect 370044 269832 370096 269884
rect 523408 269900 523460 269952
rect 202972 269764 203024 269816
rect 208400 269764 208452 269816
rect 212448 269764 212500 269816
rect 247592 269764 247644 269816
rect 280528 269764 280580 269816
rect 299940 269764 299992 269816
rect 307208 269764 307260 269816
rect 370872 269764 370924 269816
rect 109592 269696 109644 269748
rect 95424 269628 95476 269680
rect 203524 269628 203576 269680
rect 102508 269560 102560 269612
rect 206192 269560 206244 269612
rect 207756 269696 207808 269748
rect 245752 269696 245804 269748
rect 280068 269696 280120 269748
rect 298744 269696 298796 269748
rect 308128 269696 308180 269748
rect 373264 269764 373316 269816
rect 530492 269832 530544 269884
rect 537576 269764 537628 269816
rect 375380 269696 375432 269748
rect 206560 269628 206612 269680
rect 224132 269628 224184 269680
rect 234620 269628 234672 269680
rect 239128 269628 239180 269680
rect 281816 269628 281868 269680
rect 303436 269628 303488 269680
rect 328644 269628 328696 269680
rect 351920 269628 351972 269680
rect 361580 269628 361632 269680
rect 382280 269628 382332 269680
rect 382464 269696 382516 269748
rect 544660 269696 544712 269748
rect 703544 269696 703596 269748
rect 704004 269696 704056 269748
rect 708880 269696 708932 269748
rect 708972 269696 709024 269748
rect 551744 269628 551796 269680
rect 208860 269560 208912 269612
rect 209136 269560 209188 269612
rect 246212 269560 246264 269612
rect 281448 269560 281500 269612
rect 302332 269560 302384 269612
rect 310796 269560 310848 269612
rect 380348 269560 380400 269612
rect 380716 269560 380768 269612
rect 565912 269560 565964 269612
rect 708052 269628 708104 269680
rect 704924 269560 704976 269612
rect 707960 269560 708012 269612
rect 94228 269492 94280 269544
rect 202604 269492 202656 269544
rect 204168 269492 204220 269544
rect 244464 269492 244516 269544
rect 280988 269492 281040 269544
rect 301136 269492 301188 269544
rect 312084 269492 312136 269544
rect 383844 269492 383896 269544
rect 386052 269492 386104 269544
rect 580080 269492 580132 269544
rect 704832 269492 704884 269544
rect 74080 269424 74132 269476
rect 195888 269424 195940 269476
rect 198648 269424 198700 269476
rect 80060 269356 80112 269408
rect 197268 269356 197320 269408
rect 197360 269356 197412 269408
rect 208400 269424 208452 269476
rect 244004 269424 244056 269476
rect 282736 269424 282788 269476
rect 305828 269424 305880 269476
rect 313464 269424 313516 269476
rect 387432 269424 387484 269476
rect 388720 269424 388772 269476
rect 587164 269424 587216 269476
rect 707040 269492 707092 269544
rect 706672 269424 706724 269476
rect 82360 269288 82412 269340
rect 198556 269288 198608 269340
rect 239956 269356 240008 269408
rect 282276 269356 282328 269408
rect 304632 269356 304684 269408
rect 314844 269356 314896 269408
rect 390928 269356 390980 269408
rect 394056 269356 394108 269408
rect 601424 269356 601476 269408
rect 705752 269356 705804 269408
rect 706212 269356 706264 269408
rect 706304 269356 706356 269408
rect 706580 269356 706632 269408
rect 241796 269288 241848 269340
rect 276940 269288 276992 269340
rect 283472 269288 283524 269340
rect 283656 269288 283708 269340
rect 308220 269288 308272 269340
rect 315212 269288 315264 269340
rect 392124 269288 392176 269340
rect 396724 269288 396776 269340
rect 608508 269288 608560 269340
rect 705844 269288 705896 269340
rect 707040 269288 707092 269340
rect 707592 269288 707644 269340
rect 81256 269220 81308 269272
rect 198096 269220 198148 269272
rect 200580 269220 200632 269272
rect 243084 269220 243136 269272
rect 283196 269220 283248 269272
rect 307024 269220 307076 269272
rect 317880 269220 317932 269272
rect 399208 269220 399260 269272
rect 399392 269220 399444 269272
rect 615592 269220 615644 269272
rect 705384 269220 705436 269272
rect 707500 269220 707552 269272
rect 71780 269152 71832 269204
rect 194600 269152 194652 269204
rect 195796 269152 195848 269204
rect 241336 269152 241388 269204
rect 284944 269152 284996 269204
rect 311716 269152 311768 269204
rect 320548 269152 320600 269204
rect 406292 269152 406344 269204
rect 411444 269152 411496 269204
rect 647516 269152 647568 269204
rect 705292 269152 705344 269204
rect 708512 269152 708564 269204
rect 193496 269084 193548 269136
rect 240416 269084 240468 269136
rect 269396 269084 269448 269136
rect 270408 269084 270460 269136
rect 284484 269084 284536 269136
rect 310520 269084 310572 269136
rect 323216 269084 323268 269136
rect 411812 269084 411864 269136
rect 411904 269084 411956 269136
rect 648712 269084 648764 269136
rect 704464 269084 704516 269136
rect 708420 269084 708472 269136
rect 154488 269016 154540 269068
rect 225328 269016 225380 269068
rect 292948 269016 293000 269068
rect 333060 269016 333112 269068
rect 159272 268948 159324 269000
rect 224040 268948 224092 269000
rect 224132 268948 224184 269000
rect 245292 268948 245344 269000
rect 295616 268948 295668 269000
rect 329748 268948 329800 269000
rect 330852 268948 330904 269000
rect 351828 269016 351880 269068
rect 345940 268948 345992 269000
rect 473728 269016 473780 269068
rect 704372 269016 704424 269068
rect 352012 268948 352064 269000
rect 466644 268948 466696 269000
rect 160468 268880 160520 268932
rect 161572 268812 161624 268864
rect 223764 268812 223816 268864
rect 231860 268880 231912 268932
rect 238668 268880 238720 268932
rect 309876 268880 309928 268932
rect 331128 268880 331180 268932
rect 344192 268880 344244 268932
rect 468944 268880 468996 268932
rect 228456 268812 228508 268864
rect 229100 268812 229152 268864
rect 239588 268812 239640 268864
rect 272984 268812 273036 268864
rect 279792 268812 279844 268864
rect 341524 268812 341576 268864
rect 461860 268812 461912 268864
rect 166356 268744 166408 268796
rect 167552 268676 167604 268728
rect 224040 268744 224092 268796
rect 227536 268744 227588 268796
rect 340604 268744 340656 268796
rect 459560 268744 459612 268796
rect 173440 268608 173492 268660
rect 223580 268608 223632 268660
rect 230204 268676 230256 268728
rect 273812 268676 273864 268728
rect 282184 268676 282236 268728
rect 338856 268676 338908 268728
rect 454776 268676 454828 268728
rect 231124 268608 231176 268660
rect 337936 268608 337988 268660
rect 452476 268608 452528 268660
rect 168656 268540 168708 268592
rect 230664 268540 230716 268592
rect 230756 268540 230808 268592
rect 236644 268540 236696 268592
rect 240140 268540 240192 268592
rect 244924 268540 244976 268592
rect 336188 268540 336240 268592
rect 447692 268540 447744 268592
rect 156788 268472 156840 268524
rect 212816 268472 212868 268524
rect 213644 268472 213696 268524
rect 248052 268472 248104 268524
rect 335268 268472 335320 268524
rect 445300 268472 445352 268524
rect 174636 268404 174688 268456
rect 233792 268404 233844 268456
rect 272524 268404 272576 268456
rect 278688 268404 278740 268456
rect 325976 268404 326028 268456
rect 332784 268404 332836 268456
rect 333520 268404 333572 268456
rect 440608 268404 440660 268456
rect 179328 268336 179380 268388
rect 233332 268336 233384 268388
rect 233424 268336 233476 268388
rect 237288 268336 237340 268388
rect 309416 268336 309468 268388
rect 332508 268336 332560 268388
rect 332600 268336 332652 268388
rect 438216 268336 438268 268388
rect 181720 268268 181772 268320
rect 223580 268268 223632 268320
rect 223672 268268 223724 268320
rect 232872 268268 232924 268320
rect 232964 268268 233016 268320
rect 236000 268268 236052 268320
rect 275192 268268 275244 268320
rect 285772 268268 285824 268320
rect 312544 268268 312596 268320
rect 180524 268200 180576 268252
rect 235540 268200 235592 268252
rect 270684 268200 270736 268252
rect 273904 268200 273956 268252
rect 275652 268200 275704 268252
rect 286876 268200 286928 268252
rect 316132 268200 316184 268252
rect 184112 268132 184164 268184
rect 236920 268132 236972 268184
rect 316592 268132 316644 268184
rect 326436 268132 326488 268184
rect 197176 268064 197228 268116
rect 216864 268064 216916 268116
rect 218336 268064 218388 268116
rect 189264 267996 189316 268048
rect 200764 267996 200816 268048
rect 201316 267996 201368 268048
rect 203892 267996 203944 268048
rect 208124 267996 208176 268048
rect 222660 267996 222712 268048
rect 223580 268064 223632 268116
rect 236460 268064 236512 268116
rect 249800 268064 249852 268116
rect 236644 267996 236696 268048
rect 238208 267996 238260 268048
rect 271604 267996 271656 268048
rect 276296 267996 276348 268048
rect 276388 267996 276440 268048
rect 288072 267996 288124 268048
rect 298744 267996 298796 268048
rect 307852 267996 307904 268048
rect 319260 267996 319312 268048
rect 326712 267996 326764 268048
rect 88340 267928 88392 267980
rect 201224 267928 201276 267980
rect 211252 267928 211304 267980
rect 208032 267860 208084 267912
rect 224868 267860 224920 267912
rect 202512 267792 202564 267844
rect 217324 267792 217376 267844
rect 223764 267792 223816 267844
rect 227996 267792 228048 267844
rect 232688 267792 232740 267844
rect 235080 267792 235132 267844
rect 247132 267928 247184 267980
rect 297916 267928 297968 267980
rect 304908 267928 304960 267980
rect 321928 267928 321980 267980
rect 325608 267928 325660 267980
rect 351828 268268 351880 268320
rect 433524 268268 433576 268320
rect 332692 268200 332744 268252
rect 426440 268200 426492 268252
rect 351920 268132 351972 268184
rect 427636 268132 427688 268184
rect 332784 268064 332836 268116
rect 420552 268064 420604 268116
rect 666468 268064 666520 268116
rect 676220 268064 676272 268116
rect 357440 267996 357492 268048
rect 357532 267996 357584 268048
rect 358728 267996 358780 268048
rect 372712 267996 372764 268048
rect 382464 267996 382516 268048
rect 390008 267996 390060 268048
rect 394608 267996 394660 268048
rect 400772 267996 400824 268048
rect 402888 267996 402940 268048
rect 406108 267996 406160 268048
rect 411996 267996 412048 268048
rect 351736 267928 351788 267980
rect 661132 267928 661184 267980
rect 676036 267928 676088 267980
rect 276480 267860 276532 267912
rect 289268 267860 289320 267912
rect 328000 267860 328052 267912
rect 332692 267860 332744 267912
rect 343272 267860 343324 267912
rect 352012 267860 352064 267912
rect 304540 267792 304592 267844
rect 363788 267792 363840 267844
rect 202788 267724 202840 267776
rect 206560 267724 206612 267776
rect 206652 267724 206704 267776
rect 212356 267724 212408 267776
rect 227628 267724 227680 267776
rect 234160 267724 234212 267776
rect 234712 267724 234764 267776
rect 237748 267724 237800 267776
rect 332508 267724 332560 267776
rect 376760 267724 376812 267776
rect 660948 267724 661000 267776
rect 676128 267724 676180 267776
rect 359740 267656 359792 267708
rect 510344 267656 510396 267708
rect 674748 267656 674800 267708
rect 676036 267656 676088 267708
rect 362408 267588 362460 267640
rect 517428 267588 517480 267640
rect 365076 267520 365128 267572
rect 524512 267520 524564 267572
rect 367744 267452 367796 267504
rect 531596 267452 531648 267504
rect 672264 267452 672316 267504
rect 675944 267452 675996 267504
rect 370504 267384 370556 267436
rect 538772 267384 538824 267436
rect 373540 267316 373592 267368
rect 547052 267316 547104 267368
rect 374460 267248 374512 267300
rect 549352 267248 549404 267300
rect 376208 267180 376260 267232
rect 554136 267180 554188 267232
rect 299664 267112 299716 267164
rect 350724 267112 350776 267164
rect 375840 267112 375892 267164
rect 552940 267112 552992 267164
rect 300952 267044 301004 267096
rect 354312 267044 354364 267096
rect 377128 267044 377180 267096
rect 556436 267044 556488 267096
rect 302332 266976 302384 267028
rect 357900 266976 357952 267028
rect 378508 266976 378560 267028
rect 560024 266976 560076 267028
rect 303712 266908 303764 266960
rect 361396 266908 361448 266960
rect 378876 266908 378928 266960
rect 561220 266908 561272 266960
rect 305000 266840 305052 266892
rect 364984 266840 365036 266892
rect 379796 266840 379848 266892
rect 563520 266840 563572 266892
rect 306380 266772 306432 266824
rect 368480 266772 368532 266824
rect 381636 266772 381688 266824
rect 568304 266772 568356 266824
rect 307668 266704 307720 266756
rect 372068 266704 372120 266756
rect 381176 266704 381228 266756
rect 567108 266704 567160 266756
rect 309048 266636 309100 266688
rect 375564 266636 375616 266688
rect 382464 266636 382516 266688
rect 570696 266636 570748 266688
rect 123760 266568 123812 266620
rect 214196 266568 214248 266620
rect 310336 266568 310388 266620
rect 379152 266568 379204 266620
rect 384304 266568 384356 266620
rect 575388 266568 575440 266620
rect 116676 266500 116728 266552
rect 211528 266500 211580 266552
rect 311716 266500 311768 266552
rect 382648 266500 382700 266552
rect 383844 266500 383896 266552
rect 574192 266500 574244 266552
rect 72976 266432 73028 266484
rect 195060 266432 195112 266484
rect 313004 266432 313056 266484
rect 386236 266432 386288 266484
rect 389180 266432 389232 266484
rect 588360 266432 588412 266484
rect 113180 266364 113232 266416
rect 210148 266364 210200 266416
rect 315672 266364 315724 266416
rect 68192 266296 68244 266348
rect 193220 266296 193272 266348
rect 317052 266296 317104 266348
rect 382188 266296 382240 266348
rect 392308 266364 392360 266416
rect 596640 266364 596692 266416
rect 393320 266296 393372 266348
rect 394976 266296 395028 266348
rect 603724 266296 603776 266348
rect 652944 266296 652996 266348
rect 675668 266296 675720 266348
rect 357072 266228 357124 266280
rect 503260 266228 503312 266280
rect 353208 266160 353260 266212
rect 492588 266160 492640 266212
rect 351736 266092 351788 266144
rect 489092 266092 489144 266144
rect 671896 266092 671948 266144
rect 676220 266092 676272 266144
rect 347780 266024 347832 266076
rect 478420 266024 478472 266076
rect 346400 265956 346452 266008
rect 474924 265956 474976 266008
rect 339776 265888 339828 265940
rect 457168 265888 457220 265940
rect 338396 265820 338448 265872
rect 453580 265820 453632 265872
rect 317512 265752 317564 265804
rect 382096 265752 382148 265804
rect 382188 265752 382240 265804
rect 396908 265752 396960 265804
rect 397644 265752 397696 265804
rect 511632 265752 511684 265804
rect 329472 265684 329524 265736
rect 429936 265684 429988 265736
rect 382280 265616 382332 265668
rect 398012 265616 398064 265668
rect 400312 265616 400364 265668
rect 498844 265616 498896 265668
rect 325516 265548 325568 265600
rect 419356 265548 419408 265600
rect 324136 265480 324188 265532
rect 415768 265480 415820 265532
rect 322848 265412 322900 265464
rect 412272 265412 412324 265464
rect 321468 265344 321520 265396
rect 408684 265344 408736 265396
rect 674748 265344 674800 265396
rect 676036 265344 676088 265396
rect 318340 265276 318392 265328
rect 400404 265276 400456 265328
rect 402980 265276 403032 265328
rect 471980 265276 472032 265328
rect 314384 265208 314436 265260
rect 389732 265208 389784 265260
rect 319720 265140 319772 265192
rect 403992 265140 404044 265192
rect 658280 264936 658332 264988
rect 675760 265004 675812 265056
rect 673184 264936 673236 264988
rect 676220 264936 676272 264988
rect 674196 263032 674248 263084
rect 676036 263032 676088 263084
rect 673736 262352 673788 262404
rect 675944 262352 675996 262404
rect 674012 262284 674064 262336
rect 676128 262284 676180 262336
rect 418068 262216 418120 262268
rect 571708 262216 571760 262268
rect 674288 262216 674340 262268
rect 676036 262216 676088 262268
rect 674104 261808 674156 261860
rect 676036 261808 676088 261860
rect 673460 260176 673512 260228
rect 675576 260176 675628 260228
rect 673552 259700 673604 259752
rect 675576 259700 675628 259752
rect 674472 259632 674524 259684
rect 676128 259632 676180 259684
rect 674380 259564 674432 259616
rect 675944 259564 675996 259616
rect 675024 259496 675076 259548
rect 676128 259496 676180 259548
rect 52276 259428 52328 259480
rect 184940 259428 184992 259480
rect 417792 259428 417844 259480
rect 571800 259428 571852 259480
rect 675208 259428 675260 259480
rect 676036 259428 676088 259480
rect 41512 258340 41564 258392
rect 48412 258340 48464 258392
rect 41788 257796 41840 257848
rect 53932 257796 53984 257848
rect 41512 257524 41564 257576
rect 50988 257524 51040 257576
rect 41788 256844 41840 256896
rect 45836 256844 45888 256896
rect 672816 256844 672868 256896
rect 678980 256844 679032 256896
rect 673644 256776 673696 256828
rect 676128 256776 676180 256828
rect 418344 256708 418396 256760
rect 571524 256708 571576 256760
rect 673828 256708 673880 256760
rect 676036 256708 676088 256760
rect 674748 255280 674800 255332
rect 675668 255280 675720 255332
rect 674656 255212 674708 255264
rect 675760 255212 675812 255264
rect 416780 253920 416832 253972
rect 574100 253920 574152 253972
rect 52184 251200 52236 251252
rect 184940 251200 184992 251252
rect 416780 251200 416832 251252
rect 572628 251200 572680 251252
rect 675760 251200 675812 251252
rect 675760 250928 675812 250980
rect 675208 250384 675260 250436
rect 675484 250384 675536 250436
rect 33048 249772 33100 249824
rect 43628 249772 43680 249824
rect 674196 249568 674248 249620
rect 675392 249568 675444 249620
rect 416780 248412 416832 248464
rect 569868 248412 569920 248464
rect 674288 247868 674340 247920
rect 675484 247868 675536 247920
rect 41512 247664 41564 247716
rect 45928 247664 45980 247716
rect 41512 247256 41564 247308
rect 45836 247256 45888 247308
rect 674472 247256 674524 247308
rect 675392 247256 675444 247308
rect 674012 247120 674064 247172
rect 674472 247120 674524 247172
rect 41512 246848 41564 246900
rect 45744 246848 45796 246900
rect 674380 246508 674432 246560
rect 675392 246508 675444 246560
rect 675116 246032 675168 246084
rect 675392 246032 675444 246084
rect 43628 244740 43680 244792
rect 43904 244740 43956 244792
rect 43352 244604 43404 244656
rect 43628 244604 43680 244656
rect 42892 244536 42944 244588
rect 43536 244536 43588 244588
rect 42708 244468 42760 244520
rect 43352 244468 43404 244520
rect 33048 244400 33100 244452
rect 42892 244400 42944 244452
rect 32864 244332 32916 244384
rect 43168 244332 43220 244384
rect 32956 244264 33008 244316
rect 42984 244264 43036 244316
rect 31668 244196 31720 244248
rect 42708 244196 42760 244248
rect 673736 243584 673788 243636
rect 675300 243584 675352 243636
rect 52092 242904 52144 242956
rect 184940 242904 184992 242956
rect 673828 242904 673880 242956
rect 675300 242904 675352 242956
rect 38292 242836 38344 242888
rect 42800 242836 42852 242888
rect 673552 242156 673604 242208
rect 675392 242156 675444 242208
rect 674472 241884 674524 241936
rect 675300 241884 675352 241936
rect 673644 241544 673696 241596
rect 675392 241544 675444 241596
rect 673460 240524 673512 240576
rect 675392 240524 675444 240576
rect 42156 240320 42208 240372
rect 43720 240320 43772 240372
rect 224132 238552 224184 238604
rect 42156 238416 42208 238468
rect 42708 238416 42760 238468
rect 224132 238348 224184 238400
rect 161388 237328 161440 237380
rect 237196 237328 237248 237380
rect 238944 237328 238996 237380
rect 266728 237328 266780 237380
rect 329196 237328 329248 237380
rect 375748 237328 375800 237380
rect 395436 237328 395488 237380
rect 533988 237328 534040 237380
rect 165436 237260 165488 237312
rect 240416 237260 240468 237312
rect 241612 237260 241664 237312
rect 269580 237260 269632 237312
rect 314936 237260 314988 237312
rect 342720 237260 342772 237312
rect 397276 237260 397328 237312
rect 535460 237260 535512 237312
rect 142160 237192 142212 237244
rect 218980 237192 219032 237244
rect 254860 237192 254912 237244
rect 263876 237192 263928 237244
rect 312084 237192 312136 237244
rect 334440 237192 334492 237244
rect 399392 237192 399444 237244
rect 539508 237192 539560 237244
rect 159824 237124 159876 237176
rect 237564 237124 237616 237176
rect 238852 237124 238904 237176
rect 265348 237124 265400 237176
rect 302424 237124 302476 237176
rect 312820 237124 312872 237176
rect 317420 237124 317472 237176
rect 329748 237124 329800 237176
rect 400496 237124 400548 237176
rect 542268 237124 542320 237176
rect 153200 237056 153252 237108
rect 234344 237056 234396 237108
rect 242808 237056 242860 237108
rect 272156 237056 272208 237108
rect 401140 237056 401192 237108
rect 545120 237056 545172 237108
rect 147588 236988 147640 237040
rect 229008 236988 229060 237040
rect 245476 236988 245528 237040
rect 273536 236988 273588 237040
rect 302792 236988 302844 237040
rect 309784 236988 309836 237040
rect 405096 236988 405148 237040
rect 413468 236988 413520 237040
rect 413560 236988 413612 237040
rect 545028 236988 545080 237040
rect 136548 236920 136600 236972
rect 216128 236920 216180 236972
rect 223488 236920 223540 236972
rect 254860 236920 254912 236972
rect 258080 236920 258132 236972
rect 128268 236852 128320 236904
rect 197268 236852 197320 236904
rect 206376 236852 206428 236904
rect 226156 236852 226208 236904
rect 226248 236852 226300 236904
rect 258172 236852 258224 236904
rect 264704 236920 264756 236972
rect 280988 236920 281040 236972
rect 301688 236920 301740 236972
rect 309968 236920 310020 236972
rect 325976 236920 326028 236972
rect 343364 236920 343416 236972
rect 399024 236920 399076 236972
rect 542360 236920 542412 236972
rect 277492 236852 277544 236904
rect 318800 236852 318852 236904
rect 338120 236852 338172 236904
rect 402980 236852 403032 236904
rect 550364 236852 550416 236904
rect 674380 236852 674432 236904
rect 675392 236852 675444 236904
rect 155868 236784 155920 236836
rect 234712 236784 234764 236836
rect 241428 236784 241480 236836
rect 271052 236784 271104 236836
rect 320272 236784 320324 236836
rect 340880 236784 340932 236836
rect 403348 236784 403400 236836
rect 550548 236784 550600 236836
rect 139308 236716 139360 236768
rect 218612 236716 218664 236768
rect 220728 236716 220780 236768
rect 264244 236716 264296 236768
rect 264888 236716 264940 236768
rect 281724 236716 281776 236768
rect 324504 236716 324556 236768
rect 343272 236716 343324 236768
rect 405464 236716 405516 236768
rect 413652 236716 413704 236768
rect 413744 236716 413796 236768
rect 547788 236716 547840 236768
rect 42156 236648 42208 236700
rect 42892 236648 42944 236700
rect 117228 236648 117280 236700
rect 199752 236648 199804 236700
rect 200856 236648 200908 236700
rect 252468 236648 252520 236700
rect 253204 236648 253256 236700
rect 263232 236648 263284 236700
rect 150348 236580 150400 236632
rect 231860 236580 231912 236632
rect 237288 236580 237340 236632
rect 269304 236648 269356 236700
rect 303160 236648 303212 236700
rect 312636 236648 312688 236700
rect 404728 236648 404780 236700
rect 552296 236648 552348 236700
rect 270408 236580 270460 236632
rect 284576 236580 284628 236632
rect 406844 236580 406896 236632
rect 557540 236580 557592 236632
rect 142068 236512 142120 236564
rect 206376 236512 206428 236564
rect 119988 236444 120040 236496
rect 202604 236444 202656 236496
rect 203248 236444 203300 236496
rect 209688 236444 209740 236496
rect 226156 236444 226208 236496
rect 239956 236512 240008 236564
rect 270684 236512 270736 236564
rect 407212 236512 407264 236564
rect 413376 236512 413428 236564
rect 413468 236512 413520 236564
rect 556160 236512 556212 236564
rect 255320 236444 255372 236496
rect 259276 236444 259328 236496
rect 279976 236444 280028 236496
rect 317788 236444 317840 236496
rect 348148 236444 348200 236496
rect 407580 236444 407632 236496
rect 413560 236444 413612 236496
rect 413652 236444 413704 236496
rect 556068 236444 556120 236496
rect 125508 236376 125560 236428
rect 215760 236376 215812 236428
rect 220636 236376 220688 236428
rect 253204 236376 253256 236428
rect 122748 236308 122800 236360
rect 213276 236308 213328 236360
rect 216680 236308 216732 236360
rect 261024 236376 261076 236428
rect 264796 236376 264848 236428
rect 282828 236376 282880 236428
rect 302056 236376 302108 236428
rect 312268 236376 312320 236428
rect 316316 236376 316368 236428
rect 345388 236376 345440 236428
rect 401508 236376 401560 236428
rect 406384 236376 406436 236428
rect 409052 236376 409104 236428
rect 563152 236376 563204 236428
rect 260840 236308 260892 236360
rect 278872 236308 278924 236360
rect 303528 236308 303580 236360
rect 315028 236308 315080 236360
rect 319168 236308 319220 236360
rect 351092 236308 351144 236360
rect 396172 236308 396224 236360
rect 399300 236308 399352 236360
rect 409328 236308 409380 236360
rect 565544 236308 565596 236360
rect 103428 236240 103480 236292
rect 196900 236240 196952 236292
rect 205732 236240 205784 236292
rect 254308 236240 254360 236292
rect 256516 236240 256568 236292
rect 278504 236240 278556 236292
rect 320640 236240 320692 236292
rect 356428 236240 356480 236292
rect 387616 236240 387668 236292
rect 401508 236240 401560 236292
rect 413376 236240 413428 236292
rect 561588 236240 561640 236292
rect 111708 236172 111760 236224
rect 197176 236172 197228 236224
rect 197268 236172 197320 236224
rect 207204 236172 207256 236224
rect 210976 236172 211028 236224
rect 260012 236172 260064 236224
rect 260748 236172 260800 236224
rect 280344 236172 280396 236224
rect 303804 236172 303856 236224
rect 317972 236172 318024 236224
rect 322020 236172 322072 236224
rect 359188 236172 359240 236224
rect 379428 236172 379480 236224
rect 390376 236172 390428 236224
rect 400772 236172 400824 236224
rect 413284 236172 413336 236224
rect 413560 236172 413612 236224
rect 561680 236172 561732 236224
rect 86868 236104 86920 236156
rect 203340 236104 203392 236156
rect 204168 236104 204220 236156
rect 257160 236104 257212 236156
rect 259368 236104 259420 236156
rect 279240 236104 279292 236156
rect 309232 236104 309284 236156
rect 328644 236104 328696 236156
rect 377956 236104 378008 236156
rect 387616 236104 387668 236156
rect 390836 236104 390888 236156
rect 401600 236104 401652 236156
rect 410064 236104 410116 236156
rect 565820 236104 565872 236156
rect 67548 236036 67600 236088
rect 192944 236036 192996 236088
rect 193036 236036 193088 236088
rect 251824 236036 251876 236088
rect 253756 236036 253808 236088
rect 276388 236036 276440 236088
rect 300952 236036 301004 236088
rect 309416 236036 309468 236088
rect 330576 236036 330628 236088
rect 378508 236036 378560 236088
rect 410432 236036 410484 236088
rect 568028 236036 568080 236088
rect 73160 235968 73212 236020
rect 200120 235968 200172 236020
rect 201408 235968 201460 236020
rect 254676 235968 254728 236020
rect 255412 235968 255464 236020
rect 277124 235968 277176 236020
rect 298100 235968 298152 236020
rect 303804 235968 303856 236020
rect 313464 235968 313516 236020
rect 337108 235968 337160 236020
rect 338396 235968 338448 236020
rect 395160 235968 395212 236020
rect 410800 235968 410852 236020
rect 569960 235968 570012 236020
rect 168104 235900 168156 235952
rect 241152 235900 241204 235952
rect 245568 235900 245620 235952
rect 248328 235900 248380 235952
rect 273904 235900 273956 235952
rect 310612 235900 310664 235952
rect 331772 235900 331824 235952
rect 334532 235900 334584 235952
rect 346492 235900 346544 235952
rect 397644 235900 397696 235952
rect 536748 235900 536800 235952
rect 165344 235832 165396 235884
rect 239772 235832 239824 235884
rect 272432 235832 272484 235884
rect 299940 235832 299992 235884
rect 304080 235832 304132 235884
rect 393320 235832 393372 235884
rect 528468 235832 528520 235884
rect 173716 235764 173768 235816
rect 244280 235764 244332 235816
rect 250996 235764 251048 235816
rect 275284 235764 275336 235816
rect 395068 235764 395120 235816
rect 529940 235764 529992 235816
rect 173808 235696 173860 235748
rect 243268 235696 243320 235748
rect 247316 235696 247368 235748
rect 261392 235696 261444 235748
rect 267188 235696 267240 235748
rect 281356 235696 281408 235748
rect 299204 235696 299256 235748
rect 303712 235696 303764 235748
rect 197268 235628 197320 235680
rect 246120 235628 246172 235680
rect 251088 235628 251140 235680
rect 275008 235628 275060 235680
rect 301320 235628 301372 235680
rect 307300 235696 307352 235748
rect 392952 235696 393004 235748
rect 524420 235696 524472 235748
rect 306656 235628 306708 235680
rect 308772 235628 308824 235680
rect 401600 235628 401652 235680
rect 520188 235628 520240 235680
rect 158628 235560 158680 235612
rect 208124 235560 208176 235612
rect 155960 235492 156012 235544
rect 222936 235560 222988 235612
rect 224040 235560 224092 235612
rect 224684 235560 224736 235612
rect 161572 235424 161624 235476
rect 208216 235424 208268 235476
rect 223304 235492 223356 235544
rect 42156 235356 42208 235408
rect 42800 235356 42852 235408
rect 156052 235356 156104 235408
rect 208400 235356 208452 235408
rect 231492 235356 231544 235408
rect 183468 235288 183520 235340
rect 247132 235560 247184 235612
rect 244280 235492 244332 235544
rect 249984 235492 250036 235544
rect 236092 235424 236144 235476
rect 259644 235560 259696 235612
rect 261944 235560 261996 235612
rect 279608 235560 279660 235612
rect 299572 235560 299624 235612
rect 307208 235560 307260 235612
rect 331680 235560 331732 235612
rect 346400 235560 346452 235612
rect 386236 235560 386288 235612
rect 393780 235560 393832 235612
rect 393964 235560 394016 235612
rect 512000 235560 512052 235612
rect 674748 235560 674800 235612
rect 675668 235560 675720 235612
rect 258172 235492 258224 235544
rect 276020 235492 276072 235544
rect 300308 235492 300360 235544
rect 306656 235492 306708 235544
rect 394056 235492 394108 235544
rect 401416 235492 401468 235544
rect 401508 235492 401560 235544
rect 513472 235492 513524 235544
rect 674656 235492 674708 235544
rect 675760 235492 675812 235544
rect 256608 235424 256660 235476
rect 277860 235424 277912 235476
rect 388720 235424 388772 235476
rect 511908 235424 511960 235476
rect 233424 235356 233476 235408
rect 244188 235356 244240 235408
rect 245752 235356 245804 235408
rect 255320 235356 255372 235408
rect 274272 235356 274324 235408
rect 333060 235356 333112 235408
rect 346216 235356 346268 235408
rect 385500 235356 385552 235408
rect 507952 235356 508004 235408
rect 190368 235220 190420 235272
rect 251456 235220 251508 235272
rect 255228 235288 255280 235340
rect 275652 235288 275704 235340
rect 306380 235288 306432 235340
rect 321008 235288 321060 235340
rect 384028 235288 384080 235340
rect 506388 235288 506440 235340
rect 256792 235220 256844 235272
rect 262036 235220 262088 235272
rect 267188 235220 267240 235272
rect 267280 235220 267332 235272
rect 280712 235220 280764 235272
rect 304908 235220 304960 235272
rect 317880 235220 317932 235272
rect 383384 235220 383436 235272
rect 502800 235220 502852 235272
rect 187608 235152 187660 235204
rect 169668 235084 169720 235136
rect 208400 235084 208452 235136
rect 179328 235016 179380 235068
rect 197268 235016 197320 235068
rect 236276 235152 236328 235204
rect 253940 235152 253992 235204
rect 259184 235152 259236 235204
rect 278136 235152 278188 235204
rect 306012 235152 306064 235204
rect 317788 235152 317840 235204
rect 381912 235152 381964 235204
rect 500868 235152 500920 235204
rect 236000 235084 236052 235136
rect 246948 235084 247000 235136
rect 247132 235084 247184 235136
rect 258540 235084 258592 235136
rect 262128 235084 262180 235136
rect 267280 235084 267332 235136
rect 267372 235084 267424 235136
rect 276756 235084 276808 235136
rect 305644 235084 305696 235136
rect 317696 235084 317748 235136
rect 379060 235084 379112 235136
rect 495348 235084 495400 235136
rect 161480 234948 161532 235000
rect 193036 234880 193088 234932
rect 198648 234880 198700 234932
rect 205732 234880 205784 234932
rect 208124 234948 208176 235000
rect 225788 234948 225840 235000
rect 248972 235016 249024 235068
rect 257988 235016 258040 235068
rect 274640 235016 274692 235068
rect 300676 235016 300728 235068
rect 306748 235016 306800 235068
rect 307024 235016 307076 235068
rect 320824 235016 320876 235068
rect 328828 235016 328880 235068
rect 343640 235016 343692 235068
rect 380808 235016 380860 235068
rect 489828 235016 489880 235068
rect 250812 234948 250864 235000
rect 263508 234948 263560 235000
rect 267464 234948 267516 235000
rect 304172 234948 304224 235000
rect 315396 234948 315448 235000
rect 323124 234948 323176 235000
rect 340788 234948 340840 235000
rect 376576 234948 376628 235000
rect 481548 234948 481600 235000
rect 212908 234880 212960 234932
rect 233148 234880 233200 234932
rect 236276 234880 236328 234932
rect 233240 234812 233292 234864
rect 249616 234880 249668 234932
rect 255504 234880 255556 234932
rect 273168 234880 273220 234932
rect 304540 234880 304592 234932
rect 315304 234880 315356 234932
rect 336280 234880 336332 234932
rect 336648 234880 336700 234932
rect 347044 234880 347096 234932
rect 347688 234880 347740 234932
rect 402612 234880 402664 234932
rect 413744 234880 413796 234932
rect 247040 234812 247092 234864
rect 255688 234812 255740 234864
rect 197176 234676 197228 234728
rect 210424 234744 210476 234796
rect 212540 234744 212592 234796
rect 217232 234744 217284 234796
rect 246948 234744 247000 234796
rect 208216 234676 208268 234728
rect 228640 234676 228692 234728
rect 244464 234676 244516 234728
rect 248604 234676 248656 234728
rect 252560 234744 252612 234796
rect 272800 234812 272852 234864
rect 297824 234812 297876 234864
rect 300860 234812 300912 234864
rect 309508 234812 309560 234864
rect 311716 234812 311768 234864
rect 312360 234812 312412 234864
rect 314016 234812 314068 234864
rect 315212 234812 315264 234864
rect 317144 234812 317196 234864
rect 320916 234812 320968 234864
rect 322848 234812 322900 234864
rect 324136 234812 324188 234864
rect 325516 234812 325568 234864
rect 326344 234812 326396 234864
rect 328184 234812 328236 234864
rect 328460 234812 328512 234864
rect 330852 234812 330904 234864
rect 331312 234812 331364 234864
rect 333796 234812 333848 234864
rect 343088 234812 343140 234864
rect 349068 234812 349120 234864
rect 386512 234812 386564 234864
rect 390560 234812 390612 234864
rect 267464 234744 267516 234796
rect 283196 234744 283248 234796
rect 296352 234744 296404 234796
rect 298192 234744 298244 234796
rect 307392 234744 307444 234796
rect 308956 234744 309008 234796
rect 309876 234744 309928 234796
rect 311808 234744 311860 234796
rect 313096 234744 313148 234796
rect 314476 234744 314528 234796
rect 315948 234744 316000 234796
rect 317328 234744 317380 234796
rect 318064 234744 318116 234796
rect 320088 234744 320140 234796
rect 321652 234744 321704 234796
rect 322756 234744 322808 234796
rect 324872 234744 324924 234796
rect 325608 234744 325660 234796
rect 326988 234744 327040 234796
rect 328276 234744 328328 234796
rect 329472 234744 329524 234796
rect 331128 234744 331180 234796
rect 332692 234744 332744 234796
rect 333888 234744 333940 234796
rect 337016 234744 337068 234796
rect 339224 234744 339276 234796
rect 339500 234744 339552 234796
rect 341800 234744 341852 234796
rect 342352 234744 342404 234796
rect 344376 234744 344428 234796
rect 345204 234744 345256 234796
rect 347136 234744 347188 234796
rect 347320 234744 347372 234796
rect 347688 234744 347740 234796
rect 348056 234744 348108 234796
rect 349896 234744 349948 234796
rect 350908 234744 350960 234796
rect 353024 234744 353076 234796
rect 353392 234744 353444 234796
rect 355784 234744 355836 234796
rect 356244 234744 356296 234796
rect 358544 234744 358596 234796
rect 359096 234744 359148 234796
rect 361212 234744 361264 234796
rect 384396 234744 384448 234796
rect 387800 234744 387852 234796
rect 42156 234608 42208 234660
rect 43260 234608 43312 234660
rect 215300 234608 215352 234660
rect 220084 234608 220136 234660
rect 241796 234608 241848 234660
rect 242900 234608 242952 234660
rect 246948 234608 247000 234660
rect 252836 234608 252888 234660
rect 253848 234676 253900 234728
rect 267372 234676 267424 234728
rect 267556 234676 267608 234728
rect 282460 234676 282512 234728
rect 292580 234676 292632 234728
rect 294604 234676 294656 234728
rect 295248 234676 295300 234728
rect 295892 234676 295944 234728
rect 296720 234676 296772 234728
rect 298284 234676 298336 234728
rect 298468 234676 298520 234728
rect 301044 234676 301096 234728
rect 308128 234676 308180 234728
rect 308864 234676 308916 234728
rect 310244 234676 310296 234728
rect 311440 234676 311492 234728
rect 312728 234676 312780 234728
rect 314108 234676 314160 234728
rect 314200 234676 314252 234728
rect 314568 234676 314620 234728
rect 316684 234676 316736 234728
rect 317236 234676 317288 234728
rect 318432 234676 318484 234728
rect 319904 234676 319956 234728
rect 321284 234676 321336 234728
rect 322480 234676 322532 234728
rect 323768 234676 323820 234728
rect 325332 234676 325384 234728
rect 327356 234676 327408 234728
rect 328368 234676 328420 234728
rect 330208 234676 330260 234728
rect 331036 234676 331088 234728
rect 332048 234676 332100 234728
rect 333520 234676 333572 234728
rect 334164 234676 334216 234728
rect 336096 234676 336148 234728
rect 337384 234676 337436 234728
rect 338856 234676 338908 234728
rect 340604 234676 340656 234728
rect 341984 234676 342036 234728
rect 343456 234676 343508 234728
rect 344652 234676 344704 234728
rect 346308 234676 346360 234728
rect 347596 234676 347648 234728
rect 349160 234676 349212 234728
rect 350264 234676 350316 234728
rect 350540 234676 350592 234728
rect 352564 234676 352616 234728
rect 353760 234676 353812 234728
rect 355416 234676 355468 234728
rect 356612 234676 356664 234728
rect 358084 234676 358136 234728
rect 359464 234676 359516 234728
rect 361396 234676 361448 234728
rect 362316 234676 362368 234728
rect 364064 234676 364116 234728
rect 375472 234676 375524 234728
rect 379428 234676 379480 234728
rect 384764 234676 384816 234728
rect 386236 234676 386288 234728
rect 387248 234676 387300 234728
rect 389088 234676 389140 234728
rect 398288 234676 398340 234728
rect 403808 234676 403860 234728
rect 411536 234676 411588 234728
rect 413836 234676 413888 234728
rect 262496 234608 262548 234660
rect 267648 234608 267700 234660
rect 282092 234608 282144 234660
rect 289820 234608 289872 234660
rect 292396 234608 292448 234660
rect 292672 234608 292724 234660
rect 293868 234608 293920 234660
rect 294972 234608 295024 234660
rect 295432 234608 295484 234660
rect 295800 234608 295852 234660
rect 297088 234608 297140 234660
rect 298836 234608 298888 234660
rect 300952 234608 301004 234660
rect 305276 234608 305328 234660
rect 306288 234608 306340 234660
rect 307760 234608 307812 234660
rect 308496 234608 308548 234660
rect 310980 234608 311032 234660
rect 311624 234608 311676 234660
rect 313832 234608 313884 234660
rect 314384 234608 314436 234660
rect 315580 234608 315632 234660
rect 316960 234608 317012 234660
rect 319536 234608 319588 234660
rect 319996 234608 320048 234660
rect 322388 234608 322440 234660
rect 322664 234608 322716 234660
rect 323492 234608 323544 234660
rect 325148 234608 325200 234660
rect 326620 234608 326672 234660
rect 327908 234608 327960 234660
rect 329840 234608 329892 234660
rect 330760 234608 330812 234660
rect 332324 234608 332376 234660
rect 333612 234608 333664 234660
rect 335544 234608 335596 234660
rect 336464 234608 336516 234660
rect 338028 234608 338080 234660
rect 338948 234608 339000 234660
rect 340236 234608 340288 234660
rect 341616 234608 341668 234660
rect 343732 234608 343784 234660
rect 344836 234608 344888 234660
rect 346584 234608 346636 234660
rect 347504 234608 347556 234660
rect 349436 234608 349488 234660
rect 350356 234608 350408 234660
rect 352012 234608 352064 234660
rect 352656 234608 352708 234660
rect 354864 234608 354916 234660
rect 355692 234608 355744 234660
rect 357716 234608 357768 234660
rect 358452 234608 358504 234660
rect 360568 234608 360620 234660
rect 361304 234608 361356 234660
rect 361948 234608 362000 234660
rect 363512 234608 363564 234660
rect 364800 234608 364852 234660
rect 367008 234608 367060 234660
rect 367652 234608 367704 234660
rect 369124 234608 369176 234660
rect 370504 234608 370556 234660
rect 371976 234608 372028 234660
rect 373356 234608 373408 234660
rect 374736 234608 374788 234660
rect 376944 234608 376996 234660
rect 377956 234608 378008 234660
rect 379796 234608 379848 234660
rect 380624 234608 380676 234660
rect 382280 234608 382332 234660
rect 384948 234608 385000 234660
rect 385132 234608 385184 234660
rect 386328 234608 386380 234660
rect 386880 234608 386932 234660
rect 388996 234608 389048 234660
rect 390100 234608 390152 234660
rect 391848 234608 391900 234660
rect 391940 234608 391992 234660
rect 403072 234608 403124 234660
rect 403624 234608 403676 234660
rect 407396 234608 407448 234660
rect 411904 234608 411956 234660
rect 413928 234608 413980 234660
rect 42156 234200 42208 234252
rect 43076 234200 43128 234252
rect 389732 233724 389784 233776
rect 401324 233724 401376 233776
rect 377680 233452 377732 233504
rect 489920 233452 489972 233504
rect 393688 233384 393740 233436
rect 528560 233384 528612 233436
rect 42156 233316 42208 233368
rect 43904 233316 43956 233368
rect 396908 233316 396960 233368
rect 536840 233316 536892 233368
rect 397920 233248 397972 233300
rect 539600 233248 539652 233300
rect 287244 233180 287296 233232
rect 287888 233180 287940 233232
rect 400128 233180 400180 233232
rect 542452 233180 542504 233232
rect 284392 233112 284444 233164
rect 285036 233112 285088 233164
rect 287060 233112 287112 233164
rect 287612 233112 287664 233164
rect 193680 233044 193732 233096
rect 195520 233044 195572 233096
rect 196164 233044 196216 233096
rect 198372 233044 198424 233096
rect 226616 233044 226668 233096
rect 227628 233044 227680 233096
rect 229284 233044 229336 233096
rect 230480 233044 230532 233096
rect 232044 233044 232096 233096
rect 233332 233044 233384 233096
rect 234804 233044 234856 233096
rect 236184 233044 236236 233096
rect 240324 233044 240376 233096
rect 241888 233044 241940 233096
rect 243084 233044 243136 233096
rect 244740 233044 244792 233096
rect 245844 233044 245896 233096
rect 247592 233044 247644 233096
rect 251364 233044 251416 233096
rect 253296 233044 253348 233096
rect 281724 233044 281776 233096
rect 283288 233044 283340 233096
rect 290280 233044 290332 233096
rect 291108 233044 291160 233096
rect 190644 232976 190696 233028
rect 192392 232976 192444 233028
rect 193496 232976 193548 233028
rect 194876 232976 194928 233028
rect 196348 232976 196400 233028
rect 198096 232976 198148 233028
rect 218428 232976 218480 233028
rect 220176 232976 220228 233028
rect 221096 232976 221148 233028
rect 221924 232976 221976 233028
rect 223764 232976 223816 233028
rect 224776 232976 224828 233028
rect 226800 232976 226852 233028
rect 227260 232976 227312 233028
rect 229192 232976 229244 233028
rect 230112 232976 230164 233028
rect 232320 232976 232372 233028
rect 232964 232976 233016 233028
rect 235172 232976 235224 233028
rect 235816 232976 235868 233028
rect 237748 232976 237800 233028
rect 238668 232976 238720 233028
rect 240508 232976 240560 233028
rect 241520 232976 241572 233028
rect 243268 232976 243320 233028
rect 244372 232976 244424 233028
rect 246028 232976 246080 233028
rect 247224 232976 247276 233028
rect 248604 232976 248656 233028
rect 250444 232976 250496 233028
rect 251456 232976 251508 233028
rect 252928 232976 252980 233028
rect 254216 232976 254268 233028
rect 255780 232976 255832 233028
rect 257068 232976 257120 233028
rect 258632 232976 258684 233028
rect 259828 232976 259880 233028
rect 261484 232976 261536 233028
rect 262588 232976 262640 233028
rect 264336 232976 264388 233028
rect 268200 232976 268252 233028
rect 270040 232976 270092 233028
rect 282000 232976 282052 233028
rect 283656 232976 283708 233028
rect 284484 232976 284536 233028
rect 286508 232976 286560 233028
rect 287888 232976 287940 233028
rect 289360 232976 289412 233028
rect 290372 232976 290424 233028
rect 291476 232976 291528 233028
rect 292764 232976 292816 233028
rect 293960 232976 294012 233028
rect 196440 232908 196492 232960
rect 197728 232908 197780 232960
rect 237656 232908 237708 232960
rect 239036 232908 239088 232960
rect 281816 232908 281868 232960
rect 283932 232908 283984 232960
rect 287428 232908 287480 232960
rect 288624 232908 288676 232960
rect 290188 232908 290240 232960
rect 291844 232908 291896 232960
rect 314016 232908 314068 232960
rect 314476 232908 314528 232960
rect 335452 232908 335504 232960
rect 336372 232908 336424 232960
rect 196256 232840 196308 232892
rect 196624 232840 196676 232892
rect 287152 232840 287204 232892
rect 288256 232840 288308 232892
rect 284852 232636 284904 232688
rect 286140 232636 286192 232688
rect 341708 231752 341760 231804
rect 403624 231752 403676 231804
rect 363052 231684 363104 231736
rect 454132 231684 454184 231736
rect 364432 231616 364484 231668
rect 457444 231616 457496 231668
rect 367284 231548 367336 231600
rect 464252 231548 464304 231600
rect 287796 231480 287848 231532
rect 288992 231480 289044 231532
rect 365904 231480 365956 231532
rect 460940 231480 460992 231532
rect 370136 231412 370188 231464
rect 470968 231412 471020 231464
rect 368756 231344 368808 231396
rect 467564 231344 467616 231396
rect 371608 231276 371660 231328
rect 474280 231276 474332 231328
rect 372988 231208 373040 231260
rect 477684 231208 477736 231260
rect 374460 231140 374512 231192
rect 480996 231140 481048 231192
rect 42156 231072 42208 231124
rect 43628 231072 43680 231124
rect 374552 231072 374604 231124
rect 483020 231072 483072 231124
rect 186412 231004 186464 231056
rect 248236 231004 248288 231056
rect 376208 231004 376260 231056
rect 487160 231004 487212 231056
rect 179696 230936 179748 230988
rect 245384 230936 245436 230988
rect 389364 230936 389416 230988
rect 183100 230868 183152 230920
rect 246764 230868 246816 230920
rect 390468 230868 390520 230920
rect 401600 230936 401652 230988
rect 515496 230936 515548 230988
rect 172980 230800 173032 230852
rect 242532 230800 242584 230852
rect 391572 230800 391624 230852
rect 518072 230868 518124 230920
rect 176384 230732 176436 230784
rect 243912 230732 243964 230784
rect 518992 230800 519044 230852
rect 523408 230732 523460 230784
rect 166264 230664 166316 230716
rect 239680 230664 239732 230716
rect 334900 230664 334952 230716
rect 389364 230664 389416 230716
rect 392584 230664 392636 230716
rect 525892 230664 525944 230716
rect 169576 230596 169628 230648
rect 241060 230596 241112 230648
rect 336648 230596 336700 230648
rect 392676 230596 392728 230648
rect 394792 230596 394844 230648
rect 530952 230596 531004 230648
rect 42156 230528 42208 230580
rect 42984 230528 43036 230580
rect 162768 230528 162820 230580
rect 238208 230528 238260 230580
rect 337752 230528 337804 230580
rect 395712 230528 395764 230580
rect 395804 230528 395856 230580
rect 533160 230528 533212 230580
rect 46848 230460 46900 230512
rect 662880 230460 662932 230512
rect 46388 230392 46440 230444
rect 662788 230392 662840 230444
rect 339408 230324 339460 230376
rect 399484 230324 399536 230376
rect 388352 230256 388404 230308
rect 401600 230256 401652 230308
rect 42156 229848 42208 229900
rect 43168 229848 43220 229900
rect 42156 229032 42208 229084
rect 43536 229032 43588 229084
rect 353116 229032 353168 229084
rect 428924 229032 428976 229084
rect 159548 228964 159600 229016
rect 236828 228964 236880 229016
rect 354128 228964 354180 229016
rect 432236 228964 432288 229016
rect 156144 228896 156196 228948
rect 235356 228896 235408 228948
rect 355508 228896 355560 228948
rect 435640 228896 435692 228948
rect 152832 228828 152884 228880
rect 233976 228828 234028 228880
rect 354496 228828 354548 228880
rect 433892 228828 433944 228880
rect 149428 228760 149480 228812
rect 232504 228760 232556 228812
rect 353208 228760 353260 228812
rect 430580 228760 430632 228812
rect 146024 228692 146076 228744
rect 231124 228692 231176 228744
rect 357348 228692 357400 228744
rect 440700 228692 440752 228744
rect 142712 228624 142764 228676
rect 229652 228624 229704 228676
rect 355876 228624 355928 228676
rect 437296 228624 437348 228676
rect 139216 228556 139268 228608
rect 228272 228556 228324 228608
rect 356980 228556 357032 228608
rect 438952 228556 439004 228608
rect 135996 228488 136048 228540
rect 226708 228488 226760 228540
rect 358360 228488 358412 228540
rect 442356 228488 442408 228540
rect 132408 228420 132460 228472
rect 225420 228420 225472 228472
rect 359832 228420 359884 228472
rect 445668 228420 445720 228472
rect 129280 228352 129332 228404
rect 223948 228352 224000 228404
rect 358728 228352 358780 228404
rect 444380 228352 444432 228404
rect 125876 228284 125928 228336
rect 222568 228284 222620 228336
rect 360200 228284 360252 228336
rect 447416 228284 447468 228336
rect 122472 228216 122524 228268
rect 221188 228216 221240 228268
rect 361488 228216 361540 228268
rect 449072 228216 449124 228268
rect 119160 228148 119212 228200
rect 219716 228148 219768 228200
rect 361580 228148 361632 228200
rect 450728 228148 450780 228200
rect 97264 228080 97316 228132
rect 210792 228080 210844 228132
rect 248788 228080 248840 228132
rect 250076 228080 250128 228132
rect 362684 228080 362736 228132
rect 452660 228080 452712 228132
rect 93768 228012 93820 228064
rect 209412 228012 209464 228064
rect 221740 228012 221792 228064
rect 263600 228012 263652 228064
rect 365536 228012 365588 228064
rect 459192 228012 459244 228064
rect 87144 227944 87196 227996
rect 206560 227944 206612 227996
rect 218336 227944 218388 227996
rect 261852 227944 261904 227996
rect 364248 227944 364300 227996
rect 455788 227944 455840 227996
rect 90548 227876 90600 227928
rect 207940 227876 207992 227928
rect 215024 227876 215076 227928
rect 260472 227876 260524 227928
rect 363972 227876 364024 227928
rect 458364 227876 458416 227928
rect 61936 227808 61988 227860
rect 195428 227808 195480 227860
rect 211712 227808 211764 227860
rect 259000 227808 259052 227860
rect 368388 227808 368440 227860
rect 465908 227808 465960 227860
rect 58624 227740 58676 227792
rect 194048 227740 194100 227792
rect 204904 227740 204956 227792
rect 256424 227740 256476 227792
rect 365168 227740 365220 227792
rect 461676 227740 461728 227792
rect 53564 227672 53616 227724
rect 192300 227672 192352 227724
rect 208492 227672 208544 227724
rect 257896 227672 257948 227724
rect 366916 227672 366968 227724
rect 462504 227672 462556 227724
rect 349804 227604 349856 227656
rect 422300 227604 422352 227656
rect 351644 227536 351696 227588
rect 427176 227536 427228 227588
rect 350172 227468 350224 227520
rect 423864 227468 423916 227520
rect 42064 227400 42116 227452
rect 43352 227400 43404 227452
rect 351276 227400 351328 227452
rect 425520 227400 425572 227452
rect 348792 227332 348844 227384
rect 420460 227332 420512 227384
rect 347688 227264 347740 227316
rect 417148 227264 417200 227316
rect 345940 227196 345992 227248
rect 414020 227196 414072 227248
rect 290004 227128 290056 227180
rect 290740 227128 290792 227180
rect 348424 227128 348476 227180
rect 418804 227128 418856 227180
rect 346952 227060 347004 227112
rect 415400 227060 415452 227112
rect 344468 226992 344520 227044
rect 410340 226992 410392 227044
rect 345572 226924 345624 226976
rect 412088 226924 412140 226976
rect 344100 226856 344152 226908
rect 408684 226856 408736 226908
rect 42156 226788 42208 226840
rect 43812 226788 43864 226840
rect 342996 226788 343048 226840
rect 405740 226788 405792 226840
rect 341248 226720 341300 226772
rect 401968 226720 402020 226772
rect 339868 226652 339920 226704
rect 398564 226652 398616 226704
rect 137652 226244 137704 226296
rect 226616 226244 226668 226296
rect 349896 226244 349948 226296
rect 421288 226244 421340 226296
rect 134248 226176 134300 226228
rect 226524 226176 226576 226228
rect 347412 226176 347464 226228
rect 418252 226176 418304 226228
rect 130936 226108 130988 226160
rect 223764 226108 223816 226160
rect 347044 226108 347096 226160
rect 419724 226108 419776 226160
rect 127532 226040 127584 226092
rect 223856 226040 223908 226092
rect 352564 226040 352616 226092
rect 426348 226040 426400 226092
rect 124128 225972 124180 226024
rect 221096 225972 221148 226024
rect 350264 225972 350316 226024
rect 423036 225972 423088 226024
rect 114100 225904 114152 225956
rect 217600 225904 217652 225956
rect 352656 225904 352708 225956
rect 429752 225904 429804 225956
rect 117504 225836 117556 225888
rect 219072 225836 219124 225888
rect 353024 225836 353076 225888
rect 428004 225836 428056 225888
rect 120816 225768 120868 225820
rect 221004 225768 221056 225820
rect 350356 225768 350408 225820
rect 425060 225768 425112 225820
rect 110696 225700 110748 225752
rect 216220 225700 216272 225752
rect 355784 225700 355836 225752
rect 433340 225700 433392 225752
rect 115756 225632 115808 225684
rect 218244 225632 218296 225684
rect 355416 225632 355468 225684
rect 434812 225632 434864 225684
rect 112444 225564 112496 225616
rect 216588 225564 216640 225616
rect 352932 225564 352984 225616
rect 431408 225564 431460 225616
rect 109040 225496 109092 225548
rect 215668 225496 215720 225548
rect 355324 225496 355376 225548
rect 438124 225496 438176 225548
rect 105728 225428 105780 225480
rect 213736 225428 213788 225480
rect 358544 225428 358596 225480
rect 439780 225428 439832 225480
rect 107384 225360 107436 225412
rect 214840 225360 214892 225412
rect 355692 225360 355744 225412
rect 436468 225360 436520 225412
rect 100668 225292 100720 225344
rect 211988 225292 212040 225344
rect 228456 225292 228508 225344
rect 266176 225292 266228 225344
rect 358084 225292 358136 225344
rect 441620 225292 441672 225344
rect 103980 225224 104032 225276
rect 213368 225224 213420 225276
rect 231768 225224 231820 225276
rect 267832 225224 267884 225276
rect 361212 225224 361264 225276
rect 446588 225224 446640 225276
rect 95608 225156 95660 225208
rect 209504 225156 209556 225208
rect 225144 225156 225196 225208
rect 265256 225156 265308 225208
rect 358452 225156 358504 225208
rect 443184 225156 443236 225208
rect 73712 225088 73764 225140
rect 200580 225088 200632 225140
rect 201316 225088 201368 225140
rect 254768 225088 254820 225140
rect 358176 225088 358228 225140
rect 444840 225088 444892 225140
rect 66996 225020 67048 225072
rect 196440 225020 196492 225072
rect 198188 225020 198240 225072
rect 251364 225020 251416 225072
rect 361396 225020 361448 225072
rect 448244 225020 448296 225072
rect 60280 224952 60332 225004
rect 193496 224952 193548 225004
rect 194876 224952 194928 225004
rect 251916 224952 251968 225004
rect 363512 224952 363564 225004
rect 453304 224952 453356 225004
rect 55128 224884 55180 224936
rect 190644 224884 190696 224936
rect 191472 224884 191524 224936
rect 248604 224884 248656 224936
rect 361304 224884 361356 224936
rect 449900 224884 449952 224936
rect 141056 224816 141108 224868
rect 229376 224816 229428 224868
rect 347596 224816 347648 224868
rect 416228 224816 416280 224868
rect 144368 224748 144420 224800
rect 229284 224748 229336 224800
rect 344836 224748 344888 224800
rect 411260 224748 411312 224800
rect 147772 224680 147824 224732
rect 232136 224680 232188 224732
rect 344744 224680 344796 224732
rect 412916 224680 412968 224732
rect 154488 224612 154540 224664
rect 234896 224612 234948 224664
rect 347136 224612 347188 224664
rect 414572 224612 414624 224664
rect 151084 224544 151136 224596
rect 232044 224544 232096 224596
rect 344652 224544 344704 224596
rect 409512 224544 409564 224596
rect 161204 224476 161256 224528
rect 237564 224476 237616 224528
rect 341892 224476 341944 224528
rect 406200 224476 406252 224528
rect 704004 224476 704056 224528
rect 708880 224476 708932 224528
rect 157800 224408 157852 224460
rect 234804 224408 234856 224460
rect 341984 224408 342036 224460
rect 402980 224408 403032 224460
rect 704464 224408 704516 224460
rect 708420 224408 708472 224460
rect 164608 224340 164660 224392
rect 237656 224340 237708 224392
rect 341156 224340 341208 224392
rect 404452 224340 404504 224392
rect 167920 224272 167972 224324
rect 240600 224272 240652 224324
rect 344376 224272 344428 224324
rect 407856 224272 407908 224324
rect 707500 224340 707552 224392
rect 707040 224272 707092 224324
rect 171048 224204 171100 224256
rect 240324 224204 240376 224256
rect 336280 224204 336332 224256
rect 394700 224204 394752 224256
rect 705292 224204 705344 224256
rect 705752 224204 705804 224256
rect 706212 224204 706264 224256
rect 706580 224204 706632 224256
rect 174636 224136 174688 224188
rect 243452 224136 243504 224188
rect 339132 224136 339184 224188
rect 397736 224136 397788 224188
rect 705844 224136 705896 224188
rect 707040 224136 707092 224188
rect 178040 224068 178092 224120
rect 243084 224068 243136 224120
rect 341800 224068 341852 224120
rect 401140 224068 401192 224120
rect 706304 224068 706356 224120
rect 706580 224068 706632 224120
rect 181352 224000 181404 224052
rect 246212 224000 246264 224052
rect 336372 224000 336424 224052
rect 391020 224000 391072 224052
rect 705384 224000 705436 224052
rect 707500 224000 707552 224052
rect 708052 224000 708104 224052
rect 184756 223932 184808 223984
rect 245844 223932 245896 223984
rect 333428 223932 333480 223984
rect 385960 223932 386012 223984
rect 704924 223932 704976 223984
rect 707960 223932 708012 223984
rect 188160 223864 188212 223916
rect 249064 223864 249116 223916
rect 333520 223864 333572 223916
rect 382648 223864 382700 223916
rect 704832 223864 704884 223916
rect 113088 223524 113140 223576
rect 139308 223524 139360 223576
rect 141884 223524 141936 223576
rect 229192 223524 229244 223576
rect 272248 223524 272300 223576
rect 284576 223524 284628 223576
rect 325516 223524 325568 223576
rect 361764 223524 361816 223576
rect 494336 223524 494388 223576
rect 495348 223524 495400 223576
rect 607588 223524 607640 223576
rect 108212 223456 108264 223508
rect 136548 223456 136600 223508
rect 140136 223456 140188 223508
rect 229744 223456 229796 223508
rect 230940 223456 230992 223508
rect 244280 223456 244332 223508
rect 244464 223456 244516 223508
rect 273076 223456 273128 223508
rect 284760 223456 284812 223508
rect 325148 223456 325200 223508
rect 362408 223456 362460 223508
rect 499488 223456 499540 223508
rect 608048 223456 608100 223508
rect 106556 223388 106608 223440
rect 125508 223388 125560 223440
rect 135168 223388 135220 223440
rect 226800 223388 226852 223440
rect 227536 223388 227588 223440
rect 278688 223388 278740 223440
rect 287336 223388 287388 223440
rect 314200 223388 314252 223440
rect 339684 223388 339736 223440
rect 346216 223388 346268 223440
rect 383660 223388 383712 223440
rect 403808 223388 403860 223440
rect 539048 223388 539100 223440
rect 546040 223388 546092 223440
rect 616880 223388 616932 223440
rect 86316 223320 86368 223372
rect 128268 223320 128320 223372
rect 101496 223252 101548 223304
rect 122748 223252 122800 223304
rect 128360 223252 128412 223304
rect 199016 223320 199068 223372
rect 224132 223320 224184 223372
rect 229284 223320 229336 223372
rect 244188 223320 244240 223372
rect 244464 223320 244516 223372
rect 255320 223320 255372 223372
rect 278136 223320 278188 223372
rect 287152 223320 287204 223372
rect 328184 223320 328236 223372
rect 369124 223320 369176 223372
rect 500868 223320 500920 223372
rect 608508 223320 608560 223372
rect 224040 223252 224092 223304
rect 241152 223252 241204 223304
rect 252560 223252 252612 223304
rect 328276 223252 328328 223304
rect 368296 223252 368348 223304
rect 394516 223252 394568 223304
rect 530032 223252 530084 223304
rect 538864 223252 538916 223304
rect 539600 223252 539652 223304
rect 78772 223184 78824 223236
rect 119988 223184 120040 223236
rect 126704 223184 126756 223236
rect 198832 223184 198884 223236
rect 198924 223184 198976 223236
rect 207940 223184 207992 223236
rect 94780 223116 94832 223168
rect 111708 223116 111760 223168
rect 116584 223116 116636 223168
rect 215300 223184 215352 223236
rect 221280 223184 221332 223236
rect 237748 223184 237800 223236
rect 252468 223184 252520 223236
rect 325608 223184 325660 223236
rect 365812 223184 365864 223236
rect 398656 223184 398708 223236
rect 539876 223184 539928 223236
rect 542452 223184 542504 223236
rect 543648 223184 543700 223236
rect 546960 223252 547012 223304
rect 615040 223252 615092 223304
rect 72056 223048 72108 223100
rect 117228 223048 117280 223100
rect 119988 223048 120040 223100
rect 220084 223116 220136 223168
rect 235908 223116 235960 223168
rect 242716 223116 242768 223168
rect 255504 223116 255556 223168
rect 308956 223116 309008 223168
rect 323124 223116 323176 223168
rect 325424 223116 325476 223168
rect 364984 223116 365036 223168
rect 406384 223116 406436 223168
rect 546684 223116 546736 223168
rect 615500 223184 615552 223236
rect 616420 223116 616472 223168
rect 88064 222980 88116 223032
rect 106188 222980 106240 223032
rect 118332 222980 118384 223032
rect 218428 223048 218480 223100
rect 226616 223048 226668 223100
rect 230940 223048 230992 223100
rect 231032 223048 231084 223100
rect 249892 223048 249944 223100
rect 311716 223048 311768 223100
rect 330484 223048 330536 223100
rect 330852 223048 330904 223100
rect 371700 223048 371752 223100
rect 400036 223048 400088 223100
rect 542176 223048 542228 223100
rect 542360 223048 542412 223100
rect 615960 223048 616012 223100
rect 224316 222980 224368 223032
rect 250168 222980 250220 223032
rect 308772 222980 308824 223032
rect 323768 222980 323820 223032
rect 325332 222980 325384 223032
rect 364340 222980 364392 223032
rect 401876 222980 401928 223032
rect 544936 222980 544988 223032
rect 545120 222980 545172 223032
rect 546040 222980 546092 223032
rect 65340 222912 65392 222964
rect 103428 222912 103480 222964
rect 109868 222912 109920 222964
rect 198924 222912 198976 222964
rect 199016 222912 199068 222964
rect 201408 222912 201460 222964
rect 207940 222912 207992 222964
rect 212540 222912 212592 222964
rect 229376 222912 229428 222964
rect 82728 222844 82780 222896
rect 97908 222844 97960 222896
rect 103152 222844 103204 222896
rect 214104 222844 214156 222896
rect 214196 222844 214248 222896
rect 236092 222912 236144 222964
rect 268200 222912 268252 222964
rect 317236 222912 317288 222964
rect 347320 222912 347372 222964
rect 347412 222912 347464 222964
rect 386788 222912 386840 222964
rect 402520 222912 402572 222964
rect 536288 222912 536340 222964
rect 536380 222912 536432 222964
rect 536840 222912 536892 222964
rect 546960 222912 547012 222964
rect 550548 222912 550600 222964
rect 551468 222912 551520 222964
rect 617800 222912 617852 222964
rect 98092 222776 98144 222828
rect 211620 222776 211672 222828
rect 215852 222776 215904 222828
rect 235816 222776 235868 222828
rect 263508 222844 263560 222896
rect 309048 222844 309100 222896
rect 326252 222844 326304 222896
rect 328368 222844 328420 222896
rect 370044 222844 370096 222896
rect 407396 222844 407448 222896
rect 552020 222844 552072 222896
rect 247316 222776 247368 222828
rect 308680 222776 308732 222828
rect 324596 222776 324648 222828
rect 325240 222776 325292 222828
rect 367468 222776 367520 222828
rect 405832 222776 405884 222828
rect 62764 222708 62816 222760
rect 89628 222708 89680 222760
rect 189540 222708 189592 222760
rect 205180 222708 205232 222760
rect 207388 222708 207440 222760
rect 247132 222708 247184 222760
rect 281448 222708 281500 222760
rect 289912 222708 289964 222760
rect 308864 222708 308916 222760
rect 327080 222708 327132 222760
rect 327908 222708 327960 222760
rect 370872 222708 370924 222760
rect 404360 222708 404412 222760
rect 552204 222708 552256 222760
rect 555056 222708 555108 222760
rect 71228 222640 71280 222692
rect 81348 222640 81400 222692
rect 89720 222640 89772 222692
rect 208400 222640 208452 222692
rect 222568 222640 222620 222692
rect 262588 222640 262640 222692
rect 311440 222640 311492 222692
rect 329656 222640 329708 222692
rect 333796 222640 333848 222692
rect 378416 222640 378468 222692
rect 403992 222640 404044 222692
rect 552112 222640 552164 222692
rect 82176 222572 82228 222624
rect 203800 222572 203852 222624
rect 209136 222572 209188 222624
rect 85488 222504 85540 222556
rect 189540 222504 189592 222556
rect 81256 222436 81308 222488
rect 204444 222504 204496 222556
rect 212356 222504 212408 222556
rect 235816 222572 235868 222624
rect 259828 222572 259880 222624
rect 308496 222572 308548 222624
rect 325700 222572 325752 222624
rect 328000 222572 328052 222624
rect 372620 222572 372672 222624
rect 406292 222572 406344 222624
rect 557908 222844 557960 222896
rect 564072 222844 564124 222896
rect 559104 222776 559156 222828
rect 572812 222776 572864 222828
rect 189724 222436 189776 222488
rect 208768 222436 208820 222488
rect 213368 222436 213420 222488
rect 220820 222436 220872 222488
rect 257068 222504 257120 222556
rect 311532 222504 311584 222556
rect 332968 222504 333020 222556
rect 333888 222504 333940 222556
rect 381820 222504 381872 222556
rect 406476 222504 406528 222556
rect 561680 222708 561732 222760
rect 619640 222708 619692 222760
rect 556068 222640 556120 222692
rect 618720 222640 618772 222692
rect 260104 222436 260156 222488
rect 311348 222436 311400 222488
rect 331312 222436 331364 222488
rect 336096 222436 336148 222488
rect 385132 222436 385184 222488
rect 408776 222436 408828 222488
rect 563980 222572 564032 222624
rect 564072 222572 564124 222624
rect 633624 222572 633676 222624
rect 561588 222504 561640 222556
rect 634084 222504 634136 222556
rect 555424 222436 555476 222488
rect 562876 222436 562928 222488
rect 563980 222436 564032 222488
rect 620100 222436 620152 222488
rect 56048 222368 56100 222420
rect 73068 222368 73120 222420
rect 75368 222368 75420 222420
rect 200948 222368 201000 222420
rect 205824 222368 205876 222420
rect 257344 222368 257396 222420
rect 283196 222368 283248 222420
rect 290096 222368 290148 222420
rect 314108 222368 314160 222420
rect 334716 222368 334768 222420
rect 336464 222368 336516 222420
rect 388536 222368 388588 222420
rect 408132 222368 408184 222420
rect 561772 222368 561824 222420
rect 202420 222300 202472 222352
rect 254216 222300 254268 222352
rect 311624 222300 311676 222352
rect 333980 222300 334032 222352
rect 338856 222300 338908 222352
rect 393596 222300 393648 222352
rect 408224 222300 408276 222352
rect 555424 222300 555476 222352
rect 570236 222368 570288 222420
rect 194048 222232 194100 222284
rect 246948 222232 247000 222284
rect 314292 222232 314344 222284
rect 338028 222232 338080 222284
rect 339224 222232 339276 222284
rect 391940 222232 391992 222284
rect 413836 222232 413888 222284
rect 569960 222300 570012 222352
rect 621020 222300 621072 222352
rect 54392 222164 54444 222216
rect 193312 222164 193364 222216
rect 195704 222164 195756 222216
rect 251456 222164 251508 222216
rect 317052 222164 317104 222216
rect 345020 222164 345072 222216
rect 349068 222164 349120 222216
rect 407028 222164 407080 222216
rect 409696 222164 409748 222216
rect 566004 222232 566056 222284
rect 555700 222164 555752 222216
rect 556160 222164 556212 222216
rect 114928 222096 114980 222148
rect 142160 222096 142212 222148
rect 148600 222096 148652 222148
rect 232320 222096 232372 222148
rect 280620 222096 280672 222148
rect 287244 222096 287296 222148
rect 322664 222096 322716 222148
rect 360752 222096 360804 222148
rect 401416 222096 401468 222148
rect 529020 222096 529072 222148
rect 536288 222096 536340 222148
rect 548340 222096 548392 222148
rect 560760 222096 560812 222148
rect 561588 222096 561640 222148
rect 569132 222096 569184 222148
rect 569960 222096 570012 222148
rect 620560 222164 620612 222216
rect 652852 222164 652904 222216
rect 633164 222096 633216 222148
rect 674564 222164 674616 222216
rect 675760 222164 675812 222216
rect 674656 222096 674708 222148
rect 675576 222096 675628 222148
rect 146944 222028 146996 222080
rect 232596 222028 232648 222080
rect 233516 222028 233568 222080
rect 248788 222028 248840 222080
rect 322572 222028 322624 222080
rect 358268 222028 358320 222080
rect 389088 222028 389140 222080
rect 513380 222028 513432 222080
rect 544936 222028 544988 222080
rect 547512 222028 547564 222080
rect 552112 222028 552164 222080
rect 552848 222028 552900 222080
rect 632704 222028 632756 222080
rect 153660 221960 153712 222012
rect 235448 221960 235500 222012
rect 274732 221960 274784 222012
rect 287612 221960 287664 222012
rect 322756 221960 322808 222012
rect 356520 221960 356572 222012
rect 386328 221960 386380 222012
rect 507952 221960 508004 222012
rect 533160 221960 533212 222012
rect 533804 221960 533856 222012
rect 614580 221960 614632 222012
rect 93032 221892 93084 221944
rect 153108 221892 153160 221944
rect 155316 221892 155368 221944
rect 235172 221892 235224 221944
rect 319996 221892 320048 221944
rect 354036 221892 354088 221944
rect 390560 221892 390612 221944
rect 511356 221892 511408 221944
rect 530952 221892 531004 221944
rect 614028 221892 614080 221944
rect 123392 221824 123444 221876
rect 155960 221824 156012 221876
rect 160376 221824 160428 221876
rect 125048 221756 125100 221808
rect 156052 221756 156104 221808
rect 162032 221756 162084 221808
rect 232228 221756 232280 221808
rect 99840 221688 99892 221740
rect 161480 221688 161532 221740
rect 170496 221688 170548 221740
rect 234344 221824 234396 221876
rect 249708 221824 249760 221876
rect 275560 221824 275612 221876
rect 284852 221824 284904 221876
rect 322848 221824 322900 221876
rect 357348 221824 357400 221876
rect 383568 221824 383620 221876
rect 503536 221824 503588 221876
rect 541440 221824 541492 221876
rect 542360 221824 542412 221876
rect 547512 221824 547564 221876
rect 631784 221824 631836 221876
rect 232504 221756 232556 221808
rect 237656 221756 237708 221808
rect 317144 221756 317196 221808
rect 343916 221756 343968 221808
rect 346400 221756 346452 221808
rect 380072 221756 380124 221808
rect 403072 221756 403124 221808
rect 523960 221756 524012 221808
rect 528560 221756 528612 221808
rect 613568 221756 613620 221808
rect 130108 221620 130160 221672
rect 158628 221620 158680 221672
rect 168748 221620 168800 221672
rect 232228 221620 232280 221672
rect 143448 221552 143500 221604
rect 169668 221552 169720 221604
rect 175464 221552 175516 221604
rect 232136 221552 232188 221604
rect 238300 221688 238352 221740
rect 322480 221688 322532 221740
rect 354864 221688 354916 221740
rect 401324 221688 401376 221740
rect 518900 221688 518952 221740
rect 545028 221688 545080 221740
rect 631324 221688 631376 221740
rect 232412 221620 232464 221672
rect 240508 221620 240560 221672
rect 279792 221620 279844 221672
rect 287428 221620 287480 221672
rect 319812 221620 319864 221672
rect 351460 221620 351512 221672
rect 387800 221620 387852 221672
rect 506296 221620 506348 221672
rect 525892 221620 525944 221672
rect 613108 221620 613160 221672
rect 241612 221552 241664 221604
rect 276480 221552 276532 221604
rect 287060 221552 287112 221604
rect 320088 221552 320140 221604
rect 350632 221552 350684 221604
rect 380808 221552 380860 221604
rect 497372 221552 497424 221604
rect 499488 221552 499540 221604
rect 136824 221484 136876 221536
rect 161572 221484 161624 221536
rect 177212 221484 177264 221536
rect 229284 221484 229336 221536
rect 229560 221484 229612 221536
rect 236000 221484 236052 221536
rect 236920 221484 236972 221536
rect 241520 221484 241572 221536
rect 246120 221484 246172 221536
rect 257988 221484 258040 221536
rect 314384 221484 314436 221536
rect 340604 221484 340656 221536
rect 343732 221484 343784 221536
rect 373356 221484 373408 221536
rect 384948 221484 385000 221536
rect 501236 221484 501288 221536
rect 182088 221416 182140 221468
rect 57704 221348 57756 221400
rect 62028 221348 62080 221400
rect 76288 221348 76340 221400
rect 78588 221348 78640 221400
rect 138480 221348 138532 221400
rect 147588 221348 147640 221400
rect 52736 221280 52788 221332
rect 67548 221280 67600 221332
rect 77944 221280 77996 221332
rect 86868 221280 86920 221332
rect 131764 221280 131816 221332
rect 142068 221280 142120 221332
rect 145196 221280 145248 221332
rect 150348 221348 150400 221400
rect 151728 221348 151780 221400
rect 155868 221348 155920 221400
rect 158720 221348 158772 221400
rect 159824 221348 159876 221400
rect 163688 221348 163740 221400
rect 165344 221348 165396 221400
rect 172152 221348 172204 221400
rect 173808 221348 173860 221400
rect 183928 221348 183980 221400
rect 227536 221348 227588 221400
rect 227628 221348 227680 221400
rect 229008 221348 229060 221400
rect 246028 221416 246080 221468
rect 249524 221416 249576 221468
rect 258172 221416 258224 221468
rect 271420 221416 271472 221468
rect 284668 221416 284720 221468
rect 317328 221416 317380 221468
rect 232136 221348 232188 221400
rect 150256 221280 150308 221332
rect 153200 221280 153252 221332
rect 156972 221280 157024 221332
rect 161388 221280 161440 221332
rect 167092 221280 167144 221332
rect 168104 221280 168156 221332
rect 178868 221280 178920 221332
rect 179328 221280 179380 221332
rect 185584 221280 185636 221332
rect 187608 221280 187660 221332
rect 192300 221280 192352 221332
rect 192944 221280 192996 221332
rect 196532 221280 196584 221332
rect 200856 221280 200908 221332
rect 208032 221280 208084 221332
rect 233516 221280 233568 221332
rect 235264 221348 235316 221400
rect 237288 221348 237340 221400
rect 243268 221348 243320 221400
rect 247040 221348 247092 221400
rect 248328 221348 248380 221400
rect 254584 221348 254636 221400
rect 256516 221348 256568 221400
rect 257068 221348 257120 221400
rect 259184 221348 259236 221400
rect 289728 221348 289780 221400
rect 292948 221348 293000 221400
rect 298100 221348 298152 221400
rect 299388 221348 299440 221400
rect 300952 221348 301004 221400
rect 302700 221348 302752 221400
rect 309784 221348 309836 221400
rect 311164 221348 311216 221400
rect 315028 221348 315080 221400
rect 315488 221348 315540 221400
rect 317788 221348 317840 221400
rect 319536 221348 319588 221400
rect 319904 221416 319956 221468
rect 348148 221416 348200 221468
rect 379428 221416 379480 221468
rect 484400 221416 484452 221468
rect 513380 221416 513432 221468
rect 343088 221348 343140 221400
rect 343640 221348 343692 221400
rect 366640 221348 366692 221400
rect 387616 221348 387668 221400
rect 491300 221348 491352 221400
rect 507952 221348 508004 221400
rect 536748 221552 536800 221604
rect 538036 221552 538088 221604
rect 539508 221484 539560 221536
rect 541624 221484 541676 221536
rect 542268 221484 542320 221536
rect 544108 221484 544160 221536
rect 547788 221484 547840 221536
rect 549260 221484 549312 221536
rect 552296 221484 552348 221536
rect 554228 221484 554280 221536
rect 554412 221552 554464 221604
rect 630864 221552 630916 221604
rect 629944 221484 629996 221536
rect 532976 221416 533028 221468
rect 533988 221416 534040 221468
rect 628932 221416 628984 221468
rect 239404 221280 239456 221332
rect 240048 221280 240100 221332
rect 241980 221280 242032 221332
rect 242808 221280 242860 221332
rect 250352 221280 250404 221332
rect 250996 221280 251048 221332
rect 252928 221280 252980 221332
rect 258080 221280 258132 221332
rect 258816 221280 258868 221332
rect 259368 221280 259420 221332
rect 268844 221280 268896 221332
rect 281724 221280 281776 221332
rect 286508 221280 286560 221332
rect 290372 221280 290424 221332
rect 292396 221280 292448 221332
rect 293224 221280 293276 221332
rect 295800 221280 295852 221332
rect 297640 221280 297692 221332
rect 298284 221280 298336 221332
rect 300216 221280 300268 221332
rect 300860 221280 300912 221332
rect 301872 221280 301924 221332
rect 303712 221280 303764 221332
rect 305276 221280 305328 221332
rect 306748 221280 306800 221332
rect 308588 221280 308640 221332
rect 309416 221280 309468 221332
rect 310244 221280 310296 221332
rect 315304 221280 315356 221332
rect 316132 221280 316184 221332
rect 317604 221280 317656 221332
rect 317972 221280 318024 221332
rect 84660 221212 84712 221264
rect 95148 221212 95200 221264
rect 187240 221212 187292 221264
rect 226616 221212 226668 221264
rect 226708 221212 226760 221264
rect 233240 221212 233292 221264
rect 238576 221212 238628 221264
rect 239956 221212 240008 221264
rect 247868 221212 247920 221264
rect 255228 221212 255280 221264
rect 256240 221212 256292 221264
rect 260840 221212 260892 221264
rect 285680 221212 285732 221264
rect 290464 221212 290516 221264
rect 316960 221212 317012 221264
rect 59176 221144 59228 221196
rect 193680 221144 193732 221196
rect 200764 221144 200816 221196
rect 246948 221144 247000 221196
rect 252008 221144 252060 221196
rect 253756 221144 253808 221196
rect 259368 221144 259420 221196
rect 260748 221144 260800 221196
rect 263784 221144 263836 221196
rect 264704 221144 264756 221196
rect 269672 221144 269724 221196
rect 270408 221144 270460 221196
rect 283932 221144 283984 221196
rect 287888 221144 287940 221196
rect 288256 221144 288308 221196
rect 292856 221144 292908 221196
rect 314476 221144 314528 221196
rect 68652 221008 68704 221060
rect 196348 221076 196400 221128
rect 199936 221076 199988 221128
rect 208124 221076 208176 221128
rect 180524 221008 180576 221060
rect 183468 221008 183520 221060
rect 188988 221008 189040 221060
rect 208032 221008 208084 221060
rect 64512 220940 64564 220992
rect 75828 220940 75880 220992
rect 197360 220940 197412 220992
rect 198648 220940 198700 220992
rect 206652 220940 206704 220992
rect 208124 220940 208176 220992
rect 69480 220872 69532 220924
rect 73160 220872 73212 220924
rect 91376 220872 91428 220924
rect 189724 220872 189776 220924
rect 189816 220872 189868 220924
rect 226708 221076 226760 221128
rect 226800 221076 226852 221128
rect 238760 221076 238812 221128
rect 240048 221076 240100 221128
rect 241428 221076 241480 221128
rect 250996 221076 251048 221128
rect 255412 221076 255464 221128
rect 277308 221076 277360 221128
rect 284484 221076 284536 221128
rect 287336 221076 287388 221128
rect 290004 221076 290056 221128
rect 314568 221076 314620 221128
rect 336740 221144 336792 221196
rect 337108 221280 337160 221332
rect 338856 221280 338908 221332
rect 340788 221280 340840 221332
rect 340880 221212 340932 221264
rect 351092 221280 351144 221332
rect 352380 221280 352432 221332
rect 390376 221280 390428 221332
rect 494520 221280 494572 221332
rect 511908 221280 511960 221332
rect 516416 221280 516468 221332
rect 520188 221280 520240 221332
rect 521660 221280 521712 221332
rect 524420 221280 524472 221332
rect 526444 221280 526496 221332
rect 529940 221280 529992 221332
rect 531504 221280 531556 221332
rect 610808 221348 610860 221400
rect 609888 221280 609940 221332
rect 341432 221144 341484 221196
rect 359924 221212 359976 221264
rect 413928 221212 413980 221264
rect 353300 221144 353352 221196
rect 481548 221212 481600 221264
rect 487804 221212 487856 221264
rect 489828 221212 489880 221264
rect 497832 221212 497884 221264
rect 511080 221212 511132 221264
rect 512000 221212 512052 221264
rect 610348 221212 610400 221264
rect 485228 221144 485280 221196
rect 506112 221144 506164 221196
rect 609428 221144 609480 221196
rect 669688 221144 669740 221196
rect 676036 221144 676088 221196
rect 337200 221076 337252 221128
rect 338120 221076 338172 221128
rect 349804 221076 349856 221128
rect 503536 221076 503588 221128
rect 608968 221076 609020 221128
rect 208400 221008 208452 221060
rect 230204 221008 230256 221060
rect 238944 221008 238996 221060
rect 260472 221008 260524 221060
rect 261944 221008 261996 221060
rect 270408 221008 270460 221060
rect 282000 221008 282052 221060
rect 282368 221008 282420 221060
rect 208308 220872 208360 220924
rect 219256 220872 219308 220924
rect 220636 220872 220688 220924
rect 220820 220872 220872 220924
rect 229560 220872 229612 220924
rect 233148 220940 233200 220992
rect 284852 221008 284904 221060
rect 290280 221008 290332 221060
rect 306288 221008 306340 221060
rect 320364 221008 320416 221060
rect 329748 221008 329800 221060
rect 346492 221008 346544 221060
rect 399300 221008 399352 221060
rect 533988 221008 534040 221060
rect 542176 221008 542228 221060
rect 543096 221008 543148 221060
rect 554412 221008 554464 221060
rect 555056 221008 555108 221060
rect 556804 221008 556856 221060
rect 557540 221008 557592 221060
rect 559288 221008 559340 221060
rect 563152 221008 563204 221060
rect 564348 221008 564400 221060
rect 571708 221008 571760 221060
rect 572720 221008 572772 221060
rect 572812 221008 572864 221060
rect 619180 221008 619232 221060
rect 669596 221008 669648 221060
rect 675852 221008 675904 221060
rect 287796 220940 287848 220992
rect 289084 220940 289136 220992
rect 290188 220940 290240 220992
rect 291568 220940 291620 220992
rect 292764 220940 292816 220992
rect 311808 220940 311860 220992
rect 327908 220940 327960 220992
rect 343272 220940 343324 220992
rect 363236 220940 363288 220992
rect 396816 220940 396868 220992
rect 534908 220940 534960 220992
rect 552204 220940 552256 220992
rect 553676 220940 553728 220992
rect 618260 220940 618312 220992
rect 667112 220940 667164 220992
rect 675944 220940 675996 220992
rect 233424 220872 233476 220924
rect 233516 220872 233568 220924
rect 238668 220872 238720 220924
rect 255412 220872 255464 220924
rect 256608 220872 256660 220924
rect 261300 220872 261352 220924
rect 262036 220872 262088 220924
rect 266360 220872 266412 220924
rect 267464 220872 267516 220924
rect 273904 220872 273956 220924
rect 284392 220872 284444 220924
rect 392216 220872 392268 220924
rect 525064 220872 525116 220924
rect 548340 220872 548392 220924
rect 617340 220872 617392 220924
rect 133420 220804 133472 220856
rect 226892 220804 226944 220856
rect 232688 220804 232740 220856
rect 234528 220804 234580 220856
rect 243636 220804 243688 220856
rect 245568 220804 245620 220856
rect 248696 220804 248748 220856
rect 251088 220804 251140 220856
rect 257896 220804 257948 220856
rect 259276 220804 259328 220856
rect 262956 220804 263008 220856
rect 264888 220804 264940 220856
rect 265532 220804 265584 220856
rect 267648 220804 267700 220856
rect 268016 220804 268068 220856
rect 281816 220804 281868 220856
rect 490196 220804 490248 220856
rect 607128 220804 607180 220856
rect 46020 220328 46072 220380
rect 647148 220328 647200 220380
rect 48504 220260 48556 220312
rect 649908 220260 649960 220312
rect 46296 220192 46348 220244
rect 648528 220192 648580 220244
rect 48596 220124 48648 220176
rect 651288 220124 651340 220176
rect 652668 220124 652720 220176
rect 675576 220124 675628 220176
rect 676036 220124 676088 220176
rect 48688 220056 48740 220108
rect 652760 220056 652812 220108
rect 652852 220056 652904 220108
rect 674840 220056 674892 220108
rect 675944 220056 675996 220108
rect 48872 219988 48924 220040
rect 655520 219988 655572 220040
rect 48780 219920 48832 219972
rect 654140 219920 654192 219972
rect 48964 219852 49016 219904
rect 656900 219852 656952 219904
rect 46664 219784 46716 219836
rect 658280 219784 658332 219836
rect 46756 219716 46808 219768
rect 659752 219716 659804 219768
rect 46204 219648 46256 219700
rect 661132 219648 661184 219700
rect 46112 219580 46164 219632
rect 663432 219580 663484 219632
rect 45836 219512 45888 219564
rect 664352 219512 664404 219564
rect 45928 219444 45980 219496
rect 664812 219444 664864 219496
rect 45744 219376 45796 219428
rect 663892 219376 663944 219428
rect 523408 218356 523460 218408
rect 523776 218356 523828 218408
rect 612648 218356 612700 218408
rect 518992 218288 519044 218340
rect 521200 218288 521252 218340
rect 612188 218288 612240 218340
rect 673920 218288 673972 218340
rect 676036 218288 676088 218340
rect 518072 218220 518124 218272
rect 518624 218220 518676 218272
rect 611728 218220 611780 218272
rect 515496 218152 515548 218204
rect 611268 218152 611320 218204
rect 487160 218084 487212 218136
rect 606668 218084 606720 218136
rect 662788 218084 662840 218136
rect 662972 218084 663024 218136
rect 673460 218084 673512 218136
rect 675944 218084 675996 218136
rect 46940 218016 46992 218068
rect 671160 218016 671212 218068
rect 674380 218016 674432 218068
rect 676036 218016 676088 218068
rect 646964 217948 647016 218000
rect 651472 217948 651524 218000
rect 644112 217880 644164 217932
rect 651564 217880 651616 217932
rect 507860 217608 507912 217660
rect 509930 217608 509982 217660
rect 513840 217608 513892 217660
rect 514990 217608 515042 217660
rect 502708 217472 502760 217524
rect 504870 217472 504922 217524
rect 570558 217472 570610 217524
rect 635924 217472 635976 217524
rect 568304 217404 568356 217456
rect 635464 217404 635516 217456
rect 492588 217336 492640 217388
rect 500316 217336 500368 217388
rect 565728 217336 565780 217388
rect 635004 217336 635056 217388
rect 563060 217268 563112 217320
rect 634544 217268 634596 217320
rect 550640 217200 550692 217252
rect 632244 217200 632296 217252
rect 540520 217132 540572 217184
rect 630404 217132 630456 217184
rect 530308 217064 530360 217116
rect 628472 217064 628524 217116
rect 535368 216996 535420 217048
rect 629484 216996 629536 217048
rect 525432 216928 525484 216980
rect 627552 216928 627604 216980
rect 418528 216860 418580 216912
rect 639696 216860 639748 216912
rect 520372 216792 520424 216844
rect 626632 216792 626684 216844
rect 41512 216724 41564 216776
rect 59360 216724 59412 216776
rect 418436 216724 418488 216776
rect 640156 216724 640208 216776
rect 41420 216656 41472 216708
rect 59452 216656 59504 216708
rect 418068 216656 418120 216708
rect 641076 216656 641128 216708
rect 642732 216656 642784 216708
rect 651380 216656 651432 216708
rect 674012 216656 674064 216708
rect 675760 216656 675812 216708
rect 41604 216588 41656 216640
rect 59268 216588 59320 216640
rect 418160 216588 418212 216640
rect 640616 216588 640668 216640
rect 495992 216520 496044 216572
rect 497004 216452 497056 216504
rect 499304 216452 499356 216504
rect 502524 216452 502576 216504
rect 484216 216384 484268 216436
rect 486700 216384 486752 216436
rect 490104 216384 490156 216436
rect 500224 216384 500276 216436
rect 500316 216384 500368 216436
rect 505008 216520 505060 216572
rect 502708 216384 502760 216436
rect 515128 216520 515180 216572
rect 625712 216520 625764 216572
rect 510252 216452 510304 216504
rect 624792 216452 624844 216504
rect 623872 216384 623924 216436
rect 622952 216316 623004 216368
rect 622492 216248 622544 216300
rect 645584 216248 645636 216300
rect 651656 216248 651708 216300
rect 673828 216248 673880 216300
rect 676036 216248 676088 216300
rect 622032 216180 622084 216232
rect 637856 216112 637908 216164
rect 636384 216044 636436 216096
rect 638316 215976 638368 216028
rect 638776 215908 638828 215960
rect 48228 215840 48280 215892
rect 665732 215840 665784 215892
rect 673552 215840 673604 215892
rect 675944 215840 675996 215892
rect 31852 215772 31904 215824
rect 666192 215772 666244 215824
rect 31668 215704 31720 215756
rect 665272 215704 665324 215756
rect 579712 215636 579764 215688
rect 599768 215636 599820 215688
rect 674104 215432 674156 215484
rect 675852 215432 675904 215484
rect 674196 215364 674248 215416
rect 675944 215364 675996 215416
rect 675208 215296 675260 215348
rect 676036 215296 676088 215348
rect 673644 214616 673696 214668
rect 676036 214616 676088 214668
rect 41512 213868 41564 213920
rect 45560 213868 45612 213920
rect 673736 213800 673788 213852
rect 675944 213800 675996 213852
rect 41512 213664 41564 213716
rect 43444 213664 43496 213716
rect 674656 212848 674708 212900
rect 674748 212644 674800 212696
rect 582288 212576 582340 212628
rect 599952 212576 600004 212628
rect 674656 212576 674708 212628
rect 675944 212576 675996 212628
rect 580264 212508 580316 212560
rect 599860 212508 599912 212560
rect 674472 212508 674524 212560
rect 676036 212508 676088 212560
rect 651288 212440 651340 212492
rect 651380 212440 651432 212492
rect 673184 212440 673236 212492
rect 675392 212440 675444 212492
rect 581644 209856 581696 209908
rect 600044 209856 600096 209908
rect 580540 209788 580592 209840
rect 599124 209788 599176 209840
rect 674288 208360 674340 208412
rect 675576 208360 675628 208412
rect 674840 208292 674892 208344
rect 675208 208292 675260 208344
rect 582288 207068 582340 207120
rect 601148 207068 601200 207120
rect 581460 207000 581512 207052
rect 600964 207000 601016 207052
rect 675668 205980 675720 206032
rect 675760 205980 675812 206032
rect 674380 205504 674432 205556
rect 675300 205504 675352 205556
rect 674380 205368 674432 205420
rect 673920 205164 673972 205216
rect 675300 205164 675352 205216
rect 675760 204960 675812 205012
rect 582288 204280 582340 204332
rect 599952 204280 600004 204332
rect 673828 202716 673880 202768
rect 675484 202716 675536 202768
rect 673644 202580 673696 202632
rect 673828 202580 673880 202632
rect 673552 202308 673604 202360
rect 674380 202308 674432 202360
rect 674840 202036 674892 202088
rect 675392 202036 675444 202088
rect 674104 201900 674156 201952
rect 674840 201900 674892 201952
rect 581828 201560 581880 201612
rect 599032 201560 599084 201612
rect 581092 201492 581144 201544
rect 599952 201492 600004 201544
rect 674196 201492 674248 201544
rect 675392 201492 675444 201544
rect 674472 200880 674524 200932
rect 675392 200880 675444 200932
rect 33048 200200 33100 200252
rect 41880 200200 41932 200252
rect 581092 200064 581144 200116
rect 599952 200064 600004 200116
rect 32956 199996 33008 200048
rect 42524 199996 42576 200048
rect 582288 198704 582340 198756
rect 599124 198704 599176 198756
rect 673644 198364 673696 198416
rect 675392 198364 675444 198416
rect 673736 197548 673788 197600
rect 675484 197548 675536 197600
rect 41880 197412 41932 197464
rect 580816 197344 580868 197396
rect 599308 197344 599360 197396
rect 581276 197276 581328 197328
rect 599952 197276 600004 197328
rect 41880 197140 41932 197192
rect 673828 197004 673880 197056
rect 675392 197004 675444 197056
rect 674656 196528 674708 196580
rect 675392 196528 675444 196580
rect 674472 196392 674524 196444
rect 674656 196392 674708 196444
rect 674840 195304 674892 195356
rect 675392 195304 675444 195356
rect 42156 195236 42208 195288
rect 42524 195236 42576 195288
rect 674380 195168 674432 195220
rect 674840 195168 674892 195220
rect 582196 194624 582248 194676
rect 599124 194624 599176 194676
rect 582288 194556 582340 194608
rect 599952 194556 600004 194608
rect 42064 193468 42116 193520
rect 42892 193468 42944 193520
rect 673460 193468 673512 193520
rect 675392 193468 675444 193520
rect 42156 192176 42208 192228
rect 42800 192176 42852 192228
rect 582288 191836 582340 191888
rect 599860 191836 599912 191888
rect 581276 191768 581328 191820
rect 599952 191768 600004 191820
rect 673552 191632 673604 191684
rect 675392 191632 675444 191684
rect 42064 191428 42116 191480
rect 43076 191428 43128 191480
rect 42156 190952 42208 191004
rect 42984 190952 43036 191004
rect 579712 190408 579764 190460
rect 599860 190408 599912 190460
rect 582196 187620 582248 187672
rect 601608 187620 601660 187672
rect 582288 187552 582340 187604
rect 600964 187552 601016 187604
rect 580264 184832 580316 184884
rect 599952 184832 600004 184884
rect 580908 184764 580960 184816
rect 601516 184764 601568 184816
rect 666744 183880 666796 183932
rect 667112 183880 667164 183932
rect 581828 182112 581880 182164
rect 599860 182112 599912 182164
rect 580540 182044 580592 182096
rect 600044 182044 600096 182096
rect 708512 179460 708564 179512
rect 704464 179392 704516 179444
rect 708420 179392 708472 179444
rect 580724 179324 580776 179376
rect 599952 179324 600004 179376
rect 666928 179324 666980 179376
rect 671436 179324 671488 179376
rect 674748 179324 674800 179376
rect 675852 179324 675904 179376
rect 704372 179324 704424 179376
rect 581092 179256 581144 179308
rect 599768 179256 599820 179308
rect 705292 179188 705344 179240
rect 707500 179324 707552 179376
rect 707040 179256 707092 179308
rect 705752 179188 705804 179240
rect 706212 179188 706264 179240
rect 706672 179188 706724 179240
rect 706304 179120 706356 179172
rect 706580 179120 706632 179172
rect 705844 179052 705896 179104
rect 707040 179052 707092 179104
rect 705384 178984 705436 179036
rect 707500 178984 707552 179036
rect 708052 178984 708104 179036
rect 704924 178916 704976 178968
rect 707960 178916 708012 178968
rect 704832 178848 704884 178900
rect 704004 178780 704056 178832
rect 708880 178780 708932 178832
rect 669412 177080 669464 177132
rect 675944 177080 675996 177132
rect 669136 176944 669188 176996
rect 676036 176944 676088 176996
rect 671436 176876 671488 176928
rect 673276 176876 673328 176928
rect 675944 176876 675996 176928
rect 667020 176808 667072 176860
rect 675760 176808 675812 176860
rect 581092 176672 581144 176724
rect 598940 176672 598992 176724
rect 581460 176604 581512 176656
rect 599860 176604 599912 176656
rect 666836 176604 666888 176656
rect 671896 176604 671948 176656
rect 674840 176604 674892 176656
rect 676036 176604 676088 176656
rect 667112 176536 667164 176588
rect 672172 176536 672224 176588
rect 674564 176332 674616 176384
rect 676036 176332 676088 176384
rect 673368 175992 673420 176044
rect 675944 175992 675996 176044
rect 674656 175516 674708 175568
rect 676036 175516 676088 175568
rect 671896 175244 671948 175296
rect 672264 175244 672316 175296
rect 675944 175244 675996 175296
rect 671896 174428 671948 174480
rect 672172 174428 672224 174480
rect 676036 174428 676088 174480
rect 580816 173884 580868 173936
rect 599952 173884 600004 173936
rect 674104 173884 674156 173936
rect 676036 173884 676088 173936
rect 579712 173816 579764 173868
rect 600044 173816 600096 173868
rect 582288 173748 582340 173800
rect 600136 173748 600188 173800
rect 674840 171640 674892 171692
rect 676036 171640 676088 171692
rect 673460 171300 673512 171352
rect 675944 171300 675996 171352
rect 582196 171164 582248 171216
rect 599952 171164 600004 171216
rect 674564 171164 674616 171216
rect 675944 171164 675996 171216
rect 579896 171096 579948 171148
rect 599860 171096 599912 171148
rect 580908 171028 580960 171080
rect 599676 171028 599728 171080
rect 676036 171096 676088 171148
rect 580080 170960 580132 171012
rect 599768 170960 599820 171012
rect 675208 170960 675260 171012
rect 673552 170008 673604 170060
rect 675944 170008 675996 170060
rect 674656 169600 674708 169652
rect 676036 169600 676088 169652
rect 673736 169192 673788 169244
rect 675944 169192 675996 169244
rect 674012 168716 674064 168768
rect 675944 168716 675996 168768
rect 674748 168648 674800 168700
rect 676036 168648 676088 168700
rect 579712 168512 579764 168564
rect 598940 168512 598992 168564
rect 673644 168512 673696 168564
rect 675852 168512 675904 168564
rect 581920 168444 581972 168496
rect 599952 168444 600004 168496
rect 580264 168376 580316 168428
rect 599492 168376 599544 168428
rect 580172 168308 580224 168360
rect 600228 168308 600280 168360
rect 672356 168240 672408 168292
rect 676036 168240 676088 168292
rect 672172 167832 672224 167884
rect 676036 167832 676088 167884
rect 672080 167424 672132 167476
rect 676036 167424 676088 167476
rect 582288 165724 582340 165776
rect 599860 165724 599912 165776
rect 580080 165656 580132 165708
rect 600044 165656 600096 165708
rect 581552 165588 581604 165640
rect 599952 165588 600004 165640
rect 581828 165520 581880 165572
rect 601424 165520 601476 165572
rect 581644 162936 581696 162988
rect 599860 162936 599912 162988
rect 581092 162868 581144 162920
rect 599952 162868 600004 162920
rect 675760 160964 675812 161016
rect 675760 160760 675812 160812
rect 582012 160216 582064 160268
rect 599952 160216 600004 160268
rect 581736 160148 581788 160200
rect 600044 160148 600096 160200
rect 581184 160080 581236 160132
rect 599860 160080 599912 160132
rect 675208 160012 675260 160064
rect 675392 160012 675444 160064
rect 674104 159332 674156 159384
rect 675484 159332 675536 159384
rect 674840 157700 674892 157752
rect 675484 157700 675536 157752
rect 580908 157496 580960 157548
rect 599952 157496 600004 157548
rect 581000 157428 581052 157480
rect 600044 157428 600096 157480
rect 580724 157360 580776 157412
rect 599860 157360 599912 157412
rect 674564 156884 674616 156936
rect 675392 156884 675444 156936
rect 674656 156476 674708 156528
rect 675392 156476 675444 156528
rect 674748 155864 674800 155916
rect 675484 155864 675536 155916
rect 582104 154640 582156 154692
rect 599952 154640 600004 154692
rect 580632 154572 580684 154624
rect 599860 154572 599912 154624
rect 673460 153348 673512 153400
rect 675392 153348 675444 153400
rect 674012 152736 674064 152788
rect 675392 152736 675444 152788
rect 673736 151988 673788 152040
rect 675392 151988 675444 152040
rect 582196 151920 582248 151972
rect 599860 151920 599912 151972
rect 581920 151852 581972 151904
rect 599952 151852 600004 151904
rect 580816 151784 580868 151836
rect 600044 151784 600096 151836
rect 673644 151376 673696 151428
rect 675392 151376 675444 151428
rect 673552 150356 673604 150408
rect 675392 150356 675444 150408
rect 581828 149200 581880 149252
rect 598940 149200 598992 149252
rect 581460 149132 581512 149184
rect 599860 149132 599912 149184
rect 581644 149064 581696 149116
rect 599952 149064 600004 149116
rect 582288 146344 582340 146396
rect 599860 146344 599912 146396
rect 581276 146276 581328 146328
rect 599952 146276 600004 146328
rect 581736 143692 581788 143744
rect 599952 143692 600004 143744
rect 579712 143624 579764 143676
rect 599584 143624 599636 143676
rect 579804 143556 579856 143608
rect 599676 143556 599728 143608
rect 581552 140904 581604 140956
rect 599860 140904 599912 140956
rect 581368 140836 581420 140888
rect 599952 140836 600004 140888
rect 581184 140768 581236 140820
rect 599308 140768 599360 140820
rect 581092 138116 581144 138168
rect 599952 138116 600004 138168
rect 581000 138048 581052 138100
rect 599860 138048 599912 138100
rect 579896 137980 579948 138032
rect 600044 137980 600096 138032
rect 580080 135328 580132 135380
rect 599860 135328 599912 135380
rect 580172 135260 580224 135312
rect 599952 135260 600004 135312
rect 704372 134308 704424 134360
rect 704464 134240 704516 134292
rect 708420 134240 708472 134292
rect 707500 134172 707552 134224
rect 708512 134172 708564 134224
rect 707040 134104 707092 134156
rect 705292 134036 705344 134088
rect 705752 134036 705804 134088
rect 706212 134036 706264 134088
rect 706580 134036 706632 134088
rect 705844 133968 705896 134020
rect 707040 133968 707092 134020
rect 706304 133900 706356 133952
rect 706580 133900 706632 133952
rect 704832 133832 704884 133884
rect 705384 133832 705436 133884
rect 707500 133832 707552 133884
rect 704924 133764 704976 133816
rect 707960 133764 708012 133816
rect 708052 133696 708104 133748
rect 704004 133628 704056 133680
rect 708880 133628 708932 133680
rect 670056 132880 670108 132932
rect 676220 132880 676272 132932
rect 669504 132744 669556 132796
rect 676128 132744 676180 132796
rect 580908 132608 580960 132660
rect 599308 132608 599360 132660
rect 669320 132608 669372 132660
rect 676036 132608 676088 132660
rect 580264 132540 580316 132592
rect 599952 132540 600004 132592
rect 579988 132472 580040 132524
rect 599860 132472 599912 132524
rect 673276 132268 673328 132320
rect 676220 132268 676272 132320
rect 670792 131656 670844 131708
rect 676036 131656 676088 131708
rect 673368 131452 673420 131504
rect 676220 131452 676272 131504
rect 672448 130840 672500 130892
rect 676036 130840 676088 130892
rect 672264 130636 672316 130688
rect 676220 130636 676272 130688
rect 670884 130024 670936 130076
rect 676036 130024 676088 130076
rect 580540 129888 580592 129940
rect 599860 129888 599912 129940
rect 580356 129820 580408 129872
rect 599952 129820 600004 129872
rect 669228 129820 669280 129872
rect 670792 129820 670844 129872
rect 580448 129752 580500 129804
rect 598940 129752 598992 129804
rect 666744 129752 666796 129804
rect 670884 129752 670936 129804
rect 671896 129684 671948 129736
rect 676036 129684 676088 129736
rect 671988 129412 672040 129464
rect 676220 129412 676272 129464
rect 674472 127712 674524 127764
rect 676036 127712 676088 127764
rect 582196 127032 582248 127084
rect 599952 127032 600004 127084
rect 673644 127032 673696 127084
rect 675944 127032 675996 127084
rect 580724 126964 580776 127016
rect 599860 126964 599912 127016
rect 674564 126964 674616 127016
rect 676036 126964 676088 127016
rect 673460 124856 673512 124908
rect 675852 124856 675904 124908
rect 674748 124448 674800 124500
rect 675944 124448 675996 124500
rect 673552 124380 673604 124432
rect 675852 124380 675904 124432
rect 582012 124312 582064 124364
rect 599952 124312 600004 124364
rect 674656 124312 674708 124364
rect 676128 124312 676180 124364
rect 580816 124244 580868 124296
rect 600044 124244 600096 124296
rect 675116 124244 675168 124296
rect 675944 124244 675996 124296
rect 580632 124176 580684 124228
rect 599860 124176 599912 124228
rect 675208 124176 675260 124228
rect 676036 124176 676088 124228
rect 673828 123224 673880 123276
rect 676036 123224 676088 123276
rect 671436 123088 671488 123140
rect 676036 123088 676088 123140
rect 672908 122680 672960 122732
rect 676036 122680 676088 122732
rect 672264 122272 672316 122324
rect 676036 122272 676088 122324
rect 582288 121592 582340 121644
rect 598940 121592 598992 121644
rect 582104 121524 582156 121576
rect 599860 121524 599912 121576
rect 581920 121456 581972 121508
rect 599952 121456 600004 121508
rect 673736 121456 673788 121508
rect 675944 121456 675996 121508
rect 583668 118804 583720 118856
rect 599860 118804 599912 118856
rect 581644 118736 581696 118788
rect 599952 118736 600004 118788
rect 581828 118668 581880 118720
rect 600044 118668 600096 118720
rect 581736 116016 581788 116068
rect 599860 116016 599912 116068
rect 581276 115948 581328 116000
rect 599952 115948 600004 116000
rect 675760 115744 675812 115796
rect 675760 115540 675812 115592
rect 675208 114996 675260 115048
rect 675392 114996 675444 115048
rect 674472 114180 674524 114232
rect 675392 114180 675444 114232
rect 581368 113228 581420 113280
rect 599952 113228 600004 113280
rect 581552 113160 581604 113212
rect 599860 113160 599912 113212
rect 674564 112344 674616 112396
rect 675392 112344 675444 112396
rect 674748 111868 674800 111920
rect 675392 111868 675444 111920
rect 674656 111120 674708 111172
rect 675392 111120 675444 111172
rect 675116 110644 675168 110696
rect 675392 110644 675444 110696
rect 581460 110508 581512 110560
rect 599952 110508 600004 110560
rect 581184 110440 581236 110492
rect 599768 110440 599820 110492
rect 673644 108196 673696 108248
rect 675484 108196 675536 108248
rect 581000 107652 581052 107704
rect 599952 107652 600004 107704
rect 673828 107516 673880 107568
rect 675392 107516 675444 107568
rect 673552 106972 673604 107024
rect 675392 106972 675444 107024
rect 673736 106360 673788 106412
rect 675392 106360 675444 106412
rect 673460 105136 673512 105188
rect 675484 105136 675536 105188
rect 581092 104864 581144 104916
rect 599952 104864 600004 104916
rect 657728 99764 657780 99816
rect 660902 99764 660954 99816
rect 580908 99356 580960 99408
rect 599952 99356 600004 99408
rect 633072 96568 633124 96620
rect 635280 96568 635332 96620
rect 636292 96568 636344 96620
rect 640984 96568 641036 96620
rect 655980 96568 656032 96620
rect 659568 96568 659620 96620
rect 661868 96568 661920 96620
rect 663064 96568 663116 96620
rect 633808 96500 633860 96552
rect 636384 96500 636436 96552
rect 637028 96500 637080 96552
rect 642364 96500 642416 96552
rect 654692 96500 654744 96552
rect 658280 96500 658332 96552
rect 659108 96500 659160 96552
rect 662512 96500 662564 96552
rect 634452 96432 634504 96484
rect 637580 96432 637632 96484
rect 652024 96432 652076 96484
rect 661960 96432 662012 96484
rect 635740 96364 635792 96416
rect 639880 96364 639932 96416
rect 631140 96024 631192 96076
rect 632106 96024 632158 96076
rect 632428 96024 632480 96076
rect 634406 96024 634458 96076
rect 635096 96024 635148 96076
rect 639006 96024 639058 96076
rect 647516 96024 647568 96076
rect 653220 96024 653272 96076
rect 631784 95888 631836 95940
rect 632980 95888 633032 95940
rect 640064 95888 640116 95940
rect 646044 95888 646096 95940
rect 638868 95820 638920 95872
rect 646228 95820 646280 95872
rect 616788 95752 616840 95804
rect 623228 95752 623280 95804
rect 639604 95752 639656 95804
rect 645952 95752 646004 95804
rect 621204 95684 621256 95736
rect 622032 95684 622084 95736
rect 637488 95684 637540 95736
rect 640524 95684 640576 95736
rect 640892 95684 640944 95736
rect 645860 95684 645912 95736
rect 603540 95616 603592 95668
rect 610440 95616 610492 95668
rect 619364 95616 619416 95668
rect 623412 95616 623464 95668
rect 641628 95616 641680 95668
rect 642824 95616 642876 95668
rect 604460 95548 604512 95600
rect 606392 95548 606444 95600
rect 607496 95548 607548 95600
rect 608968 95548 609020 95600
rect 610256 95548 610308 95600
rect 611544 95548 611596 95600
rect 612832 95548 612884 95600
rect 613568 95548 613620 95600
rect 618260 95548 618312 95600
rect 620100 95548 620152 95600
rect 621480 95548 621532 95600
rect 623320 95548 623372 95600
rect 623780 95548 623832 95600
rect 624608 95548 624660 95600
rect 638316 95548 638368 95600
rect 642272 95548 642324 95600
rect 642916 95548 642968 95600
rect 656992 95548 657044 95600
rect 659200 95548 659252 95600
rect 610164 95480 610216 95532
rect 612188 95480 612240 95532
rect 617432 95480 617484 95532
rect 623136 95480 623188 95532
rect 642732 95480 642784 95532
rect 660580 95480 660632 95532
rect 661408 95480 661460 95532
rect 620008 95412 620060 95464
rect 622308 95412 622360 95464
rect 616144 95344 616196 95396
rect 622492 95344 622544 95396
rect 656624 95344 656676 95396
rect 663156 95344 663208 95396
rect 646780 95276 646832 95328
rect 663340 95276 663392 95328
rect 589188 95208 589240 95260
rect 610900 95208 610952 95260
rect 643560 95208 643612 95260
rect 644848 95208 644900 95260
rect 651472 95208 651524 95260
rect 653404 95208 653456 95260
rect 657084 95208 657136 95260
rect 657912 95208 657964 95260
rect 646136 95140 646188 95192
rect 663432 95140 663484 95192
rect 597468 95072 597520 95124
rect 607680 95072 607732 95124
rect 646688 95072 646740 95124
rect 648160 95072 648212 95124
rect 648896 95072 648948 95124
rect 650736 95072 650788 95124
rect 652668 95072 652720 95124
rect 663800 95072 663852 95124
rect 614856 94936 614908 94988
rect 615408 94936 615460 94988
rect 648712 94800 648764 94852
rect 650092 94800 650144 94852
rect 618720 94732 618772 94784
rect 623320 94732 623372 94784
rect 645952 94732 646004 94784
rect 646228 94732 646280 94784
rect 648804 94664 648856 94716
rect 649448 94664 649500 94716
rect 653312 94664 653364 94716
rect 663708 94664 663760 94716
rect 657268 94596 657320 94648
rect 663524 94596 663576 94648
rect 618076 94528 618128 94580
rect 621940 94528 621992 94580
rect 656900 94528 656952 94580
rect 658556 94528 658608 94580
rect 648068 94460 648120 94512
rect 659844 94460 659896 94512
rect 660396 94460 660448 94512
rect 643468 94188 643520 94240
rect 644204 94052 644256 94104
rect 654048 94052 654100 94104
rect 649356 93984 649408 94036
rect 656900 93984 656952 94036
rect 644756 93848 644808 93900
rect 653496 93848 653548 93900
rect 613016 91672 613068 91724
rect 614948 91672 615000 91724
rect 590660 89632 590712 89684
rect 603540 89632 603592 89684
rect 657084 88816 657136 88868
rect 658004 88816 658056 88868
rect 659476 88816 659528 88868
rect 663616 88816 663668 88868
rect 578148 85552 578200 85604
rect 589188 85552 589240 85604
rect 648896 85484 648948 85536
rect 657176 85484 657228 85536
rect 651472 85416 651524 85468
rect 658832 85416 658884 85468
rect 648804 85348 648856 85400
rect 660672 85348 660724 85400
rect 648712 85280 648764 85332
rect 657728 85280 657780 85332
rect 643560 85212 643612 85264
rect 660120 85212 660172 85264
rect 646688 85144 646740 85196
rect 661408 85144 661460 85196
rect 586428 84600 586480 84652
rect 600320 84600 600372 84652
rect 583852 84532 583904 84584
rect 600504 84532 600556 84584
rect 583760 84464 583812 84516
rect 600688 84464 600740 84516
rect 582288 84396 582340 84448
rect 600228 84396 600280 84448
rect 582012 84328 582064 84380
rect 600412 84328 600464 84380
rect 582196 84260 582248 84312
rect 600596 84260 600648 84312
rect 582104 84192 582156 84244
rect 600780 84192 600832 84244
rect 581920 84124 581972 84176
rect 600872 84124 600924 84176
rect 607220 83784 607272 83836
rect 612924 83784 612976 83836
rect 598940 82764 598992 82816
rect 610164 82900 610216 82952
rect 605748 82832 605800 82884
rect 610348 82832 610400 82884
rect 579620 82628 579672 82680
rect 583668 82628 583720 82680
rect 580816 81472 580868 81524
rect 581092 81472 581144 81524
rect 578240 75760 578292 75812
rect 590660 75760 590712 75812
rect 600320 75352 600372 75404
rect 607220 75352 607272 75404
rect 581000 72156 581052 72208
rect 598848 72156 598900 72208
rect 629300 71952 629352 72004
rect 631508 71952 631560 72004
rect 602620 71748 602672 71800
rect 612832 71748 612884 71800
rect 578332 69028 578384 69080
rect 581000 69028 581052 69080
rect 594708 66240 594760 66292
rect 600320 66240 600372 66292
rect 587900 66172 587952 66224
rect 597468 66172 597520 66224
rect 580724 65968 580776 66020
rect 586428 65968 586480 66020
rect 594340 63724 594392 63776
rect 605748 63724 605800 63776
rect 597560 63520 597612 63572
rect 602620 63520 602672 63572
rect 579620 59848 579672 59900
rect 583760 59848 583812 59900
rect 579804 59032 579856 59084
rect 594340 59032 594392 59084
rect 579620 58624 579672 58676
rect 583852 58624 583904 58676
rect 599124 55496 599176 55548
rect 604460 55496 604512 55548
rect 576768 55156 576820 55208
rect 579804 55224 579856 55276
rect 587900 53660 587952 53712
rect 571340 53592 571392 53644
rect 346860 52368 346912 52420
rect 642916 52368 642968 52420
rect 230388 51416 230440 51468
rect 642824 51416 642876 51468
rect 212448 51348 212500 51400
rect 639328 51348 639380 51400
rect 559472 51008 559524 51060
rect 578240 51008 578292 51060
rect 565820 49648 565872 49700
rect 578332 49716 578384 49768
rect 590660 49716 590712 49768
rect 597560 49716 597612 49768
rect 478144 48492 478196 48544
rect 526168 48492 526220 48544
rect 215208 48424 215260 48476
rect 346492 48424 346544 48476
rect 412640 48424 412692 48476
rect 494060 48424 494112 48476
rect 149980 48356 150032 48408
rect 150256 48356 150308 48408
rect 218060 48356 218112 48408
rect 281448 48356 281500 48408
rect 506388 48356 506440 48408
rect 216128 48288 216180 48340
rect 518532 48288 518584 48340
rect 590752 48288 590804 48340
rect 599124 48288 599176 48340
rect 535460 47200 535512 47252
rect 543004 47200 543056 47252
rect 52092 47064 52144 47116
rect 213828 47064 213880 47116
rect 215208 47064 215260 47116
rect 52276 46996 52328 47048
rect 149980 46996 150032 47048
rect 494060 46860 494112 46912
rect 502248 46860 502300 46912
rect 646320 46860 646372 46912
rect 666560 46860 666612 46912
rect 460664 45772 460716 45824
rect 610256 45772 610308 45824
rect 367100 45704 367152 45756
rect 607312 45704 607364 45756
rect 312820 45636 312872 45688
rect 607588 45636 607640 45688
rect 230848 45568 230900 45620
rect 613016 45568 613068 45620
rect 85120 45500 85172 45552
rect 475660 45500 475712 45552
rect 524052 45500 524104 45552
rect 559472 45500 559524 45552
rect 312820 44140 312872 44192
rect 367100 44140 367152 44192
rect 565820 44140 565872 44192
rect 571340 44140 571392 44192
rect 310428 44072 310480 44124
rect 365168 44072 365220 44124
rect 444564 44072 444616 44124
rect 576768 44140 576820 44192
rect 474464 44004 474516 44056
rect 590660 44140 590712 44192
rect 419724 43936 419776 43988
rect 578148 43936 578200 43988
rect 405556 43868 405608 43920
rect 607496 43868 607548 43920
rect 230572 43800 230624 43852
rect 618260 43800 618312 43852
rect 231032 43732 231084 43784
rect 621480 43732 621532 43784
rect 230940 43664 230992 43716
rect 621204 43664 621256 43716
rect 230756 43596 230808 43648
rect 621572 43596 621624 43648
rect 230664 43528 230716 43580
rect 621296 43528 621348 43580
rect 230480 43460 230532 43512
rect 621388 43460 621440 43512
rect 226248 43392 226300 43444
rect 622492 43392 622544 43444
rect 223488 43324 223540 43376
rect 622308 43324 622360 43376
rect 209688 43256 209740 43308
rect 629300 43256 629352 43308
rect 615408 42916 615460 42968
rect 641168 42916 641220 42968
rect 52184 42848 52236 42900
rect 215300 42848 215352 42900
rect 507860 42236 507912 42288
rect 530676 42236 530728 42288
rect 531044 42236 531096 42288
rect 565728 42236 565780 42288
rect 506388 41896 506440 41948
rect 520372 41896 520424 41948
rect 502248 41828 502300 41880
rect 518532 41828 518584 41880
rect 416688 41760 416740 41812
rect 420736 41760 420788 41812
rect 471704 41760 471756 41812
rect 475568 41760 475620 41812
rect 514024 41760 514076 41812
rect 514852 41760 514904 41812
rect 141792 41488 141844 41540
rect 207020 41488 207072 41540
rect 209688 41488 209740 41540
rect 420736 38564 420788 38616
rect 444564 38632 444616 38684
rect 475568 38564 475620 38616
rect 507860 38564 507912 38616
rect 475660 38496 475712 38548
rect 514024 38496 514076 38548
rect 213184 24760 213236 24812
rect 213828 24760 213880 24812
rect 224592 22992 224644 23044
rect 226248 22992 226300 23044
rect 221740 22516 221792 22568
rect 223488 22516 223540 22568
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366284 1027806 366496 1027834
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366284 1027752 366312 1027806
rect 366468 1027752 366496 1027806
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366284 1024434 366312 1024488
rect 366468 1024434 366496 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366284 1024406 366496 1024434
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 425978 1006088 426034 1006097
rect 425978 1006023 425980 1006032
rect 426032 1006023 426034 1006032
rect 458916 1006052 458968 1006058
rect 425980 1005994 426032 1006000
rect 458916 1005994 458968 1006000
rect 424322 1005952 424378 1005961
rect 424322 1005887 424324 1005896
rect 424376 1005887 424378 1005896
rect 440424 1005916 440476 1005922
rect 424324 1005858 424376 1005864
rect 440424 1005858 440476 1005864
rect 423864 1005848 423916 1005854
rect 423862 1005816 423864 1005825
rect 440240 1005848 440292 1005854
rect 423916 1005816 423918 1005825
rect 440240 1005790 440292 1005796
rect 423862 1005751 423918 1005760
rect 356058 1005680 356114 1005689
rect 356058 1005615 356060 1005624
rect 356112 1005615 356114 1005624
rect 373172 1005644 373224 1005650
rect 356060 1005586 356112 1005592
rect 373172 1005586 373224 1005592
rect 356888 1005576 356940 1005582
rect 356886 1005544 356888 1005553
rect 356940 1005544 356942 1005553
rect 356886 1005479 356942 1005488
rect 144828 1005440 144880 1005446
rect 160284 1005440 160336 1005446
rect 144828 1005382 144880 1005388
rect 160282 1005408 160284 1005417
rect 356520 1005440 356572 1005446
rect 160336 1005408 160338 1005417
rect 92664 1005304 92716 1005310
rect 109316 1005304 109368 1005310
rect 92664 1005246 92716 1005252
rect 106462 1005272 106518 1005281
rect 92572 999932 92624 999938
rect 92572 999874 92624 999880
rect 92480 999864 92532 999870
rect 92480 999806 92532 999812
rect 92296 999796 92348 999802
rect 92296 999738 92348 999744
rect 86040 995852 86092 995858
rect 86040 995794 86092 995800
rect 86052 995738 86080 995794
rect 92308 995790 92336 999738
rect 92388 999660 92440 999666
rect 92388 999602 92440 999608
rect 91560 995784 91612 995790
rect 86590 995752 86646 995761
rect 85698 995710 86080 995738
rect 86342 995710 86590 995738
rect 89378 995722 89760 995738
rect 91218 995732 91560 995738
rect 91218 995726 91612 995732
rect 92296 995784 92348 995790
rect 92296 995726 92348 995732
rect 89378 995716 89772 995722
rect 89378 995710 89720 995716
rect 86590 995687 86646 995696
rect 91218 995710 91600 995726
rect 89720 995658 89772 995664
rect 92400 995654 92428 999602
rect 92492 995722 92520 999806
rect 92480 995716 92532 995722
rect 92480 995658 92532 995664
rect 77944 995648 77996 995654
rect 77694 995596 77944 995602
rect 92388 995648 92440 995654
rect 87786 995616 87842 995625
rect 77694 995590 77996 995596
rect 77694 995574 77984 995590
rect 87538 995574 87786 995602
rect 88734 995586 89024 995602
rect 92388 995590 92440 995596
rect 92584 995586 92612 999874
rect 88734 995580 89036 995586
rect 88734 995574 88984 995580
rect 87786 995551 87842 995560
rect 88984 995522 89036 995528
rect 92572 995580 92624 995586
rect 92572 995522 92624 995528
rect 81622 995480 81678 995489
rect 77036 993682 77064 995452
rect 78324 993721 78352 995452
rect 80164 993857 80192 995452
rect 80716 995217 80744 995452
rect 81374 995438 81622 995466
rect 85302 995480 85358 995489
rect 81622 995415 81678 995424
rect 82004 995353 82032 995452
rect 81990 995344 82046 995353
rect 81990 995279 82046 995288
rect 84488 995217 84516 995452
rect 85054 995438 85302 995466
rect 85302 995415 85358 995424
rect 80702 995208 80758 995217
rect 80702 995143 80758 995152
rect 84474 995208 84530 995217
rect 84474 995143 84530 995152
rect 80150 993848 80206 993857
rect 80150 993783 80206 993792
rect 78310 993712 78366 993721
rect 77024 993676 77076 993682
rect 78310 993647 78366 993656
rect 77024 993618 77076 993624
rect 92676 990854 92704 1005246
rect 106462 1005207 106464 1005216
rect 106516 1005207 106518 1005216
rect 109314 1005272 109316 1005281
rect 109368 1005272 109370 1005281
rect 109314 1005207 109370 1005216
rect 125784 1005236 125836 1005242
rect 106464 1005178 106516 1005184
rect 125784 1005178 125836 1005184
rect 105636 1005168 105688 1005174
rect 105634 1005136 105636 1005145
rect 125600 1005168 125652 1005174
rect 105688 1005136 105690 1005145
rect 125600 1005110 125652 1005116
rect 105634 1005071 105690 1005080
rect 108028 1004896 108080 1004902
rect 108026 1004864 108028 1004873
rect 109684 1004896 109736 1004902
rect 108080 1004864 108082 1004873
rect 108026 1004799 108082 1004808
rect 109682 1004864 109684 1004873
rect 109736 1004864 109738 1004873
rect 109682 1004799 109738 1004808
rect 114650 1004864 114706 1004873
rect 114650 1004799 114652 1004808
rect 114704 1004799 114706 1004808
rect 114652 1004770 114704 1004776
rect 99472 1004760 99524 1004766
rect 98274 1004728 98330 1004737
rect 92940 1004692 92992 1004698
rect 98642 1004728 98698 1004737
rect 98330 1004686 98642 1004714
rect 98274 1004663 98330 1004672
rect 98642 1004663 98698 1004672
rect 99470 1004728 99472 1004737
rect 99524 1004728 99526 1004737
rect 99470 1004663 99526 1004672
rect 108854 1004728 108910 1004737
rect 108854 1004663 108856 1004672
rect 92940 1004634 92992 1004640
rect 108908 1004663 108910 1004672
rect 125508 1004692 125560 1004698
rect 108856 1004634 108908 1004640
rect 125508 1004634 125560 1004640
rect 92756 999524 92808 999530
rect 92756 999466 92808 999472
rect 92768 995081 92796 999466
rect 92754 995072 92810 995081
rect 92754 995007 92810 995016
rect 92492 990826 92704 990854
rect 92492 990146 92520 990826
rect 89628 990140 89680 990146
rect 89628 990082 89680 990088
rect 92480 990140 92532 990146
rect 92480 990082 92532 990088
rect 73436 989460 73488 989466
rect 73436 989402 73488 989408
rect 45468 988032 45520 988038
rect 45468 987974 45520 987980
rect 42340 972936 42392 972942
rect 42340 972878 42392 972884
rect 41800 968833 41828 969272
rect 41786 968824 41842 968833
rect 41786 968759 41842 968768
rect 42076 967094 42104 967405
rect 42352 967298 42380 972878
rect 42156 967292 42208 967298
rect 42156 967234 42208 967240
rect 42340 967292 42392 967298
rect 42340 967234 42392 967240
rect 42064 967088 42116 967094
rect 42064 967030 42116 967036
rect 42168 966756 42196 967234
rect 42800 967088 42852 967094
rect 42800 967030 42852 967036
rect 41800 965161 41828 965565
rect 41786 965152 41842 965161
rect 41786 965087 41842 965096
rect 42168 964034 42196 964376
rect 42156 964028 42208 964034
rect 42156 963970 42208 963976
rect 41800 963393 41828 963725
rect 41786 963384 41842 963393
rect 41786 963319 41842 963328
rect 42168 962674 42196 963084
rect 42156 962668 42208 962674
rect 42156 962610 42208 962616
rect 42168 962130 42196 962540
rect 42156 962124 42208 962130
rect 42156 962066 42208 962072
rect 42076 959546 42104 960024
rect 42064 959540 42116 959546
rect 42064 959482 42116 959488
rect 42168 959138 42196 959412
rect 42156 959132 42208 959138
rect 42156 959074 42208 959080
rect 42076 958390 42104 958732
rect 42064 958384 42116 958390
rect 42064 958326 42116 958332
rect 42076 957778 42104 958188
rect 42064 957772 42116 957778
rect 42064 957714 42116 957720
rect 42182 956338 42380 956366
rect 42168 955398 42196 955740
rect 42156 955392 42208 955398
rect 42156 955334 42208 955340
rect 42168 955182 42288 955210
rect 42168 955060 42196 955182
rect 35624 949612 35676 949618
rect 35624 949554 35676 949560
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 35636 934153 35664 949554
rect 35716 949544 35768 949550
rect 35716 949486 35768 949492
rect 35806 949512 35862 949521
rect 35728 934561 35756 949486
rect 35806 949447 35862 949456
rect 41512 949476 41564 949482
rect 35820 934969 35848 949447
rect 41512 949418 41564 949424
rect 41524 943945 41552 949418
rect 41510 943936 41566 943945
rect 41510 943871 41566 943880
rect 41972 943288 42024 943294
rect 41972 943230 42024 943236
rect 41786 943120 41842 943129
rect 41786 943055 41788 943064
rect 41840 943055 41842 943064
rect 41788 943026 41840 943032
rect 41788 942744 41840 942750
rect 41786 942712 41788 942721
rect 41840 942712 41842 942721
rect 41786 942647 41842 942656
rect 41878 942304 41934 942313
rect 41878 942239 41934 942248
rect 41788 941520 41840 941526
rect 41786 941488 41788 941497
rect 41840 941488 41842 941497
rect 41786 941423 41842 941432
rect 41788 941384 41840 941390
rect 41788 941326 41840 941332
rect 41694 940536 41750 940545
rect 41694 940471 41750 940480
rect 41708 936562 41736 940471
rect 41800 936601 41828 941326
rect 41892 941254 41920 942239
rect 41984 941905 42012 943230
rect 41970 941896 42026 941905
rect 41970 941831 42026 941840
rect 41880 941248 41932 941254
rect 41880 941190 41932 941196
rect 41878 941080 41934 941089
rect 41878 941015 41934 941024
rect 41786 936592 41842 936601
rect 41144 936556 41196 936562
rect 41144 936498 41196 936504
rect 41696 936556 41748 936562
rect 41786 936527 41842 936536
rect 41696 936498 41748 936504
rect 35806 934960 35862 934969
rect 35806 934895 35862 934904
rect 35714 934552 35770 934561
rect 35714 934487 35770 934496
rect 35622 934144 35678 934153
rect 35622 934079 35678 934088
rect 41156 819806 41184 936498
rect 41892 936442 41920 941015
rect 41970 940264 42026 940273
rect 41970 940199 42026 940208
rect 41984 938505 42012 940199
rect 41970 938496 42026 938505
rect 41970 938431 42026 938440
rect 42260 938233 42288 955182
rect 42352 939049 42380 956338
rect 42708 955392 42760 955398
rect 42708 955334 42760 955340
rect 42720 941390 42748 955334
rect 42708 941384 42760 941390
rect 42708 941326 42760 941332
rect 42708 941248 42760 941254
rect 42708 941190 42760 941196
rect 42338 939040 42394 939049
rect 42338 938975 42394 938984
rect 42246 938224 42302 938233
rect 42246 938159 42302 938168
rect 41708 936414 41920 936442
rect 41510 922040 41566 922049
rect 41510 921975 41566 921984
rect 41144 819800 41196 819806
rect 41144 819742 41196 819748
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 41156 814303 41184 819742
rect 41524 814450 41552 921975
rect 41708 902534 41736 936414
rect 41786 933328 41842 933337
rect 41786 933263 41842 933272
rect 41800 932521 41828 933263
rect 41786 932512 41842 932521
rect 41786 932447 41788 932456
rect 41840 932447 41842 932456
rect 41788 932418 41840 932424
rect 41800 932387 41828 932418
rect 41616 902506 41736 902534
rect 41616 844574 41644 902506
rect 41616 844546 41736 844574
rect 41708 815833 41736 844546
rect 41786 817728 41842 817737
rect 41786 817663 41842 817672
rect 41800 817494 41828 817663
rect 41788 817488 41840 817494
rect 41788 817430 41840 817436
rect 41788 817352 41840 817358
rect 41786 817320 41788 817329
rect 41840 817320 41842 817329
rect 41786 817255 41842 817264
rect 42720 817018 42748 941190
rect 42812 938641 42840 967030
rect 42984 964028 43036 964034
rect 42984 963970 43036 963976
rect 42892 962668 42944 962674
rect 42892 962610 42944 962616
rect 42904 959682 42932 962610
rect 42892 959676 42944 959682
rect 42892 959618 42944 959624
rect 42892 959540 42944 959546
rect 42892 959482 42944 959488
rect 42904 949550 42932 959482
rect 42892 949544 42944 949550
rect 42892 949486 42944 949492
rect 42996 939978 43024 963970
rect 43076 962124 43128 962130
rect 43076 962066 43128 962072
rect 42904 939950 43024 939978
rect 42798 938632 42854 938641
rect 42798 938567 42854 938576
rect 42904 933745 42932 939950
rect 42982 939856 43038 939865
rect 42982 939791 43038 939800
rect 42890 933736 42946 933745
rect 42890 933671 42946 933680
rect 42798 922040 42854 922049
rect 42798 921975 42854 921984
rect 42708 817012 42760 817018
rect 42708 816954 42760 816960
rect 41970 816504 42026 816513
rect 41970 816439 42026 816448
rect 41694 815824 41750 815833
rect 41694 815759 41750 815768
rect 41524 814422 41920 814450
rect 41142 814294 41198 814303
rect 41142 814229 41198 814238
rect 41788 814292 41840 814298
rect 41788 814234 41840 814240
rect 41800 813657 41828 814234
rect 41892 814065 41920 814422
rect 41984 814201 42012 816439
rect 42720 816105 42748 816954
rect 42706 816096 42762 816105
rect 42706 816031 42762 816040
rect 41970 814192 42026 814201
rect 41970 814127 42026 814136
rect 41878 814056 41934 814065
rect 41878 813991 41934 814000
rect 42338 814056 42394 814065
rect 42338 813991 42394 814000
rect 41786 813648 41842 813657
rect 41786 813583 41842 813592
rect 41786 811608 41842 811617
rect 41786 811543 41842 811552
rect 41800 810082 41828 811543
rect 41970 811200 42026 811209
rect 41970 811135 42026 811144
rect 41788 810076 41840 810082
rect 41788 810018 41840 810024
rect 41786 808344 41842 808353
rect 41786 808279 41842 808288
rect 41800 807634 41828 808279
rect 41878 807936 41934 807945
rect 41878 807871 41880 807880
rect 41932 807871 41934 807880
rect 41880 807842 41932 807848
rect 41788 807628 41840 807634
rect 41788 807570 41840 807576
rect 41786 807528 41842 807537
rect 41786 807463 41842 807472
rect 41800 806721 41828 807463
rect 41786 806712 41842 806721
rect 41786 806647 41788 806656
rect 41840 806647 41842 806656
rect 41788 806618 41840 806624
rect 41984 800222 42012 811135
rect 41972 800216 42024 800222
rect 41972 800158 42024 800164
rect 41972 800012 42024 800018
rect 41972 799954 42024 799960
rect 41984 799445 42012 799954
rect 42352 799746 42380 813991
rect 42614 809568 42670 809577
rect 42614 809503 42670 809512
rect 42340 799740 42392 799746
rect 42340 799682 42392 799688
rect 42156 798176 42208 798182
rect 42156 798118 42208 798124
rect 42168 797605 42196 798118
rect 42628 797858 42656 809503
rect 42708 807628 42760 807634
rect 42708 807570 42760 807576
rect 42720 797978 42748 807570
rect 42708 797972 42760 797978
rect 42708 797914 42760 797920
rect 42628 797830 42748 797858
rect 42432 797632 42484 797638
rect 42432 797574 42484 797580
rect 42156 797292 42208 797298
rect 42156 797234 42208 797240
rect 42168 796960 42196 797234
rect 42156 796340 42208 796346
rect 42156 796282 42208 796288
rect 42168 795765 42196 796282
rect 42156 795048 42208 795054
rect 42156 794990 42208 794996
rect 42168 794580 42196 794990
rect 42156 794300 42208 794306
rect 42156 794242 42208 794248
rect 42168 793900 42196 794242
rect 42444 793830 42472 797574
rect 42720 796346 42748 797830
rect 42708 796340 42760 796346
rect 42708 796282 42760 796288
rect 42156 793824 42208 793830
rect 42156 793766 42208 793772
rect 42432 793824 42484 793830
rect 42432 793766 42484 793772
rect 42168 793288 42196 793766
rect 42156 793008 42208 793014
rect 42156 792950 42208 792956
rect 42168 792744 42196 792950
rect 42156 790696 42208 790702
rect 42156 790638 42208 790644
rect 42168 790228 42196 790638
rect 42156 790152 42208 790158
rect 42156 790094 42208 790100
rect 42168 789616 42196 790094
rect 42156 789336 42208 789342
rect 42156 789278 42208 789284
rect 42168 788936 42196 789278
rect 42156 788860 42208 788866
rect 42156 788802 42208 788808
rect 42168 788392 42196 788802
rect 42156 787024 42208 787030
rect 42156 786966 42208 786972
rect 42168 786556 42196 786966
rect 42064 786276 42116 786282
rect 42064 786218 42116 786224
rect 42076 785944 42104 786218
rect 42156 785800 42208 785806
rect 42156 785742 42208 785748
rect 42168 785264 42196 785742
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 41512 774784 41564 774790
rect 41510 774752 41512 774761
rect 41564 774752 41566 774761
rect 41510 774687 41566 774696
rect 41788 774240 41840 774246
rect 41788 774182 41840 774188
rect 41800 774081 41828 774182
rect 41786 774072 41842 774081
rect 41786 774007 41842 774016
rect 41512 773968 41564 773974
rect 41510 773936 41512 773945
rect 41564 773936 41566 773945
rect 41510 773871 41566 773880
rect 41512 773628 41564 773634
rect 41512 773570 41564 773576
rect 41524 773537 41552 773570
rect 41510 773528 41566 773537
rect 41510 773463 41566 773472
rect 42154 772032 42210 772041
rect 42154 771967 42210 771976
rect 41878 767952 41934 767961
rect 41878 767887 41934 767896
rect 41510 764144 41566 764153
rect 41510 764079 41566 764088
rect 30378 763736 30434 763745
rect 30378 763671 30434 763680
rect 30392 763337 30420 763671
rect 41524 763337 41552 764079
rect 30378 763328 30434 763337
rect 30378 763263 30434 763272
rect 41510 763328 41566 763337
rect 41510 763263 41512 763272
rect 41564 763263 41566 763272
rect 41512 763234 41564 763240
rect 41892 757042 41920 767887
rect 42062 766728 42118 766737
rect 42062 766663 42118 766672
rect 41972 760572 42024 760578
rect 41972 760514 42024 760520
rect 41984 757081 42012 760514
rect 42076 757450 42104 766663
rect 42168 757518 42196 771967
rect 42430 770808 42486 770817
rect 42430 770743 42486 770752
rect 42444 757654 42472 770743
rect 42706 769992 42762 770001
rect 42706 769927 42762 769936
rect 42432 757648 42484 757654
rect 42432 757590 42484 757596
rect 42156 757512 42208 757518
rect 42156 757454 42208 757460
rect 42064 757444 42116 757450
rect 42064 757386 42116 757392
rect 42432 757444 42484 757450
rect 42432 757386 42484 757392
rect 41970 757072 42026 757081
rect 41880 757036 41932 757042
rect 41970 757007 42026 757016
rect 41880 756978 41932 756984
rect 41880 756764 41932 756770
rect 41880 756706 41932 756712
rect 41892 756228 41920 756706
rect 42444 755546 42472 757386
rect 42720 756566 42748 769927
rect 42708 756560 42760 756566
rect 42708 756502 42760 756508
rect 42432 755540 42484 755546
rect 42432 755482 42484 755488
rect 42616 755268 42668 755274
rect 42616 755210 42668 755216
rect 42156 754928 42208 754934
rect 42156 754870 42208 754876
rect 42168 754392 42196 754870
rect 42062 754080 42118 754089
rect 42062 754015 42118 754024
rect 42076 753780 42104 754015
rect 42156 753092 42208 753098
rect 42156 753034 42208 753040
rect 42168 752556 42196 753034
rect 42156 751800 42208 751806
rect 42156 751742 42208 751748
rect 42168 751369 42196 751742
rect 42156 751120 42208 751126
rect 42156 751062 42208 751068
rect 42168 750720 42196 751062
rect 42064 750644 42116 750650
rect 42064 750586 42116 750592
rect 42076 750108 42104 750586
rect 42156 749828 42208 749834
rect 42156 749770 42208 749776
rect 42168 749529 42196 749770
rect 42628 749018 42656 755210
rect 42616 749012 42668 749018
rect 42616 748954 42668 748960
rect 42168 746978 42196 747048
rect 42156 746972 42208 746978
rect 42156 746914 42208 746920
rect 42156 746768 42208 746774
rect 42156 746710 42208 746716
rect 42168 746401 42196 746710
rect 42156 746292 42208 746298
rect 42156 746234 42208 746240
rect 42168 745756 42196 746234
rect 42156 745476 42208 745482
rect 42156 745418 42208 745424
rect 42168 745212 42196 745418
rect 42156 743776 42208 743782
rect 42156 743718 42208 743724
rect 42168 743376 42196 743718
rect 42156 743300 42208 743306
rect 42156 743242 42208 743248
rect 42168 742696 42196 743242
rect 42156 742620 42208 742626
rect 42156 742562 42208 742568
rect 42168 742084 42196 742562
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 41788 731400 41840 731406
rect 41786 731368 41788 731377
rect 41840 731368 41842 731377
rect 41786 731303 41842 731312
rect 41512 731128 41564 731134
rect 39394 731096 39450 731105
rect 39394 731031 39450 731040
rect 41510 731096 41512 731105
rect 41564 731096 41566 731105
rect 41510 731031 41566 731040
rect 39408 729881 39436 731031
rect 41512 730720 41564 730726
rect 41510 730688 41512 730697
rect 41564 730688 41566 730697
rect 41510 730623 41566 730632
rect 41512 730516 41564 730522
rect 41512 730458 41564 730464
rect 39394 729872 39450 729881
rect 39394 729807 39450 729816
rect 39408 728249 39436 729807
rect 41524 729473 41552 730458
rect 42812 730153 42840 921975
rect 42996 902534 43024 939791
rect 43088 937417 43116 962066
rect 43628 959676 43680 959682
rect 43628 959618 43680 959624
rect 43352 959132 43404 959138
rect 43352 959074 43404 959080
rect 43168 958384 43220 958390
rect 43168 958326 43220 958332
rect 43074 937408 43130 937417
rect 43074 937343 43130 937352
rect 43180 936193 43208 958326
rect 43260 957772 43312 957778
rect 43260 957714 43312 957720
rect 43272 937825 43300 957714
rect 43258 937816 43314 937825
rect 43258 937751 43314 937760
rect 43166 936184 43222 936193
rect 43166 936119 43222 936128
rect 43364 935785 43392 959074
rect 43640 949618 43668 959618
rect 43628 949612 43680 949618
rect 43628 949554 43680 949560
rect 43350 935776 43406 935785
rect 43350 935711 43406 935720
rect 43994 927208 44050 927217
rect 43994 927143 44050 927152
rect 42904 902506 43024 902534
rect 42904 814298 42932 902506
rect 43534 815280 43590 815289
rect 43534 815215 43590 815224
rect 43442 814872 43498 814881
rect 43442 814807 43498 814816
rect 42892 814292 42944 814298
rect 42892 814234 42944 814240
rect 43350 813240 43406 813249
rect 43350 813175 43406 813184
rect 42890 812832 42946 812841
rect 42890 812767 42946 812776
rect 42904 798182 42932 812767
rect 42982 812424 43038 812433
rect 42982 812359 43038 812368
rect 42892 798176 42944 798182
rect 42892 798118 42944 798124
rect 42996 798028 43024 812359
rect 43074 812016 43130 812025
rect 43074 811951 43130 811960
rect 42904 798000 43024 798028
rect 42904 785806 42932 798000
rect 42984 797904 43036 797910
rect 42984 797846 43036 797852
rect 42892 785800 42944 785806
rect 42892 785742 42944 785748
rect 42996 776914 43024 797846
rect 43088 788866 43116 811951
rect 43258 809160 43314 809169
rect 43258 809095 43314 809104
rect 43168 807900 43220 807906
rect 43168 807842 43220 807848
rect 43180 795054 43208 807842
rect 43168 795048 43220 795054
rect 43168 794990 43220 794996
rect 43272 794306 43300 809095
rect 43260 794300 43312 794306
rect 43260 794242 43312 794248
rect 43076 788860 43128 788866
rect 43076 788802 43128 788808
rect 43364 787030 43392 813175
rect 43456 797978 43484 814807
rect 43444 797972 43496 797978
rect 43444 797914 43496 797920
rect 43548 797858 43576 815215
rect 43810 810792 43866 810801
rect 43810 810727 43866 810736
rect 43720 810076 43772 810082
rect 43720 810018 43772 810024
rect 43626 808752 43682 808761
rect 43626 808687 43682 808696
rect 43456 797830 43576 797858
rect 43352 787024 43404 787030
rect 43352 786966 43404 786972
rect 42904 776886 43024 776914
rect 42904 772886 42932 776886
rect 43352 773628 43404 773634
rect 43352 773570 43404 773576
rect 42892 772880 42944 772886
rect 42892 772822 42944 772828
rect 42904 771225 42932 772822
rect 42890 771216 42946 771225
rect 42890 771151 42946 771160
rect 43074 769584 43130 769593
rect 43074 769519 43130 769528
rect 42890 764688 42946 764697
rect 42890 764623 42946 764632
rect 42904 751806 42932 764623
rect 42984 757648 43036 757654
rect 42984 757590 43036 757596
rect 42892 751800 42944 751806
rect 42892 751742 42944 751748
rect 42798 730144 42854 730153
rect 42798 730079 42854 730088
rect 41510 729464 41566 729473
rect 41510 729399 41566 729408
rect 42996 729298 43024 757590
rect 43088 754934 43116 769519
rect 43166 768360 43222 768369
rect 43166 768295 43222 768304
rect 43180 766426 43208 768295
rect 43258 767544 43314 767553
rect 43258 767479 43314 767488
rect 43168 766420 43220 766426
rect 43168 766362 43220 766368
rect 43166 766320 43222 766329
rect 43166 766255 43222 766264
rect 43076 754928 43128 754934
rect 43076 754870 43128 754876
rect 43076 754792 43128 754798
rect 43076 754734 43128 754740
rect 43088 746978 43116 754734
rect 43180 753098 43208 766255
rect 43272 757654 43300 767479
rect 43260 757648 43312 757654
rect 43260 757590 43312 757596
rect 43260 757512 43312 757518
rect 43260 757454 43312 757460
rect 43168 753092 43220 753098
rect 43168 753034 43220 753040
rect 43168 749148 43220 749154
rect 43168 749090 43220 749096
rect 43076 746972 43128 746978
rect 43076 746914 43128 746920
rect 43180 742626 43208 749090
rect 43168 742620 43220 742626
rect 43168 742562 43220 742568
rect 43272 730522 43300 757454
rect 43260 730516 43312 730522
rect 43260 730458 43312 730464
rect 43364 729745 43392 773570
rect 43456 772449 43484 797830
rect 43536 797700 43588 797706
rect 43536 797642 43588 797648
rect 43442 772440 43498 772449
rect 43442 772375 43498 772384
rect 43548 770409 43576 797642
rect 43640 790702 43668 808687
rect 43732 793014 43760 810018
rect 43824 799814 43852 810727
rect 43902 809976 43958 809985
rect 43902 809911 43958 809920
rect 43812 799808 43864 799814
rect 43812 799750 43864 799756
rect 43812 799672 43864 799678
rect 43812 799614 43864 799620
rect 43824 798182 43852 799614
rect 43812 798176 43864 798182
rect 43812 798118 43864 798124
rect 43812 798040 43864 798046
rect 43812 797982 43864 797988
rect 43720 793008 43772 793014
rect 43720 792950 43772 792956
rect 43628 790696 43680 790702
rect 43628 790638 43680 790644
rect 43824 789342 43852 797982
rect 43916 790158 43944 809911
rect 43904 790152 43956 790158
rect 43904 790094 43956 790100
rect 43812 789336 43864 789342
rect 43812 789278 43864 789284
rect 44008 773634 44036 927143
rect 44086 810384 44142 810393
rect 44086 810319 44142 810328
rect 44100 799898 44128 810319
rect 44272 800488 44324 800494
rect 44272 800430 44324 800436
rect 44100 799870 44220 799898
rect 44088 799808 44140 799814
rect 44088 799750 44140 799756
rect 44100 786282 44128 799750
rect 44192 798046 44220 799870
rect 44180 798040 44232 798046
rect 44180 797982 44232 797988
rect 44284 797298 44312 800430
rect 44272 797292 44324 797298
rect 44272 797234 44324 797240
rect 44088 786276 44140 786282
rect 44088 786218 44140 786224
rect 43996 773628 44048 773634
rect 43996 773570 44048 773576
rect 43534 770400 43590 770409
rect 43534 770335 43590 770344
rect 43718 769176 43774 769185
rect 43718 769111 43774 769120
rect 43534 765912 43590 765921
rect 43534 765847 43590 765856
rect 43442 765096 43498 765105
rect 43442 765031 43498 765040
rect 43456 750650 43484 765031
rect 43548 751126 43576 765847
rect 43628 757648 43680 757654
rect 43628 757590 43680 757596
rect 43536 751120 43588 751126
rect 43536 751062 43588 751068
rect 43444 750644 43496 750650
rect 43444 750586 43496 750592
rect 43444 750508 43496 750514
rect 43444 750450 43496 750456
rect 43456 746298 43484 750450
rect 43444 746292 43496 746298
rect 43444 746234 43496 746240
rect 43640 743306 43668 757590
rect 43732 749154 43760 769111
rect 44086 768768 44142 768777
rect 44086 768703 44142 768712
rect 44100 767294 44128 768703
rect 43916 767266 44128 767294
rect 43812 766420 43864 766426
rect 43812 766362 43864 766368
rect 43824 749834 43852 766362
rect 43812 749828 43864 749834
rect 43812 749770 43864 749776
rect 43720 749148 43772 749154
rect 43720 749090 43772 749096
rect 43720 749012 43772 749018
rect 43720 748954 43772 748960
rect 43732 746774 43760 748954
rect 43720 746768 43772 746774
rect 43720 746710 43772 746716
rect 43916 745482 43944 767266
rect 44086 767136 44142 767145
rect 44086 767071 44142 767080
rect 43994 765504 44050 765513
rect 43994 765439 44050 765448
rect 44008 754798 44036 765439
rect 43996 754792 44048 754798
rect 43996 754734 44048 754740
rect 44100 754730 44128 767071
rect 44180 756560 44232 756566
rect 44180 756502 44232 756508
rect 44088 754724 44140 754730
rect 44088 754666 44140 754672
rect 44192 754610 44220 756502
rect 44008 754582 44220 754610
rect 44008 747974 44036 754582
rect 44088 754520 44140 754526
rect 44088 754462 44140 754468
rect 44100 750514 44128 754462
rect 44088 750508 44140 750514
rect 44088 750450 44140 750456
rect 44008 747946 44128 747974
rect 43904 745476 43956 745482
rect 43904 745418 43956 745424
rect 44100 743782 44128 747946
rect 44088 743776 44140 743782
rect 44088 743718 44140 743724
rect 43628 743300 43680 743306
rect 43628 743242 43680 743248
rect 44178 730144 44234 730153
rect 44178 730079 44234 730088
rect 43350 729736 43406 729745
rect 43350 729671 43406 729680
rect 42524 729292 42576 729298
rect 42524 729234 42576 729240
rect 42984 729292 43036 729298
rect 42984 729234 43036 729240
rect 41786 728920 41842 728929
rect 41786 728855 41788 728864
rect 41840 728855 41842 728864
rect 41788 728826 41840 728832
rect 42536 728754 42564 729234
rect 42524 728748 42576 728754
rect 42524 728690 42576 728696
rect 39394 728240 39450 728249
rect 39394 728175 39450 728184
rect 42536 727297 42564 728690
rect 43718 728512 43774 728521
rect 43718 728447 43774 728456
rect 42522 727288 42578 727297
rect 42522 727223 42578 727232
rect 43626 726880 43682 726889
rect 43626 726815 43682 726824
rect 43074 726472 43130 726481
rect 43074 726407 43130 726416
rect 41878 724840 41934 724849
rect 41878 724775 41934 724784
rect 41326 723752 41382 723761
rect 41326 723687 41382 723696
rect 30378 720488 30434 720497
rect 30378 720423 30434 720432
rect 30392 720089 30420 720423
rect 30378 720080 30434 720089
rect 30378 720015 30434 720024
rect 41340 717602 41368 723687
rect 41510 720896 41566 720905
rect 41510 720831 41566 720840
rect 41524 720089 41552 720831
rect 41510 720080 41566 720089
rect 41510 720015 41512 720024
rect 41564 720015 41566 720024
rect 41512 719986 41564 719992
rect 41328 717596 41380 717602
rect 41328 717538 41380 717544
rect 41892 713862 41920 724775
rect 42890 724432 42946 724441
rect 42890 724367 42946 724376
rect 42798 723208 42854 723217
rect 42798 723143 42854 723152
rect 42524 716644 42576 716650
rect 42524 716586 42576 716592
rect 41880 713856 41932 713862
rect 41880 713798 41932 713804
rect 41880 713584 41932 713590
rect 41880 713526 41932 713532
rect 41892 713048 41920 713526
rect 42156 711680 42208 711686
rect 42156 711622 42208 711628
rect 42168 711212 42196 711622
rect 42536 711142 42564 716586
rect 42156 711136 42208 711142
rect 42156 711078 42208 711084
rect 42524 711136 42576 711142
rect 42524 711078 42576 711084
rect 42168 710561 42196 711078
rect 42812 709918 42840 723143
rect 42156 709912 42208 709918
rect 42156 709854 42208 709860
rect 42800 709912 42852 709918
rect 42800 709854 42852 709860
rect 42168 709376 42196 709854
rect 42800 709776 42852 709782
rect 42800 709718 42852 709724
rect 42156 708484 42208 708490
rect 42156 708426 42208 708432
rect 42168 708152 42196 708426
rect 42156 708076 42208 708082
rect 42156 708018 42208 708024
rect 42168 707540 42196 708018
rect 42156 707260 42208 707266
rect 42156 707202 42208 707208
rect 42168 706860 42196 707202
rect 42156 706784 42208 706790
rect 42156 706726 42208 706732
rect 42168 706316 42196 706726
rect 42248 704880 42300 704886
rect 42248 704822 42300 704828
rect 42064 704268 42116 704274
rect 42064 704210 42116 704216
rect 42076 703868 42104 704210
rect 42260 703202 42288 704822
rect 42182 703174 42288 703202
rect 42064 702908 42116 702914
rect 42064 702850 42116 702856
rect 42076 702576 42104 702850
rect 42064 702432 42116 702438
rect 42064 702374 42116 702380
rect 42076 702032 42104 702374
rect 42156 700460 42208 700466
rect 42156 700402 42208 700408
rect 42168 700165 42196 700402
rect 42156 700052 42208 700058
rect 42156 699994 42208 700000
rect 42168 699516 42196 699994
rect 42812 699446 42840 709718
rect 42904 700058 42932 724367
rect 42982 723616 43038 723625
rect 42982 723551 43038 723560
rect 42996 704886 43024 723551
rect 43088 711686 43116 726407
rect 43166 726064 43222 726073
rect 43166 725999 43222 726008
rect 43076 711680 43128 711686
rect 43076 711622 43128 711628
rect 43076 711544 43128 711550
rect 43076 711486 43128 711492
rect 43088 706790 43116 711486
rect 43180 709782 43208 725999
rect 43534 725656 43590 725665
rect 43534 725591 43590 725600
rect 43350 725248 43406 725257
rect 43350 725183 43406 725192
rect 43258 721576 43314 721585
rect 43258 721511 43314 721520
rect 43168 709776 43220 709782
rect 43168 709718 43220 709724
rect 43168 709640 43220 709646
rect 43168 709582 43220 709588
rect 43076 706784 43128 706790
rect 43076 706726 43128 706732
rect 42984 704880 43036 704886
rect 42984 704822 43036 704828
rect 42892 700052 42944 700058
rect 42892 699994 42944 700000
rect 42064 699440 42116 699446
rect 42064 699382 42116 699388
rect 42800 699440 42852 699446
rect 42800 699382 42852 699388
rect 42076 698904 42104 699382
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 41512 688424 41564 688430
rect 41510 688392 41512 688401
rect 41564 688392 41566 688401
rect 41510 688327 41566 688336
rect 41696 687880 41748 687886
rect 41696 687822 41748 687828
rect 41708 687585 41736 687822
rect 41788 687744 41840 687750
rect 41786 687712 41788 687721
rect 41840 687712 41842 687721
rect 41786 687647 41842 687656
rect 41694 687576 41750 687585
rect 41694 687511 41750 687520
rect 42798 685264 42854 685273
rect 42798 685199 42854 685208
rect 42812 684486 42840 685199
rect 43180 684865 43208 709582
rect 43272 708490 43300 721511
rect 43364 711550 43392 725183
rect 43442 722800 43498 722809
rect 43442 722735 43498 722744
rect 43352 711544 43404 711550
rect 43352 711486 43404 711492
rect 43260 708484 43312 708490
rect 43260 708426 43312 708432
rect 43456 708082 43484 722735
rect 43444 708076 43496 708082
rect 43444 708018 43496 708024
rect 43548 702438 43576 725591
rect 43536 702432 43588 702438
rect 43536 702374 43588 702380
rect 43640 700466 43668 726815
rect 43732 709646 43760 728447
rect 43902 722392 43958 722401
rect 43902 722327 43958 722336
rect 43812 717596 43864 717602
rect 43812 717538 43864 717544
rect 43720 709640 43772 709646
rect 43720 709582 43772 709588
rect 43824 702914 43852 717538
rect 43916 704274 43944 722327
rect 44086 721984 44142 721993
rect 44086 721919 44142 721928
rect 44100 707266 44128 721919
rect 44088 707260 44140 707266
rect 44088 707202 44140 707208
rect 43904 704268 43956 704274
rect 43904 704210 43956 704216
rect 43812 702908 43864 702914
rect 43812 702850 43864 702856
rect 43628 700460 43680 700466
rect 43628 700402 43680 700408
rect 44192 686497 44220 730079
rect 44272 728884 44324 728890
rect 44272 728826 44324 728832
rect 44178 686488 44234 686497
rect 44178 686423 44234 686432
rect 44284 686089 44312 728826
rect 44362 727696 44418 727705
rect 44362 727631 44418 727640
rect 44270 686080 44326 686089
rect 44270 686015 44326 686024
rect 43442 685672 43498 685681
rect 43442 685607 43498 685616
rect 43166 684856 43222 684865
rect 43166 684791 43222 684800
rect 42800 684480 42852 684486
rect 42800 684422 42852 684428
rect 42890 684448 42946 684457
rect 41694 681864 41750 681873
rect 41340 681822 41694 681850
rect 41340 673470 41368 681822
rect 41694 681799 41750 681808
rect 41878 681592 41934 681601
rect 41878 681527 41934 681536
rect 41786 678736 41842 678745
rect 41786 678671 41842 678680
rect 41800 678230 41828 678671
rect 41788 678224 41840 678230
rect 41788 678166 41840 678172
rect 41786 677920 41842 677929
rect 41786 677855 41842 677864
rect 41800 677113 41828 677855
rect 41786 677104 41842 677113
rect 41786 677039 41788 677048
rect 41840 677039 41842 677048
rect 41788 677010 41840 677016
rect 41328 673464 41380 673470
rect 41328 673406 41380 673412
rect 41892 670614 41920 681527
rect 41970 678328 42026 678337
rect 41970 678263 42026 678272
rect 41984 670614 42012 678263
rect 41880 670608 41932 670614
rect 41880 670550 41932 670556
rect 41972 670608 42024 670614
rect 41972 670550 42024 670556
rect 42708 670608 42760 670614
rect 42708 670550 42760 670556
rect 41880 670404 41932 670410
rect 41880 670346 41932 670352
rect 41892 669868 41920 670346
rect 42064 668500 42116 668506
rect 42064 668442 42116 668448
rect 42076 668032 42104 668442
rect 42156 667752 42208 667758
rect 42156 667694 42208 667700
rect 42168 667352 42196 667694
rect 42156 666732 42208 666738
rect 42156 666674 42208 666680
rect 42168 666165 42196 666674
rect 42720 665446 42748 670550
rect 42156 665440 42208 665446
rect 42156 665382 42208 665388
rect 42708 665440 42760 665446
rect 42708 665382 42760 665388
rect 42168 664972 42196 665382
rect 42156 664692 42208 664698
rect 42156 664634 42208 664640
rect 42168 664325 42196 664634
rect 42156 664216 42208 664222
rect 42156 664158 42208 664164
rect 42168 663680 42196 664158
rect 42156 663604 42208 663610
rect 42156 663546 42208 663552
rect 42168 663136 42196 663546
rect 42156 661088 42208 661094
rect 42156 661030 42208 661036
rect 42168 660620 42196 661030
rect 42156 660544 42208 660550
rect 42156 660486 42208 660492
rect 42168 660008 42196 660486
rect 42156 659932 42208 659938
rect 42156 659874 42208 659880
rect 42168 659357 42196 659874
rect 42156 659048 42208 659054
rect 42156 658990 42208 658996
rect 42168 658784 42196 658990
rect 42156 657280 42208 657286
rect 42156 657222 42208 657228
rect 42168 656948 42196 657222
rect 42156 656872 42208 656878
rect 42156 656814 42208 656820
rect 42168 656336 42196 656814
rect 42156 656192 42208 656198
rect 42156 656134 42208 656140
rect 42168 655656 42196 656134
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 41512 645176 41564 645182
rect 41510 645144 41512 645153
rect 41564 645144 41566 645153
rect 41510 645079 41566 645088
rect 41512 644768 41564 644774
rect 41510 644736 41512 644745
rect 41564 644736 41566 644745
rect 41510 644671 41566 644680
rect 41512 644632 41564 644638
rect 41512 644574 41564 644580
rect 41524 644337 41552 644574
rect 41510 644328 41566 644337
rect 41510 644263 41566 644272
rect 41510 643512 41566 643521
rect 41510 643447 41512 643456
rect 41564 643447 41566 643456
rect 41512 643418 41564 643424
rect 42812 641889 42840 684422
rect 42890 684383 42946 684392
rect 42904 643210 42932 684383
rect 43350 683632 43406 683641
rect 43350 683567 43406 683576
rect 42982 682816 43038 682825
rect 42982 682751 43038 682760
rect 42996 656198 43024 682751
rect 43166 680776 43222 680785
rect 43166 680711 43222 680720
rect 43076 673464 43128 673470
rect 43076 673406 43128 673412
rect 43088 663610 43116 673406
rect 43076 663604 43128 663610
rect 43076 663546 43128 663552
rect 43180 659938 43208 680711
rect 43260 678224 43312 678230
rect 43260 678166 43312 678172
rect 43272 664222 43300 678166
rect 43260 664216 43312 664222
rect 43260 664158 43312 664164
rect 43168 659932 43220 659938
rect 43168 659874 43220 659880
rect 43364 657286 43392 683567
rect 43352 657280 43404 657286
rect 43352 657222 43404 657228
rect 42984 656192 43036 656198
rect 42984 656134 43036 656140
rect 42892 643204 42944 643210
rect 42892 643146 42944 643152
rect 42798 641880 42854 641889
rect 42798 641815 42854 641824
rect 42904 641073 42932 643146
rect 43456 643113 43484 685607
rect 44376 684049 44404 727631
rect 44362 684040 44418 684049
rect 44362 683975 44418 683984
rect 43994 683224 44050 683233
rect 43994 683159 44050 683168
rect 43810 682408 43866 682417
rect 43810 682343 43866 682352
rect 43718 681184 43774 681193
rect 43718 681119 43774 681128
rect 43626 680368 43682 680377
rect 43626 680303 43682 680312
rect 43534 679552 43590 679561
rect 43534 679487 43590 679496
rect 43548 664698 43576 679487
rect 43536 664692 43588 664698
rect 43536 664634 43588 664640
rect 43640 660550 43668 680303
rect 43628 660544 43680 660550
rect 43628 660486 43680 660492
rect 43732 656878 43760 681119
rect 43824 659054 43852 682343
rect 43902 679960 43958 679969
rect 43902 679895 43958 679904
rect 43916 666738 43944 679895
rect 44008 668506 44036 683159
rect 44086 679144 44142 679153
rect 44086 679079 44142 679088
rect 44100 670682 44128 679079
rect 44180 670744 44232 670750
rect 44180 670686 44232 670692
rect 44088 670676 44140 670682
rect 44088 670618 44140 670624
rect 44192 670290 44220 670686
rect 44100 670262 44220 670290
rect 43996 668500 44048 668506
rect 43996 668442 44048 668448
rect 44100 667758 44128 670262
rect 44180 670200 44232 670206
rect 44180 670142 44232 670148
rect 44088 667752 44140 667758
rect 44088 667694 44140 667700
rect 44192 667570 44220 670142
rect 44100 667542 44220 667570
rect 43904 666732 43956 666738
rect 43904 666674 43956 666680
rect 44100 661094 44128 667542
rect 44088 661088 44140 661094
rect 44088 661030 44140 661036
rect 43812 659048 43864 659054
rect 43812 658990 43864 658996
rect 43720 656872 43772 656878
rect 43720 656814 43772 656820
rect 44364 643476 44416 643482
rect 44364 643418 44416 643424
rect 43442 643104 43498 643113
rect 43442 643039 43498 643048
rect 44270 642016 44326 642025
rect 44270 641951 44326 641960
rect 42890 641064 42946 641073
rect 42890 640999 42946 641008
rect 43074 640384 43130 640393
rect 43074 640319 43130 640328
rect 42798 639432 42854 639441
rect 42798 639367 42854 639376
rect 41786 638412 41842 638421
rect 41786 638347 41842 638356
rect 33046 634944 33102 634953
rect 33046 634879 33102 634888
rect 30378 634128 30434 634137
rect 30378 634063 30434 634072
rect 30392 633729 30420 634063
rect 30378 633720 30434 633729
rect 30378 633655 30434 633664
rect 33060 627910 33088 634879
rect 41510 634536 41566 634545
rect 41510 634471 41566 634480
rect 41524 633729 41552 634471
rect 41510 633720 41566 633729
rect 41510 633655 41512 633664
rect 41564 633655 41566 633664
rect 41512 633626 41564 633632
rect 33048 627904 33100 627910
rect 33048 627846 33100 627852
rect 41800 627434 41828 638347
rect 42524 627904 42576 627910
rect 42524 627846 42576 627852
rect 41788 627428 41840 627434
rect 41788 627370 41840 627376
rect 41788 627088 41840 627094
rect 41788 627030 41840 627036
rect 41800 626620 41828 627030
rect 42156 625320 42208 625326
rect 42156 625262 42208 625268
rect 42168 624784 42196 625262
rect 42156 624708 42208 624714
rect 42156 624650 42208 624656
rect 42168 624172 42196 624650
rect 42156 623484 42208 623490
rect 42156 623426 42208 623432
rect 42168 622948 42196 623426
rect 42536 622198 42564 627846
rect 42064 622192 42116 622198
rect 42064 622134 42116 622140
rect 42524 622192 42576 622198
rect 42524 622134 42576 622140
rect 42076 621792 42104 622134
rect 42156 621512 42208 621518
rect 42156 621454 42208 621460
rect 42168 621112 42196 621454
rect 42064 621036 42116 621042
rect 42064 620978 42116 620984
rect 42076 620500 42104 620978
rect 42064 620220 42116 620226
rect 42064 620162 42116 620168
rect 42076 619956 42104 620162
rect 42248 619064 42300 619070
rect 42248 619006 42300 619012
rect 42156 617908 42208 617914
rect 42156 617850 42208 617856
rect 42168 617440 42196 617850
rect 42064 617160 42116 617166
rect 42064 617102 42116 617108
rect 42076 616828 42104 617102
rect 42156 616684 42208 616690
rect 42156 616626 42208 616632
rect 42168 616148 42196 616626
rect 42260 615618 42288 619006
rect 42182 615590 42288 615618
rect 42156 614236 42208 614242
rect 42156 614178 42208 614184
rect 42168 613768 42196 614178
rect 42156 613692 42208 613698
rect 42156 613634 42208 613640
rect 42168 613121 42196 613634
rect 42812 613018 42840 639367
rect 42982 637800 43038 637809
rect 42982 637735 43038 637744
rect 42890 636576 42946 636585
rect 42890 636511 42946 636520
rect 42904 623490 42932 636511
rect 42892 623484 42944 623490
rect 42892 623426 42944 623432
rect 42996 613698 43024 637735
rect 43088 614242 43116 640319
rect 43534 639840 43590 639849
rect 43534 639775 43590 639784
rect 43166 639024 43222 639033
rect 43166 638959 43222 638968
rect 43180 619070 43208 638959
rect 43442 638616 43498 638625
rect 43442 638551 43498 638560
rect 43350 636168 43406 636177
rect 43350 636103 43406 636112
rect 43258 635352 43314 635361
rect 43258 635287 43314 635296
rect 43272 621042 43300 635287
rect 43364 621518 43392 636103
rect 43352 621512 43404 621518
rect 43352 621454 43404 621460
rect 43260 621036 43312 621042
rect 43260 620978 43312 620984
rect 43456 620226 43484 638551
rect 43548 625326 43576 639775
rect 43718 637664 43774 637673
rect 43718 637599 43774 637608
rect 43626 635760 43682 635769
rect 43626 635695 43682 635704
rect 43536 625320 43588 625326
rect 43536 625262 43588 625268
rect 43444 620220 43496 620226
rect 43444 620162 43496 620168
rect 43168 619064 43220 619070
rect 43168 619006 43220 619012
rect 43640 617914 43668 635695
rect 43628 617908 43680 617914
rect 43628 617850 43680 617856
rect 43732 616690 43760 637599
rect 43810 636984 43866 636993
rect 43810 636919 43866 636928
rect 43824 617166 43852 636919
rect 43904 629332 43956 629338
rect 43904 629274 43956 629280
rect 43916 624714 43944 629274
rect 43904 624708 43956 624714
rect 43904 624650 43956 624656
rect 43812 617160 43864 617166
rect 43812 617102 43864 617108
rect 43720 616684 43772 616690
rect 43720 616626 43772 616632
rect 43076 614236 43128 614242
rect 43076 614178 43128 614184
rect 42984 613692 43036 613698
rect 42984 613634 43036 613640
rect 42156 613012 42208 613018
rect 42156 612954 42208 612960
rect 42800 613012 42852 613018
rect 42800 612954 42852 612960
rect 42168 612476 42196 612954
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 41512 601928 41564 601934
rect 41510 601896 41512 601905
rect 41564 601896 41566 601905
rect 41510 601831 41566 601840
rect 41512 601520 41564 601526
rect 41510 601488 41512 601497
rect 41564 601488 41566 601497
rect 41510 601423 41566 601432
rect 43074 600536 43130 600545
rect 43074 600471 43130 600480
rect 41512 599888 41564 599894
rect 41510 599856 41512 599865
rect 41564 599856 41566 599865
rect 41510 599791 41566 599800
rect 41510 599040 41566 599049
rect 41510 598975 41512 598984
rect 41564 598975 41566 598984
rect 41512 598946 41564 598952
rect 42430 598088 42486 598097
rect 42430 598023 42486 598032
rect 41878 595232 41934 595241
rect 41878 595167 41934 595176
rect 41326 594144 41382 594153
rect 41326 594079 41382 594088
rect 29918 591288 29974 591297
rect 29918 591223 29974 591232
rect 29932 590889 29960 591223
rect 29918 590880 29974 590889
rect 29918 590815 29974 590824
rect 30378 590880 30434 590889
rect 30378 590815 30434 590824
rect 30392 590481 30420 590815
rect 30378 590472 30434 590481
rect 30378 590407 30434 590416
rect 41340 585206 41368 594079
rect 41328 585200 41380 585206
rect 41328 585142 41380 585148
rect 41892 584254 41920 595167
rect 41880 584248 41932 584254
rect 41880 584190 41932 584196
rect 41880 583976 41932 583982
rect 41880 583918 41932 583924
rect 41892 583440 41920 583918
rect 42444 583710 42472 598023
rect 42890 596864 42946 596873
rect 42890 596799 42946 596808
rect 42798 593600 42854 593609
rect 42798 593535 42854 593544
rect 42706 591968 42762 591977
rect 42706 591903 42762 591912
rect 42432 583704 42484 583710
rect 42432 583646 42484 583652
rect 42156 582140 42208 582146
rect 42156 582082 42208 582088
rect 42168 581604 42196 582082
rect 42156 581324 42208 581330
rect 42156 581266 42208 581272
rect 42168 580961 42196 581266
rect 42156 580304 42208 580310
rect 42156 580246 42208 580252
rect 42168 579768 42196 580246
rect 42720 579018 42748 591903
rect 42812 580310 42840 593535
rect 42904 582146 42932 596799
rect 42982 594008 43038 594017
rect 42982 593943 43038 593952
rect 42892 582140 42944 582146
rect 42892 582082 42944 582088
rect 42800 580304 42852 580310
rect 42800 580246 42852 580252
rect 42156 579012 42208 579018
rect 42156 578954 42208 578960
rect 42708 579012 42760 579018
rect 42708 578954 42760 578960
rect 42168 578544 42196 578954
rect 42156 578468 42208 578474
rect 42156 578410 42208 578416
rect 42168 577932 42196 578410
rect 42156 577856 42208 577862
rect 42156 577798 42208 577804
rect 42168 577281 42196 577798
rect 42156 576972 42208 576978
rect 42156 576914 42208 576920
rect 42168 576708 42196 576914
rect 42156 574728 42208 574734
rect 42156 574670 42208 574676
rect 42168 574260 42196 574670
rect 42996 574122 43024 593943
rect 42156 574116 42208 574122
rect 42156 574058 42208 574064
rect 42984 574116 43036 574122
rect 42984 574058 43036 574064
rect 42168 573580 42196 574058
rect 42156 573504 42208 573510
rect 42156 573446 42208 573452
rect 42168 572968 42196 573446
rect 42064 572892 42116 572898
rect 42064 572834 42116 572840
rect 42076 572424 42104 572834
rect 42064 570920 42116 570926
rect 42064 570862 42116 570868
rect 42076 570588 42104 570862
rect 42156 570444 42208 570450
rect 42156 570386 42208 570392
rect 42168 569908 42196 570386
rect 42064 569628 42116 569634
rect 42064 569570 42116 569576
rect 42076 569296 42104 569570
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 41512 558816 41564 558822
rect 41510 558784 41512 558793
rect 41564 558784 41566 558793
rect 41510 558719 41566 558728
rect 41512 558340 41564 558346
rect 41512 558282 41564 558288
rect 41524 557977 41552 558282
rect 41788 558272 41840 558278
rect 41788 558214 41840 558220
rect 41800 558113 41828 558214
rect 41786 558104 41842 558113
rect 41786 558039 41842 558048
rect 41510 557968 41566 557977
rect 41510 557903 41566 557912
rect 43088 556889 43116 600471
rect 43352 599004 43404 599010
rect 43352 598946 43404 598952
rect 43258 596456 43314 596465
rect 43258 596391 43314 596400
rect 43166 594824 43222 594833
rect 43166 594759 43222 594768
rect 43180 583914 43208 594759
rect 43272 592482 43300 596391
rect 43260 592476 43312 592482
rect 43260 592418 43312 592424
rect 43258 592376 43314 592385
rect 43258 592311 43314 592320
rect 43168 583908 43220 583914
rect 43168 583850 43220 583856
rect 43272 583794 43300 592311
rect 43180 583766 43300 583794
rect 43180 577862 43208 583766
rect 43260 583704 43312 583710
rect 43260 583646 43312 583652
rect 43168 577856 43220 577862
rect 43168 577798 43220 577804
rect 43074 556880 43130 556889
rect 43074 556815 43130 556824
rect 43272 554774 43300 583646
rect 43364 556481 43392 598946
rect 44284 598505 44312 641951
rect 44376 600137 44404 643418
rect 44454 642288 44510 642297
rect 44454 642223 44510 642232
rect 44362 600128 44418 600137
rect 44362 600063 44418 600072
rect 44468 599894 44496 642223
rect 44638 641472 44694 641481
rect 44638 641407 44694 641416
rect 44456 599888 44508 599894
rect 44456 599830 44508 599836
rect 44270 598496 44326 598505
rect 44270 598431 44326 598440
rect 44652 597689 44680 641407
rect 44638 597680 44694 597689
rect 44638 597615 44694 597624
rect 43810 597272 43866 597281
rect 43810 597207 43866 597216
rect 43442 595640 43498 595649
rect 43442 595575 43498 595584
rect 43456 592618 43484 595575
rect 43626 593192 43682 593201
rect 43626 593127 43682 593136
rect 43444 592612 43496 592618
rect 43444 592554 43496 592560
rect 43444 592476 43496 592482
rect 43444 592418 43496 592424
rect 43456 585134 43484 592418
rect 43456 585106 43576 585134
rect 43444 583908 43496 583914
rect 43444 583850 43496 583856
rect 43456 570450 43484 583850
rect 43444 570444 43496 570450
rect 43444 570386 43496 570392
rect 43548 569634 43576 585106
rect 43640 578474 43668 593127
rect 43718 592784 43774 592793
rect 43718 592719 43774 592728
rect 43628 578468 43680 578474
rect 43628 578410 43680 578416
rect 43732 574734 43760 592719
rect 43720 574728 43772 574734
rect 43720 574670 43772 574676
rect 43824 570926 43852 597207
rect 43902 596048 43958 596057
rect 43902 595983 43958 595992
rect 43916 572898 43944 595983
rect 43996 592612 44048 592618
rect 43996 592554 44048 592560
rect 44008 576978 44036 592554
rect 44088 585200 44140 585206
rect 44088 585142 44140 585148
rect 44180 585200 44232 585206
rect 44180 585142 44232 585148
rect 43996 576972 44048 576978
rect 43996 576914 44048 576920
rect 44100 573510 44128 585142
rect 44192 581330 44220 585142
rect 44180 581324 44232 581330
rect 44180 581266 44232 581272
rect 44088 573504 44140 573510
rect 44088 573446 44140 573452
rect 43904 572892 43956 572898
rect 43904 572834 43956 572840
rect 43812 570920 43864 570926
rect 43812 570862 43864 570868
rect 43536 569628 43588 569634
rect 43536 569570 43588 569576
rect 43350 556472 43406 556481
rect 43350 556407 43406 556416
rect 43180 554746 43300 554774
rect 43180 554441 43208 554746
rect 43166 554432 43222 554441
rect 43166 554367 43222 554376
rect 43534 554024 43590 554033
rect 43534 553959 43590 553968
rect 42706 553616 42762 553625
rect 42706 553551 42762 553560
rect 41786 551984 41842 551993
rect 41786 551919 41842 551928
rect 41602 548992 41658 549001
rect 41602 548927 41658 548936
rect 41510 548584 41566 548593
rect 41510 548519 41566 548528
rect 41418 548176 41474 548185
rect 41418 548111 41474 548120
rect 30470 547768 30526 547777
rect 30470 547703 30526 547712
rect 30484 547369 30512 547703
rect 41432 547369 41460 548111
rect 30470 547360 30526 547369
rect 30470 547295 30526 547304
rect 41418 547360 41474 547369
rect 41418 547295 41420 547304
rect 41472 547295 41474 547304
rect 41420 547266 41472 547272
rect 41524 542502 41552 548519
rect 41616 543182 41644 548927
rect 41604 543176 41656 543182
rect 41604 543118 41656 543124
rect 41512 542496 41564 542502
rect 41512 542438 41564 542444
rect 41800 541074 41828 551919
rect 41788 541068 41840 541074
rect 41788 541010 41840 541016
rect 41788 540796 41840 540802
rect 41788 540738 41840 540744
rect 41800 540260 41828 540738
rect 42720 538966 42748 553551
rect 43350 553208 43406 553217
rect 43350 553143 43406 553152
rect 42982 552800 43038 552809
rect 42982 552735 43038 552744
rect 42890 550352 42946 550361
rect 42890 550287 42946 550296
rect 42800 542496 42852 542502
rect 42800 542438 42852 542444
rect 42064 538960 42116 538966
rect 42064 538902 42116 538908
rect 42708 538960 42760 538966
rect 42708 538902 42760 538908
rect 42076 538424 42104 538902
rect 42156 538144 42208 538150
rect 42156 538086 42208 538092
rect 42168 537744 42196 538086
rect 42064 537124 42116 537130
rect 42064 537066 42116 537072
rect 42076 536588 42104 537066
rect 42812 535838 42840 542438
rect 42904 537130 42932 550287
rect 42892 537124 42944 537130
rect 42892 537066 42944 537072
rect 42996 537010 43024 552735
rect 43166 552392 43222 552401
rect 43166 552327 43222 552336
rect 43074 551168 43130 551177
rect 43074 551103 43130 551112
rect 42904 536982 43024 537010
rect 42156 535832 42208 535838
rect 42156 535774 42208 535780
rect 42800 535832 42852 535838
rect 42800 535774 42852 535780
rect 42168 535364 42196 535774
rect 42064 535084 42116 535090
rect 42064 535026 42116 535032
rect 42076 534752 42104 535026
rect 42156 534608 42208 534614
rect 42156 534550 42208 534556
rect 42168 534072 42196 534550
rect 42156 533792 42208 533798
rect 42156 533734 42208 533740
rect 42168 533528 42196 533734
rect 42156 531480 42208 531486
rect 42156 531422 42208 531428
rect 42168 531045 42196 531422
rect 42156 530732 42208 530738
rect 42156 530674 42208 530680
rect 42168 530400 42196 530674
rect 42156 530324 42208 530330
rect 42156 530266 42208 530272
rect 42168 529757 42196 530266
rect 42904 529650 42932 536982
rect 42984 536920 43036 536926
rect 42984 536862 43036 536868
rect 42156 529644 42208 529650
rect 42156 529586 42208 529592
rect 42892 529644 42944 529650
rect 42892 529586 42944 529592
rect 42168 529205 42196 529586
rect 42076 527270 42104 527340
rect 42064 527264 42116 527270
rect 42064 527206 42116 527212
rect 42156 527196 42208 527202
rect 42156 527138 42208 527144
rect 42168 526728 42196 527138
rect 42996 526658 43024 536862
rect 43088 530330 43116 551103
rect 43180 533798 43208 552327
rect 43260 543176 43312 543182
rect 43260 543118 43312 543124
rect 43272 534614 43300 543118
rect 43364 536926 43392 553143
rect 43442 549944 43498 549953
rect 43442 549879 43498 549888
rect 43352 536920 43404 536926
rect 43352 536862 43404 536868
rect 43352 536784 43404 536790
rect 43352 536726 43404 536732
rect 43260 534608 43312 534614
rect 43260 534550 43312 534556
rect 43168 533792 43220 533798
rect 43168 533734 43220 533740
rect 43076 530324 43128 530330
rect 43076 530266 43128 530272
rect 43364 527270 43392 536726
rect 43456 535090 43484 549879
rect 43548 536790 43576 553959
rect 43626 551576 43682 551585
rect 43626 551511 43682 551520
rect 43536 536784 43588 536790
rect 43536 536726 43588 536732
rect 43444 535084 43496 535090
rect 43444 535026 43496 535032
rect 43352 527264 43404 527270
rect 43352 527206 43404 527212
rect 43640 527202 43668 551511
rect 43718 550760 43774 550769
rect 43718 550695 43774 550704
rect 43732 530738 43760 550695
rect 43810 549536 43866 549545
rect 43810 549471 43866 549480
rect 43824 531486 43852 549471
rect 43904 541068 43956 541074
rect 43904 541010 43956 541016
rect 43916 538150 43944 541010
rect 44086 540968 44142 540977
rect 44086 540903 44142 540912
rect 43994 540832 44050 540841
rect 43994 540767 44050 540776
rect 43904 538144 43956 538150
rect 43904 538086 43956 538092
rect 43812 531480 43864 531486
rect 43812 531422 43864 531428
rect 43720 530732 43772 530738
rect 43720 530674 43772 530680
rect 43628 527196 43680 527202
rect 43628 527138 43680 527144
rect 42156 526652 42208 526658
rect 42156 526594 42208 526600
rect 42984 526652 43036 526658
rect 42984 526594 43036 526600
rect 42168 526077 42196 526594
rect 8588 431596 8616 431732
rect 9048 431596 9076 431732
rect 9508 431596 9536 431732
rect 9968 431596 9996 431732
rect 10428 431596 10456 431732
rect 10888 431596 10916 431732
rect 11348 431596 11376 431732
rect 11808 431596 11836 431732
rect 12268 431596 12296 431732
rect 12728 431596 12756 431732
rect 13188 431596 13216 431732
rect 13648 431596 13676 431732
rect 14108 431596 14136 431732
rect 41786 430944 41842 430953
rect 41786 430879 41842 430888
rect 41800 430642 41828 430879
rect 44008 430710 44036 540767
rect 43996 430704 44048 430710
rect 43996 430646 44048 430652
rect 41788 430636 41840 430642
rect 41788 430578 41840 430584
rect 43534 429720 43590 429729
rect 43534 429655 43590 429664
rect 41788 427848 41840 427854
rect 41788 427790 41840 427796
rect 41800 426873 41828 427790
rect 41786 426864 41842 426873
rect 41786 426799 41842 426808
rect 43258 426456 43314 426465
rect 43258 426391 43314 426400
rect 42798 426048 42854 426057
rect 42798 425983 42854 425992
rect 41878 424416 41934 424425
rect 41878 424351 41934 424360
rect 41786 421560 41842 421569
rect 41786 421495 41842 421504
rect 41800 416362 41828 421495
rect 41788 416356 41840 416362
rect 41788 416298 41840 416304
rect 41892 413438 41920 424351
rect 42522 421152 42578 421161
rect 42522 421087 42578 421096
rect 41880 413432 41932 413438
rect 41880 413374 41932 413380
rect 41880 413160 41932 413166
rect 41880 413102 41932 413108
rect 41892 412624 41920 413102
rect 42156 411324 42208 411330
rect 42156 411266 42208 411272
rect 42168 410788 42196 411266
rect 42156 410712 42208 410718
rect 42156 410654 42208 410660
rect 42168 410176 42196 410654
rect 42156 409420 42208 409426
rect 42156 409362 42208 409368
rect 42168 408952 42196 409362
rect 42536 408202 42564 421087
rect 42812 411398 42840 425983
rect 42890 425640 42946 425649
rect 42890 425575 42946 425584
rect 42800 411392 42852 411398
rect 42800 411334 42852 411340
rect 42798 411268 42854 411277
rect 42798 411203 42854 411212
rect 42064 408196 42116 408202
rect 42064 408138 42116 408144
rect 42524 408196 42576 408202
rect 42524 408138 42576 408144
rect 42076 407796 42104 408138
rect 42156 407516 42208 407522
rect 42156 407458 42208 407464
rect 42168 407116 42196 407458
rect 42064 407040 42116 407046
rect 42064 406982 42116 406988
rect 42076 406504 42104 406982
rect 42156 406224 42208 406230
rect 42156 406166 42208 406172
rect 42168 405929 42196 406166
rect 42156 403912 42208 403918
rect 42156 403854 42208 403860
rect 42168 403444 42196 403854
rect 42156 403368 42208 403374
rect 42156 403310 42208 403316
rect 42168 402801 42196 403310
rect 42156 402552 42208 402558
rect 42156 402494 42208 402500
rect 42168 402152 42196 402494
rect 42156 402076 42208 402082
rect 42156 402018 42208 402024
rect 42168 401608 42196 402018
rect 42156 400036 42208 400042
rect 42156 399978 42208 399984
rect 42168 399772 42196 399978
rect 42156 399492 42208 399498
rect 42156 399434 42208 399440
rect 42168 399121 42196 399434
rect 42156 399016 42208 399022
rect 42156 398958 42208 398964
rect 42168 398480 42196 398958
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41512 388000 41564 388006
rect 41510 387968 41512 387977
rect 41564 387968 41566 387977
rect 41510 387903 41566 387912
rect 41788 387456 41840 387462
rect 41788 387398 41840 387404
rect 41800 387297 41828 387398
rect 41786 387288 41842 387297
rect 41786 387223 41842 387232
rect 41512 387184 41564 387190
rect 41510 387152 41512 387161
rect 41564 387152 41566 387161
rect 41510 387087 41566 387096
rect 42812 386442 42840 411203
rect 42904 399022 42932 425575
rect 43166 425232 43222 425241
rect 43166 425167 43222 425176
rect 42982 422784 43038 422793
rect 42982 422719 43038 422728
rect 42996 409426 43024 422719
rect 43076 416356 43128 416362
rect 43076 416298 43128 416304
rect 42984 409420 43036 409426
rect 42984 409362 43036 409368
rect 43088 407046 43116 416298
rect 43076 407040 43128 407046
rect 43076 406982 43128 406988
rect 43180 402082 43208 425167
rect 43168 402076 43220 402082
rect 43168 402018 43220 402024
rect 43272 400042 43300 426391
rect 43442 424824 43498 424833
rect 43442 424759 43498 424768
rect 43350 422376 43406 422385
rect 43350 422311 43406 422320
rect 43364 407522 43392 422311
rect 43352 407516 43404 407522
rect 43352 407458 43404 407464
rect 43456 406230 43484 424759
rect 43548 411505 43576 429655
rect 44008 429321 44036 430646
rect 43994 429312 44050 429321
rect 43994 429247 44050 429256
rect 43718 428496 43774 428505
rect 43718 428431 43774 428440
rect 43626 423192 43682 423201
rect 43626 423127 43682 423136
rect 43534 411496 43590 411505
rect 43534 411431 43590 411440
rect 43444 406224 43496 406230
rect 43444 406166 43496 406172
rect 43640 403374 43668 423127
rect 43628 403368 43680 403374
rect 43628 403310 43680 403316
rect 43260 400036 43312 400042
rect 43260 399978 43312 399984
rect 42892 399016 42944 399022
rect 42892 398958 42944 398964
rect 42800 386436 42852 386442
rect 42800 386378 42852 386384
rect 42812 386073 42840 386378
rect 42798 386064 42854 386073
rect 42798 385999 42854 386008
rect 43732 385665 43760 428431
rect 44100 427854 44128 540903
rect 44088 427848 44140 427854
rect 44088 427790 44140 427796
rect 43902 424008 43958 424017
rect 43902 423943 43958 423952
rect 43810 423600 43866 423609
rect 43810 423535 43866 423544
rect 43824 402558 43852 423535
rect 43812 402552 43864 402558
rect 43812 402494 43864 402500
rect 43916 400214 43944 423943
rect 43994 421968 44050 421977
rect 43994 421903 44050 421912
rect 44008 403918 44036 421903
rect 43996 403912 44048 403918
rect 43996 403854 44048 403860
rect 43824 400186 43944 400214
rect 43824 399498 43852 400186
rect 43812 399492 43864 399498
rect 43812 399434 43864 399440
rect 43718 385656 43774 385665
rect 43718 385591 43774 385600
rect 43534 385248 43590 385257
rect 43534 385183 43590 385192
rect 42982 383208 43038 383217
rect 42982 383143 43038 383152
rect 42706 382800 42762 382809
rect 42706 382735 42762 382744
rect 42338 381168 42394 381177
rect 42338 381103 42394 381112
rect 41510 377768 41566 377777
rect 41510 377703 41566 377712
rect 41418 377360 41474 377369
rect 41418 377295 41474 377304
rect 30470 376952 30526 376961
rect 30470 376887 30526 376896
rect 30484 376553 30512 376887
rect 41432 376553 41460 377295
rect 30470 376544 30526 376553
rect 30470 376479 30526 376488
rect 41418 376544 41474 376553
rect 41418 376479 41420 376488
rect 41472 376479 41474 376488
rect 41420 376450 41472 376456
rect 41524 371482 41552 377703
rect 41512 371476 41564 371482
rect 41512 371418 41564 371424
rect 42352 369986 42380 381103
rect 42156 369980 42208 369986
rect 42156 369922 42208 369928
rect 42340 369980 42392 369986
rect 42340 369922 42392 369928
rect 42168 369444 42196 369922
rect 42720 368150 42748 382735
rect 42890 381984 42946 381993
rect 42890 381919 42946 381928
rect 42798 381576 42854 381585
rect 42798 381511 42854 381520
rect 42812 371822 42840 381511
rect 42800 371816 42852 371822
rect 42800 371758 42852 371764
rect 42800 371476 42852 371482
rect 42800 371418 42852 371424
rect 42156 368144 42208 368150
rect 42156 368086 42208 368092
rect 42708 368144 42760 368150
rect 42708 368086 42760 368092
rect 42168 367608 42196 368086
rect 42168 366858 42196 366961
rect 42156 366852 42208 366858
rect 42156 366794 42208 366800
rect 42156 366308 42208 366314
rect 42156 366250 42208 366256
rect 42168 365772 42196 366250
rect 42812 365022 42840 371418
rect 42156 365016 42208 365022
rect 42156 364958 42208 364964
rect 42800 365016 42852 365022
rect 42800 364958 42852 364964
rect 42168 364548 42196 364958
rect 42156 364472 42208 364478
rect 42156 364414 42208 364420
rect 42168 363936 42196 364414
rect 42156 363860 42208 363866
rect 42156 363802 42208 363808
rect 42168 363256 42196 363802
rect 42156 363180 42208 363186
rect 42156 363122 42208 363128
rect 42168 362712 42196 363122
rect 42064 360732 42116 360738
rect 42064 360674 42116 360680
rect 42076 360264 42104 360674
rect 42156 359984 42208 359990
rect 42156 359926 42208 359932
rect 42168 359584 42196 359926
rect 42156 359508 42208 359514
rect 42156 359450 42208 359456
rect 42168 358972 42196 359450
rect 42904 358834 42932 381919
rect 42064 358828 42116 358834
rect 42064 358770 42116 358776
rect 42892 358828 42944 358834
rect 42892 358770 42944 358776
rect 42076 358428 42104 358770
rect 42996 356998 43024 383143
rect 43074 379536 43130 379545
rect 43074 379471 43130 379480
rect 43088 366314 43116 379471
rect 43258 379128 43314 379137
rect 43258 379063 43314 379072
rect 43166 378312 43222 378321
rect 43166 378247 43222 378256
rect 43076 366308 43128 366314
rect 43076 366250 43128 366256
rect 43180 363866 43208 378247
rect 43272 364478 43300 379063
rect 43442 378720 43498 378729
rect 43442 378655 43498 378664
rect 43352 371816 43404 371822
rect 43352 371758 43404 371764
rect 43260 364472 43312 364478
rect 43260 364414 43312 364420
rect 43168 363860 43220 363866
rect 43168 363802 43220 363808
rect 43364 363186 43392 371758
rect 43352 363180 43404 363186
rect 43352 363122 43404 363128
rect 43456 362930 43484 378655
rect 43088 362902 43484 362930
rect 43088 360738 43116 362902
rect 43168 362840 43220 362846
rect 43168 362782 43220 362788
rect 43076 360732 43128 360738
rect 43076 360674 43128 360680
rect 42064 356992 42116 356998
rect 42064 356934 42116 356940
rect 42984 356992 43036 356998
rect 42984 356934 43036 356940
rect 42076 356592 42104 356934
rect 43180 356318 43208 362782
rect 42156 356312 42208 356318
rect 42156 356254 42208 356260
rect 43168 356312 43220 356318
rect 43168 356254 43220 356260
rect 42168 355912 42196 356254
rect 41786 355736 41842 355745
rect 41786 355671 41842 355680
rect 41800 355300 41828 355671
rect 33046 351928 33102 351937
rect 33046 351863 33102 351872
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 33060 343097 33088 351863
rect 41510 344312 41566 344321
rect 41510 344247 41512 344256
rect 41564 344247 41566 344256
rect 41512 344218 41564 344224
rect 41788 344208 41840 344214
rect 41786 344176 41788 344185
rect 41840 344176 41842 344185
rect 41512 344140 41564 344146
rect 43548 344146 43576 385183
rect 43626 380760 43682 380769
rect 43626 380695 43682 380704
rect 43640 362846 43668 380695
rect 43718 380352 43774 380361
rect 43718 380287 43774 380296
rect 43628 362840 43680 362846
rect 43628 362782 43680 362788
rect 43732 361574 43760 380287
rect 43810 379944 43866 379953
rect 43810 379879 43866 379888
rect 43640 361546 43760 361574
rect 43640 359514 43668 361546
rect 43824 359990 43852 379879
rect 43812 359984 43864 359990
rect 43812 359926 43864 359932
rect 43628 359508 43680 359514
rect 43628 359450 43680 359456
rect 44364 345024 44416 345030
rect 44364 344966 44416 344972
rect 41786 344111 41842 344120
rect 43536 344140 43588 344146
rect 41512 344082 41564 344088
rect 43536 344082 43588 344088
rect 33046 343088 33102 343097
rect 33046 343023 33102 343032
rect 41524 342689 41552 344082
rect 41604 343936 41656 343942
rect 41602 343904 41604 343913
rect 41656 343904 41658 343913
rect 41602 343839 41658 343848
rect 44376 343398 44404 344966
rect 41788 343392 41840 343398
rect 41786 343360 41788 343369
rect 44364 343392 44416 343398
rect 41840 343360 41842 343369
rect 44364 343334 44416 343340
rect 41786 343295 41842 343304
rect 41510 342680 41566 342689
rect 41510 342615 41566 342624
rect 43258 342136 43314 342145
rect 43258 342071 43314 342080
rect 32678 339824 32734 339833
rect 32678 339759 32734 339768
rect 32586 338600 32642 338609
rect 32586 338535 32642 338544
rect 30378 333704 30434 333713
rect 30378 333639 30434 333648
rect 30392 333305 30420 333639
rect 30378 333296 30434 333305
rect 30378 333231 30434 333240
rect 32600 329769 32628 338535
rect 32692 329934 32720 339759
rect 32770 338192 32826 338201
rect 32770 338127 32826 338136
rect 32680 329928 32732 329934
rect 32784 329905 32812 338127
rect 33046 337784 33102 337793
rect 33046 337719 33102 337728
rect 32954 336152 33010 336161
rect 32954 336087 33010 336096
rect 32862 335744 32918 335753
rect 32862 335679 32918 335688
rect 32680 329870 32732 329876
rect 32770 329896 32826 329905
rect 32876 329866 32904 335679
rect 32968 330002 32996 336087
rect 33060 330138 33088 337719
rect 43074 335608 43130 335617
rect 43074 335543 43130 335552
rect 42982 335200 43038 335209
rect 42982 335135 43038 335144
rect 41510 334112 41566 334121
rect 41510 334047 41566 334056
rect 41524 333305 41552 334047
rect 41510 333296 41566 333305
rect 41510 333231 41512 333240
rect 41564 333231 41566 333240
rect 41512 333202 41564 333208
rect 33048 330132 33100 330138
rect 33048 330074 33100 330080
rect 41880 330132 41932 330138
rect 41880 330074 41932 330080
rect 32956 329996 33008 330002
rect 32956 329938 33008 329944
rect 32770 329831 32826 329840
rect 32864 329860 32916 329866
rect 32864 329802 32916 329808
rect 32586 329760 32642 329769
rect 32586 329695 32642 329704
rect 41892 327010 41920 330074
rect 42892 329996 42944 330002
rect 42892 329938 42944 329944
rect 42800 329928 42852 329934
rect 42800 329870 42852 329876
rect 41880 327004 41932 327010
rect 41880 326946 41932 326952
rect 41880 326800 41932 326806
rect 41880 326742 41932 326748
rect 41892 326264 41920 326742
rect 42812 324970 42840 329870
rect 42064 324964 42116 324970
rect 42064 324906 42116 324912
rect 42800 324964 42852 324970
rect 42800 324906 42852 324912
rect 42076 324428 42104 324906
rect 42800 324828 42852 324834
rect 42800 324770 42852 324776
rect 42168 323338 42196 323748
rect 42156 323332 42208 323338
rect 42156 323274 42208 323280
rect 42616 323332 42668 323338
rect 42616 323274 42668 323280
rect 42064 323128 42116 323134
rect 42064 323070 42116 323076
rect 42076 322592 42104 323070
rect 42156 321836 42208 321842
rect 42156 321778 42208 321784
rect 42168 321368 42196 321778
rect 42156 321088 42208 321094
rect 42156 321030 42208 321036
rect 42168 320725 42196 321030
rect 42156 320612 42208 320618
rect 42156 320554 42208 320560
rect 42168 320076 42196 320554
rect 42628 320142 42656 323274
rect 42616 320136 42668 320142
rect 42616 320078 42668 320084
rect 41786 319968 41842 319977
rect 41786 319903 41842 319912
rect 41800 319532 41828 319903
rect 42812 317490 42840 324770
rect 42904 323134 42932 329938
rect 42892 323128 42944 323134
rect 42892 323070 42944 323076
rect 42996 320618 43024 335135
rect 43088 324834 43116 335543
rect 43166 334792 43222 334801
rect 43166 334727 43222 334736
rect 43076 324828 43128 324834
rect 43076 324770 43128 324776
rect 43180 321842 43208 334727
rect 43168 321836 43220 321842
rect 43168 321778 43220 321784
rect 42984 320612 43036 320618
rect 42984 320554 43036 320560
rect 42156 317484 42208 317490
rect 42156 317426 42208 317432
rect 42800 317484 42852 317490
rect 42800 317426 42852 317432
rect 42168 317045 42196 317426
rect 41970 316976 42026 316985
rect 41970 316911 42026 316920
rect 41984 316404 42012 316911
rect 42154 316024 42210 316033
rect 42154 315959 42210 315968
rect 42168 315757 42196 315959
rect 42154 315480 42210 315489
rect 42154 315415 42210 315424
rect 42168 315180 42196 315415
rect 42154 313848 42210 313857
rect 42154 313783 42210 313792
rect 42168 313344 42196 313783
rect 41786 313168 41842 313177
rect 41786 313103 41842 313112
rect 41800 312732 41828 313103
rect 41786 312352 41842 312361
rect 41786 312287 41842 312296
rect 41800 312052 41828 312287
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41512 301640 41564 301646
rect 41510 301608 41512 301617
rect 41564 301608 41566 301617
rect 41510 301543 41566 301552
rect 41788 300960 41840 300966
rect 41786 300928 41788 300937
rect 41840 300928 41842 300937
rect 41786 300863 41842 300872
rect 43272 299305 43300 342071
rect 44270 341728 44326 341737
rect 44270 341663 44326 341672
rect 44178 340912 44234 340921
rect 44178 340847 44234 340856
rect 43352 329860 43404 329866
rect 43352 329802 43404 329808
rect 43364 321094 43392 329802
rect 43352 321088 43404 321094
rect 43352 321030 43404 321036
rect 43258 299296 43314 299305
rect 43258 299231 43314 299240
rect 43534 298888 43590 298897
rect 43534 298823 43590 298832
rect 32770 296848 32826 296857
rect 32770 296783 32826 296792
rect 32586 296032 32642 296041
rect 32586 295967 32642 295976
rect 32600 285705 32628 295967
rect 32678 294808 32734 294817
rect 32678 294743 32734 294752
rect 32586 285696 32642 285705
rect 32692 285666 32720 294743
rect 32784 285841 32812 296783
rect 35806 296440 35862 296449
rect 35806 296375 35862 296384
rect 32862 295216 32918 295225
rect 32862 295151 32918 295160
rect 32770 285832 32826 285841
rect 32876 285802 32904 295151
rect 33046 294400 33102 294409
rect 33046 294335 33102 294344
rect 32954 293992 33010 294001
rect 32954 293927 33010 293936
rect 32770 285767 32826 285776
rect 32864 285796 32916 285802
rect 32864 285738 32916 285744
rect 32968 285734 32996 293927
rect 33060 285977 33088 294335
rect 35820 287026 35848 296375
rect 42890 293584 42946 293593
rect 42890 293519 42946 293528
rect 35808 287020 35860 287026
rect 35808 286962 35860 286968
rect 42708 287020 42760 287026
rect 42708 286962 42760 286968
rect 33046 285968 33102 285977
rect 33046 285903 33102 285912
rect 32956 285728 33008 285734
rect 32956 285670 33008 285676
rect 32586 285631 32642 285640
rect 32680 285660 32732 285666
rect 32680 285602 32732 285608
rect 41880 285660 41932 285666
rect 41880 285602 41932 285608
rect 41892 283830 41920 285602
rect 41880 283824 41932 283830
rect 41880 283766 41932 283772
rect 41880 283620 41932 283626
rect 41880 283562 41932 283568
rect 41892 283045 41920 283562
rect 42720 281790 42748 286962
rect 42800 285796 42852 285802
rect 42800 285738 42852 285744
rect 42156 281784 42208 281790
rect 42156 281726 42208 281732
rect 42708 281784 42760 281790
rect 42708 281726 42760 281732
rect 42168 281180 42196 281726
rect 42156 281104 42208 281110
rect 42156 281046 42208 281052
rect 42168 280568 42196 281046
rect 42156 279880 42208 279886
rect 42156 279822 42208 279828
rect 42168 279344 42196 279822
rect 42064 278656 42116 278662
rect 42064 278598 42116 278604
rect 42076 278188 42104 278598
rect 42156 278044 42208 278050
rect 42156 277986 42208 277992
rect 42168 277508 42196 277986
rect 42156 277432 42208 277438
rect 42156 277374 42208 277380
rect 42168 276896 42196 277374
rect 42812 276758 42840 285738
rect 42064 276752 42116 276758
rect 42064 276694 42116 276700
rect 42800 276752 42852 276758
rect 42800 276694 42852 276700
rect 42076 276352 42104 276694
rect 42156 274304 42208 274310
rect 42156 274246 42208 274252
rect 42168 273836 42196 274246
rect 42904 273766 42932 293519
rect 42982 293176 43038 293185
rect 42982 293111 43038 293120
rect 42996 279886 43024 293111
rect 43166 292768 43222 292777
rect 43166 292703 43222 292712
rect 43074 292360 43130 292369
rect 43074 292295 43130 292304
rect 42984 279880 43036 279886
rect 42984 279822 43036 279828
rect 43088 274310 43116 292295
rect 43180 278050 43208 292703
rect 43350 291544 43406 291553
rect 43350 291479 43406 291488
rect 43260 285728 43312 285734
rect 43260 285670 43312 285676
rect 43168 278044 43220 278050
rect 43168 277986 43220 277992
rect 43076 274304 43128 274310
rect 43076 274246 43128 274252
rect 42064 273760 42116 273766
rect 42064 273702 42116 273708
rect 42892 273760 42944 273766
rect 42892 273702 42944 273708
rect 42076 273224 42104 273702
rect 43272 272950 43300 285670
rect 43364 278662 43392 291479
rect 43352 278656 43404 278662
rect 43352 278598 43404 278604
rect 42156 272944 42208 272950
rect 42156 272886 42208 272892
rect 43260 272944 43312 272950
rect 43260 272886 43312 272892
rect 42168 272544 42196 272886
rect 41970 272368 42026 272377
rect 41970 272303 42026 272312
rect 41984 272000 42012 272303
rect 42154 270464 42210 270473
rect 42154 270399 42210 270408
rect 42168 270164 42196 270399
rect 42154 270056 42210 270065
rect 42154 269991 42210 270000
rect 42168 269521 42196 269991
rect 42154 269240 42210 269249
rect 42154 269175 42210 269184
rect 42168 268872 42196 269175
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 41512 258392 41564 258398
rect 41510 258360 41512 258369
rect 41564 258360 41566 258369
rect 41510 258295 41566 258304
rect 41788 257848 41840 257854
rect 41788 257790 41840 257796
rect 41800 257689 41828 257790
rect 41786 257680 41842 257689
rect 41786 257615 41842 257624
rect 41512 257576 41564 257582
rect 41510 257544 41512 257553
rect 41564 257544 41566 257553
rect 41510 257479 41566 257488
rect 41788 256896 41840 256902
rect 41786 256864 41788 256873
rect 41840 256864 41842 256873
rect 41786 256799 41842 256808
rect 43548 256057 43576 298823
rect 44192 297265 44220 340847
rect 44284 340105 44312 341663
rect 44270 340096 44326 340105
rect 44270 340031 44326 340040
rect 44284 298081 44312 340031
rect 44376 299713 44404 343334
rect 44362 299704 44418 299713
rect 44362 299639 44418 299648
rect 44270 298072 44326 298081
rect 44270 298007 44326 298016
rect 44178 297256 44234 297265
rect 44178 297191 44234 297200
rect 43626 291952 43682 291961
rect 43626 291887 43682 291896
rect 43640 277438 43668 291887
rect 43628 277432 43680 277438
rect 43628 277374 43680 277380
rect 43534 256048 43590 256057
rect 43534 255983 43590 255992
rect 43442 255640 43498 255649
rect 43442 255575 43498 255584
rect 42706 253600 42762 253609
rect 42706 253535 42762 253544
rect 31666 253056 31722 253065
rect 31666 252991 31722 253000
rect 31680 244254 31708 252991
rect 33046 251832 33102 251841
rect 33046 251767 33102 251776
rect 32770 250608 32826 250617
rect 32770 250543 32826 250552
rect 32784 245654 32812 250543
rect 32862 250200 32918 250209
rect 32862 250135 32918 250144
rect 32876 247602 32904 250135
rect 33060 249830 33088 251767
rect 33048 249824 33100 249830
rect 32954 249792 33010 249801
rect 33048 249766 33100 249772
rect 32954 249727 33010 249736
rect 32968 247738 32996 249727
rect 38290 248160 38346 248169
rect 38290 248095 38346 248104
rect 32968 247710 33088 247738
rect 32876 247574 32996 247602
rect 32784 245626 32904 245654
rect 32876 244390 32904 245626
rect 32864 244384 32916 244390
rect 32864 244326 32916 244332
rect 32968 244322 32996 247574
rect 33060 244458 33088 247710
rect 33048 244452 33100 244458
rect 33048 244394 33100 244400
rect 32956 244316 33008 244322
rect 32956 244258 33008 244264
rect 31668 244248 31720 244254
rect 31668 244190 31720 244196
rect 38304 242894 38332 248095
rect 41510 247752 41566 247761
rect 41510 247687 41512 247696
rect 41564 247687 41566 247696
rect 41512 247658 41564 247664
rect 41510 247344 41566 247353
rect 41510 247279 41512 247288
rect 41564 247279 41566 247288
rect 41512 247250 41564 247256
rect 41510 246936 41566 246945
rect 41510 246871 41512 246880
rect 41564 246871 41566 246880
rect 41512 246842 41564 246848
rect 42720 244526 42748 253535
rect 42890 252376 42946 252385
rect 42890 252311 42946 252320
rect 42904 244594 42932 252311
rect 43258 249520 43314 249529
rect 43258 249455 43314 249464
rect 43074 248704 43130 248713
rect 43074 248639 43130 248648
rect 42892 244588 42944 244594
rect 42892 244530 42944 244536
rect 42708 244520 42760 244526
rect 42708 244462 42760 244468
rect 42892 244452 42944 244458
rect 42892 244394 42944 244400
rect 42708 244248 42760 244254
rect 42708 244190 42760 244196
rect 38292 242888 38344 242894
rect 38292 242830 38344 242836
rect 42156 240372 42208 240378
rect 42156 240314 42208 240320
rect 42168 239836 42196 240314
rect 42720 238474 42748 244190
rect 42800 242888 42852 242894
rect 42800 242830 42852 242836
rect 42156 238468 42208 238474
rect 42156 238410 42208 238416
rect 42708 238468 42760 238474
rect 42708 238410 42760 238416
rect 42168 238000 42196 238410
rect 42156 236700 42208 236706
rect 42156 236642 42208 236648
rect 42168 236164 42196 236642
rect 42812 235414 42840 242830
rect 42904 236706 42932 244394
rect 42984 244316 43036 244322
rect 42984 244258 43036 244264
rect 42892 236700 42944 236706
rect 42892 236642 42944 236648
rect 42156 235408 42208 235414
rect 42156 235350 42208 235356
rect 42800 235408 42852 235414
rect 42800 235350 42852 235356
rect 42168 234969 42196 235350
rect 42156 234660 42208 234666
rect 42156 234602 42208 234608
rect 42168 234328 42196 234602
rect 42156 234252 42208 234258
rect 42156 234194 42208 234200
rect 42168 233681 42196 234194
rect 42156 233368 42208 233374
rect 42156 233310 42208 233316
rect 42168 233104 42196 233310
rect 42156 231124 42208 231130
rect 42156 231066 42208 231072
rect 42168 230656 42196 231066
rect 42996 230586 43024 244258
rect 43088 234258 43116 248639
rect 43168 244384 43220 244390
rect 43168 244326 43220 244332
rect 43076 234252 43128 234258
rect 43076 234194 43128 234200
rect 42156 230580 42208 230586
rect 42156 230522 42208 230528
rect 42984 230580 43036 230586
rect 42984 230522 43036 230528
rect 42168 229976 42196 230522
rect 43180 229906 43208 244326
rect 43272 234666 43300 249455
rect 43350 249112 43406 249121
rect 43350 249047 43406 249056
rect 43364 244662 43392 249047
rect 43352 244656 43404 244662
rect 43352 244598 43404 244604
rect 43352 244520 43404 244526
rect 43352 244462 43404 244468
rect 43260 234660 43312 234666
rect 43260 234602 43312 234608
rect 42156 229900 42208 229906
rect 42156 229842 42208 229848
rect 43168 229900 43220 229906
rect 43168 229842 43220 229848
rect 42168 229364 42196 229842
rect 42156 229084 42208 229090
rect 42156 229026 42208 229032
rect 42168 228820 42196 229026
rect 43364 227458 43392 244462
rect 42064 227452 42116 227458
rect 42064 227394 42116 227400
rect 43352 227452 43404 227458
rect 43352 227394 43404 227400
rect 42076 226984 42104 227394
rect 42156 226840 42208 226846
rect 42156 226782 42208 226788
rect 42168 226304 42196 226782
rect 41970 225992 42026 226001
rect 41970 225927 42026 225936
rect 41984 225692 42012 225927
rect 41512 216776 41564 216782
rect 41512 216718 41564 216724
rect 41420 216708 41472 216714
rect 41420 216650 41472 216656
rect 31852 215824 31904 215830
rect 31852 215766 31904 215772
rect 31668 215756 31720 215762
rect 31668 215698 31720 215704
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 31680 204105 31708 215698
rect 31864 204921 31892 215766
rect 41432 214713 41460 216650
rect 41524 215121 41552 216718
rect 41604 216640 41656 216646
rect 41604 216582 41656 216588
rect 41510 215112 41566 215121
rect 41510 215047 41566 215056
rect 41418 214704 41474 214713
rect 41418 214639 41474 214648
rect 41616 214305 41644 216582
rect 41602 214296 41658 214305
rect 41602 214231 41658 214240
rect 41512 213920 41564 213926
rect 41510 213888 41512 213897
rect 41564 213888 41566 213897
rect 41510 213823 41566 213832
rect 43456 213722 43484 255575
rect 43718 251560 43774 251569
rect 43718 251495 43774 251504
rect 43628 249824 43680 249830
rect 43628 249766 43680 249772
rect 43640 244798 43668 249766
rect 43628 244792 43680 244798
rect 43628 244734 43680 244740
rect 43628 244656 43680 244662
rect 43628 244598 43680 244604
rect 43536 244588 43588 244594
rect 43536 244530 43588 244536
rect 43548 229090 43576 244530
rect 43640 231130 43668 244598
rect 43732 240378 43760 251495
rect 43810 251152 43866 251161
rect 43810 251087 43866 251096
rect 43720 240372 43772 240378
rect 43720 240314 43772 240320
rect 43628 231124 43680 231130
rect 43628 231066 43680 231072
rect 43536 229084 43588 229090
rect 43536 229026 43588 229032
rect 43824 226846 43852 251087
rect 43904 244792 43956 244798
rect 43904 244734 43956 244740
rect 43916 233374 43944 244734
rect 43904 233368 43956 233374
rect 43904 233310 43956 233316
rect 43812 226840 43864 226846
rect 43812 226782 43864 226788
rect 41512 213716 41564 213722
rect 41512 213658 41564 213664
rect 43444 213716 43496 213722
rect 43444 213658 43496 213664
rect 41524 213081 41552 213658
rect 41510 213072 41566 213081
rect 41510 213007 41566 213016
rect 45480 211313 45508 987974
rect 45744 987964 45796 987970
rect 45744 987906 45796 987912
rect 45560 987896 45612 987902
rect 45560 987838 45612 987844
rect 45572 213926 45600 987838
rect 45652 985108 45704 985114
rect 45652 985050 45704 985056
rect 45560 213920 45612 213926
rect 45560 213862 45612 213868
rect 45664 212129 45692 985050
rect 45756 254425 45784 987906
rect 48228 987352 48280 987358
rect 48228 987294 48280 987300
rect 46480 985380 46532 985386
rect 46480 985322 46532 985328
rect 45928 985040 45980 985046
rect 45928 984982 45980 984988
rect 45836 984972 45888 984978
rect 45836 984914 45888 984920
rect 45848 256902 45876 984914
rect 45836 256896 45888 256902
rect 45836 256838 45888 256844
rect 45940 255241 45968 984982
rect 46112 984700 46164 984706
rect 46112 984642 46164 984648
rect 46020 984156 46072 984162
rect 46020 984098 46072 984104
rect 46032 941526 46060 984098
rect 46020 941520 46072 941526
rect 46020 941462 46072 941468
rect 46020 932476 46072 932482
rect 46020 932418 46072 932424
rect 45926 255232 45982 255241
rect 45926 255167 45982 255176
rect 45742 254416 45798 254425
rect 45742 254351 45798 254360
rect 45928 247716 45980 247722
rect 45928 247658 45980 247664
rect 45836 247308 45888 247314
rect 45836 247250 45888 247256
rect 45744 246900 45796 246906
rect 45744 246842 45796 246848
rect 45756 219434 45784 246842
rect 45848 219570 45876 247250
rect 45836 219564 45888 219570
rect 45836 219506 45888 219512
rect 45940 219502 45968 247658
rect 46032 220386 46060 932418
rect 46124 298489 46152 984642
rect 46388 984496 46440 984502
rect 46388 984438 46440 984444
rect 46204 984428 46256 984434
rect 46204 984370 46256 984376
rect 46216 340921 46244 984370
rect 46296 806676 46348 806682
rect 46296 806618 46348 806624
rect 46202 340912 46258 340921
rect 46202 340847 46258 340856
rect 46204 333260 46256 333266
rect 46204 333202 46256 333208
rect 46110 298480 46166 298489
rect 46110 298415 46166 298424
rect 46110 291136 46166 291145
rect 46110 291071 46166 291080
rect 46020 220380 46072 220386
rect 46020 220322 46072 220328
rect 46124 219638 46152 291071
rect 46216 219706 46244 333202
rect 46308 220250 46336 806618
rect 46400 340105 46428 984438
rect 46492 641481 46520 985322
rect 46478 641472 46534 641481
rect 46478 641407 46534 641416
rect 46478 600128 46534 600137
rect 46478 600063 46534 600072
rect 46386 340096 46442 340105
rect 46386 340031 46442 340040
rect 46386 290728 46442 290737
rect 46386 290663 46442 290672
rect 46400 230450 46428 290663
rect 46492 278594 46520 600063
rect 46570 598496 46626 598505
rect 46570 598431 46626 598440
rect 46480 278588 46532 278594
rect 46480 278530 46532 278536
rect 46584 278526 46612 598431
rect 46662 419928 46718 419937
rect 46662 419863 46718 419872
rect 46572 278520 46624 278526
rect 46572 278462 46624 278468
rect 46388 230444 46440 230450
rect 46388 230386 46440 230392
rect 46296 220244 46348 220250
rect 46296 220186 46348 220192
rect 46676 219842 46704 419863
rect 46756 376508 46808 376514
rect 46756 376450 46808 376456
rect 46664 219836 46716 219842
rect 46664 219778 46716 219784
rect 46768 219774 46796 376450
rect 48240 297673 48268 987294
rect 62672 986876 62724 986882
rect 62672 986818 62724 986824
rect 62304 986808 62356 986814
rect 62304 986750 62356 986756
rect 48320 984632 48372 984638
rect 48320 984574 48372 984580
rect 48332 300121 48360 984574
rect 48412 984360 48464 984366
rect 48412 984302 48464 984308
rect 48424 345030 48452 984302
rect 62028 984088 62080 984094
rect 62028 984030 62080 984036
rect 58438 976032 58494 976041
rect 58438 975967 58494 975976
rect 58452 972942 58480 975967
rect 58440 972936 58492 972942
rect 58440 972878 58492 972884
rect 57978 962976 58034 962985
rect 57978 962911 58034 962920
rect 57992 960566 58020 962911
rect 48504 960560 48556 960566
rect 48504 960502 48556 960508
rect 57980 960560 58032 960566
rect 57980 960502 58032 960508
rect 48516 942750 48544 960502
rect 58438 949920 58494 949929
rect 58438 949855 58494 949864
rect 58452 949482 58480 949855
rect 58440 949476 58492 949482
rect 58440 949418 58492 949424
rect 49700 943084 49752 943090
rect 49700 943026 49752 943032
rect 48504 942744 48556 942750
rect 48504 942686 48556 942692
rect 49712 938398 49740 943026
rect 49700 938392 49752 938398
rect 49700 938334 49752 938340
rect 58440 938392 58492 938398
rect 58440 938334 58492 938340
rect 58452 937009 58480 938334
rect 58438 937000 58494 937009
rect 58438 936935 58494 936944
rect 58438 923808 58494 923817
rect 58438 923743 58494 923752
rect 58452 921874 58480 923743
rect 48504 921868 48556 921874
rect 48504 921810 48556 921816
rect 58440 921868 58492 921874
rect 58440 921810 58492 921816
rect 48516 800494 48544 921810
rect 58070 910752 58126 910761
rect 58070 910687 58126 910696
rect 58084 908138 58112 910687
rect 53840 908132 53892 908138
rect 53840 908074 53892 908080
rect 58072 908132 58124 908138
rect 58072 908074 58124 908080
rect 51080 883244 51132 883250
rect 51080 883186 51132 883192
rect 50988 869440 51040 869446
rect 50988 869382 51040 869388
rect 48596 858424 48648 858430
rect 48596 858366 48648 858372
rect 48504 800488 48556 800494
rect 48504 800430 48556 800436
rect 48608 773974 48636 858366
rect 48688 844620 48740 844626
rect 48688 844562 48740 844568
rect 48700 774790 48728 844562
rect 48872 778388 48924 778394
rect 48872 778330 48924 778336
rect 48688 774784 48740 774790
rect 48688 774726 48740 774732
rect 48596 773968 48648 773974
rect 48596 773910 48648 773916
rect 48780 767372 48832 767378
rect 48780 767314 48832 767320
rect 48504 763292 48556 763298
rect 48504 763234 48556 763240
rect 48412 345024 48464 345030
rect 48412 344966 48464 344972
rect 48412 336796 48464 336802
rect 48412 336738 48464 336744
rect 48318 300112 48374 300121
rect 48318 300047 48374 300056
rect 48226 297664 48282 297673
rect 48226 297599 48282 297608
rect 46846 290320 46902 290329
rect 46846 290255 46902 290264
rect 46860 230518 46888 290255
rect 48424 258398 48452 336738
rect 48412 258392 48464 258398
rect 48412 258334 48464 258340
rect 46848 230512 46900 230518
rect 46848 230454 46900 230460
rect 48516 220318 48544 763234
rect 48688 739764 48740 739770
rect 48688 739706 48740 739712
rect 48596 720044 48648 720050
rect 48596 719986 48648 719992
rect 48504 220312 48556 220318
rect 48504 220254 48556 220260
rect 48608 220182 48636 719986
rect 48700 688430 48728 739706
rect 48688 688424 48740 688430
rect 48688 688366 48740 688372
rect 48688 677068 48740 677074
rect 48688 677010 48740 677016
rect 48596 220176 48648 220182
rect 48596 220118 48648 220124
rect 48700 220114 48728 677010
rect 48792 670750 48820 767314
rect 48884 731134 48912 778330
rect 51000 760578 51028 869382
rect 51092 817358 51120 883186
rect 51080 817352 51132 817358
rect 51080 817294 51132 817300
rect 53748 817080 53800 817086
rect 53748 817022 53800 817028
rect 51080 805996 51132 806002
rect 51080 805938 51132 805944
rect 50988 760572 51040 760578
rect 50988 760514 51040 760520
rect 48872 731128 48924 731134
rect 48872 731070 48924 731076
rect 51092 730726 51120 805938
rect 51172 792192 51224 792198
rect 51172 792134 51224 792140
rect 51184 731406 51212 792134
rect 51172 731400 51224 731406
rect 51172 731342 51224 731348
rect 51080 730720 51132 730726
rect 51080 730662 51132 730668
rect 51172 725960 51224 725966
rect 51172 725902 51224 725908
rect 50988 714876 51040 714882
rect 50988 714818 51040 714824
rect 48872 673532 48924 673538
rect 48872 673474 48924 673480
rect 48780 670744 48832 670750
rect 48780 670686 48832 670692
rect 48884 644774 48912 673474
rect 48964 662448 49016 662454
rect 48964 662390 49016 662396
rect 48872 644768 48924 644774
rect 48872 644710 48924 644716
rect 48872 634840 48924 634846
rect 48872 634782 48924 634788
rect 48780 633684 48832 633690
rect 48780 633626 48832 633632
rect 48688 220108 48740 220114
rect 48688 220050 48740 220056
rect 48792 219978 48820 633626
rect 48884 601934 48912 634782
rect 48872 601928 48924 601934
rect 48872 601870 48924 601876
rect 48870 590744 48926 590753
rect 48870 590679 48926 590688
rect 48884 220046 48912 590679
rect 48976 585206 49004 662390
rect 51000 629338 51028 714818
rect 51184 687750 51212 725902
rect 53760 716650 53788 817022
rect 53852 816921 53880 908074
rect 58530 897832 58586 897841
rect 58530 897767 58586 897776
rect 58544 897054 58572 897767
rect 53932 897048 53984 897054
rect 53932 896990 53984 896996
rect 58532 897048 58584 897054
rect 58532 896990 58584 896996
rect 53944 817494 53972 896990
rect 58438 884776 58494 884785
rect 58438 884711 58494 884720
rect 58452 883250 58480 884711
rect 58440 883244 58492 883250
rect 58440 883186 58492 883192
rect 58438 871720 58494 871729
rect 58438 871655 58494 871664
rect 58452 869446 58480 871655
rect 58440 869440 58492 869446
rect 58440 869382 58492 869388
rect 58438 858664 58494 858673
rect 58438 858599 58494 858608
rect 58452 858430 58480 858599
rect 58440 858424 58492 858430
rect 58440 858366 58492 858372
rect 58438 845608 58494 845617
rect 58438 845543 58494 845552
rect 58452 844626 58480 845543
rect 58440 844620 58492 844626
rect 58440 844562 58492 844568
rect 57978 832552 58034 832561
rect 57978 832487 58034 832496
rect 57992 830822 58020 832487
rect 54024 830816 54076 830822
rect 54024 830758 54076 830764
rect 57980 830816 58032 830822
rect 57980 830758 58032 830764
rect 53932 817488 53984 817494
rect 53932 817430 53984 817436
rect 53838 816912 53894 816921
rect 53838 816847 53894 816856
rect 54036 774246 54064 830758
rect 59174 819496 59230 819505
rect 59174 819431 59230 819440
rect 59188 817086 59216 819431
rect 59176 817080 59228 817086
rect 59176 817022 59228 817028
rect 58438 806576 58494 806585
rect 58438 806511 58494 806520
rect 58452 806002 58480 806511
rect 58440 805996 58492 806002
rect 58440 805938 58492 805944
rect 58070 793520 58126 793529
rect 58070 793455 58126 793464
rect 58084 792198 58112 793455
rect 58072 792192 58124 792198
rect 58072 792134 58124 792140
rect 58438 780464 58494 780473
rect 58438 780399 58494 780408
rect 58452 778394 58480 780399
rect 58440 778388 58492 778394
rect 58440 778330 58492 778336
rect 54024 774240 54076 774246
rect 54024 774182 54076 774188
rect 58438 767408 58494 767417
rect 58438 767343 58440 767352
rect 58492 767343 58494 767352
rect 58440 767314 58492 767320
rect 58346 754352 58402 754361
rect 58346 754287 58402 754296
rect 58360 753574 58388 754287
rect 53840 753568 53892 753574
rect 53840 753510 53892 753516
rect 58348 753568 58400 753574
rect 58348 753510 58400 753516
rect 53748 716644 53800 716650
rect 53748 716586 53800 716592
rect 53748 701072 53800 701078
rect 53748 701014 53800 701020
rect 51172 687744 51224 687750
rect 51172 687686 51224 687692
rect 51080 687268 51132 687274
rect 51080 687210 51132 687216
rect 51092 645182 51120 687210
rect 51080 645176 51132 645182
rect 51080 645118 51132 645124
rect 53760 644638 53788 701014
rect 53852 687886 53880 753510
rect 58438 741296 58494 741305
rect 58438 741231 58494 741240
rect 58452 739770 58480 741231
rect 58440 739764 58492 739770
rect 58440 739706 58492 739712
rect 58438 728240 58494 728249
rect 58438 728175 58494 728184
rect 58452 725966 58480 728175
rect 58440 725960 58492 725966
rect 58440 725902 58492 725908
rect 58438 715320 58494 715329
rect 58438 715255 58494 715264
rect 58452 714882 58480 715255
rect 58440 714876 58492 714882
rect 58440 714818 58492 714824
rect 58162 702264 58218 702273
rect 58162 702199 58218 702208
rect 58176 701078 58204 702199
rect 58164 701072 58216 701078
rect 58164 701014 58216 701020
rect 58438 689208 58494 689217
rect 58438 689143 58494 689152
rect 53840 687880 53892 687886
rect 53840 687822 53892 687828
rect 58452 687274 58480 689143
rect 58440 687268 58492 687274
rect 58440 687210 58492 687216
rect 58438 676152 58494 676161
rect 58438 676087 58494 676096
rect 58452 673538 58480 676087
rect 58440 673532 58492 673538
rect 58440 673474 58492 673480
rect 58438 663096 58494 663105
rect 58438 663031 58494 663040
rect 58452 662454 58480 663031
rect 58440 662448 58492 662454
rect 58440 662390 58492 662396
rect 59174 650040 59230 650049
rect 59174 649975 59230 649984
rect 59188 648650 59216 649975
rect 53840 648644 53892 648650
rect 53840 648586 53892 648592
rect 59176 648644 59228 648650
rect 59176 648586 59228 648592
rect 53748 644632 53800 644638
rect 53748 644574 53800 644580
rect 50988 629332 51040 629338
rect 50988 629274 51040 629280
rect 51080 623824 51132 623830
rect 51080 623766 51132 623772
rect 50988 610020 51040 610026
rect 50988 609962 51040 609968
rect 48964 585200 49016 585206
rect 48964 585142 49016 585148
rect 48964 582412 49016 582418
rect 48964 582354 49016 582360
rect 48976 558822 49004 582354
rect 48964 558816 49016 558822
rect 48964 558758 49016 558764
rect 49056 557592 49108 557598
rect 49056 557534 49108 557540
rect 48964 547324 49016 547330
rect 48964 547266 49016 547272
rect 48872 220040 48924 220046
rect 48872 219982 48924 219988
rect 48780 219972 48832 219978
rect 48780 219914 48832 219920
rect 48976 219910 49004 547266
rect 49068 410718 49096 557534
rect 51000 541074 51028 609962
rect 51092 601526 51120 623766
rect 51080 601520 51132 601526
rect 51080 601462 51132 601468
rect 53852 600953 53880 648586
rect 58438 637120 58494 637129
rect 58438 637055 58494 637064
rect 58452 634846 58480 637055
rect 58440 634840 58492 634846
rect 58440 634782 58492 634788
rect 58438 624064 58494 624073
rect 58438 623999 58494 624008
rect 58452 623830 58480 623999
rect 58440 623824 58492 623830
rect 58440 623766 58492 623772
rect 58438 611008 58494 611017
rect 58438 610943 58494 610952
rect 58452 610026 58480 610943
rect 58440 610020 58492 610026
rect 58440 609962 58492 609968
rect 53838 600944 53894 600953
rect 53838 600879 53894 600888
rect 59174 597952 59230 597961
rect 59174 597887 59230 597896
rect 59188 596222 59216 597887
rect 53748 596216 53800 596222
rect 53748 596158 53800 596164
rect 59176 596216 59228 596222
rect 59176 596158 59228 596164
rect 53760 558346 53788 596158
rect 58438 584896 58494 584905
rect 58438 584831 58494 584840
rect 58452 582418 58480 584831
rect 58440 582412 58492 582418
rect 58440 582354 58492 582360
rect 58438 571840 58494 571849
rect 58438 571775 58494 571784
rect 57978 558784 58034 558793
rect 57978 558719 58034 558728
rect 53748 558340 53800 558346
rect 53748 558282 53800 558288
rect 57992 557598 58020 558719
rect 58452 558278 58480 571775
rect 58440 558272 58492 558278
rect 58440 558214 58492 558220
rect 57980 557592 58032 557598
rect 57980 557534 58032 557540
rect 59174 545864 59230 545873
rect 59174 545799 59230 545808
rect 59188 543794 59216 545799
rect 53840 543788 53892 543794
rect 53840 543730 53892 543736
rect 59176 543788 59228 543794
rect 59176 543730 59228 543736
rect 50988 541068 51040 541074
rect 50988 541010 51040 541016
rect 51264 518968 51316 518974
rect 51264 518910 51316 518916
rect 50988 505164 51040 505170
rect 50988 505106 51040 505112
rect 49148 491360 49200 491366
rect 49148 491302 49200 491308
rect 49056 410712 49108 410718
rect 49056 410654 49108 410660
rect 49056 400240 49108 400246
rect 49056 400182 49108 400188
rect 49068 281110 49096 400182
rect 49160 387190 49188 491302
rect 49240 414044 49292 414050
rect 49240 413986 49292 413992
rect 49148 387184 49200 387190
rect 49148 387126 49200 387132
rect 49148 375420 49200 375426
rect 49148 375362 49200 375368
rect 49160 301646 49188 375362
rect 49252 344214 49280 413986
rect 51000 366858 51028 505106
rect 51172 480276 51224 480282
rect 51172 480218 51224 480224
rect 51080 438932 51132 438938
rect 51080 438874 51132 438880
rect 50988 366852 51040 366858
rect 50988 366794 51040 366800
rect 50988 347812 51040 347818
rect 50988 347754 51040 347760
rect 49240 344208 49292 344214
rect 49240 344150 49292 344156
rect 49148 301640 49200 301646
rect 49148 301582 49200 301588
rect 49056 281104 49108 281110
rect 49056 281046 49108 281052
rect 51000 257582 51028 347754
rect 51092 343942 51120 438874
rect 51184 388006 51212 480218
rect 51276 430545 51304 518910
rect 53748 452668 53800 452674
rect 53748 452610 53800 452616
rect 51262 430536 51318 430545
rect 51262 430471 51318 430480
rect 51172 388000 51224 388006
rect 51172 387942 51224 387948
rect 51172 361616 51224 361622
rect 51172 361558 51224 361564
rect 51080 343936 51132 343942
rect 51080 343878 51132 343884
rect 51184 300966 51212 361558
rect 53760 320142 53788 452610
rect 53852 430137 53880 543730
rect 59266 532808 59322 532817
rect 59266 532743 59322 532752
rect 58438 519752 58494 519761
rect 58438 519687 58494 519696
rect 58452 518974 58480 519687
rect 58440 518968 58492 518974
rect 58440 518910 58492 518916
rect 58438 506696 58494 506705
rect 58438 506631 58494 506640
rect 58452 505170 58480 506631
rect 58440 505164 58492 505170
rect 58440 505106 58492 505112
rect 57978 493640 58034 493649
rect 57978 493575 58034 493584
rect 57992 491366 58020 493575
rect 57980 491360 58032 491366
rect 57980 491302 58032 491308
rect 58438 480584 58494 480593
rect 58438 480519 58494 480528
rect 58452 480282 58480 480519
rect 58440 480276 58492 480282
rect 58440 480218 58492 480224
rect 58622 467528 58678 467537
rect 58622 467463 58678 467472
rect 58636 466478 58664 467463
rect 54024 466472 54076 466478
rect 54024 466414 54076 466420
rect 58624 466472 58676 466478
rect 58624 466414 58676 466420
rect 53838 430128 53894 430137
rect 53838 430063 53894 430072
rect 53932 427916 53984 427922
rect 53932 427858 53984 427864
rect 53840 389224 53892 389230
rect 53840 389166 53892 389172
rect 53748 320136 53800 320142
rect 53748 320078 53800 320084
rect 51172 300960 51224 300966
rect 51172 300902 51224 300908
rect 53852 300529 53880 389166
rect 53944 344282 53972 427858
rect 54036 387462 54064 466414
rect 59174 454608 59230 454617
rect 59174 454543 59230 454552
rect 59188 452674 59216 454543
rect 59176 452668 59228 452674
rect 59176 452610 59228 452616
rect 58438 441552 58494 441561
rect 58438 441487 58494 441496
rect 58452 438938 58480 441487
rect 58440 438932 58492 438938
rect 58440 438874 58492 438880
rect 59280 430642 59308 532743
rect 59268 430636 59320 430642
rect 59268 430578 59320 430584
rect 57978 428496 58034 428505
rect 57978 428431 58034 428440
rect 57992 427922 58020 428431
rect 57980 427916 58032 427922
rect 57980 427858 58032 427864
rect 58438 415440 58494 415449
rect 58438 415375 58494 415384
rect 58452 414050 58480 415375
rect 58440 414044 58492 414050
rect 58440 413986 58492 413992
rect 58438 402384 58494 402393
rect 58438 402319 58494 402328
rect 58452 400246 58480 402319
rect 58440 400240 58492 400246
rect 58440 400182 58492 400188
rect 57978 389328 58034 389337
rect 57978 389263 58034 389272
rect 57992 389230 58020 389263
rect 57980 389224 58032 389230
rect 57980 389166 58032 389172
rect 54024 387456 54076 387462
rect 54024 387398 54076 387404
rect 62040 383489 62068 984030
rect 62120 984020 62172 984026
rect 62120 983962 62172 983968
rect 62132 386345 62160 983962
rect 62212 983952 62264 983958
rect 62212 983894 62264 983900
rect 62118 386336 62174 386345
rect 62118 386271 62174 386280
rect 62026 383480 62082 383489
rect 62026 383415 62082 383424
rect 62224 383081 62252 983894
rect 62316 939457 62344 986750
rect 62488 986740 62540 986746
rect 62488 986682 62540 986688
rect 62396 983000 62448 983006
rect 62396 982942 62448 982948
rect 62302 939448 62358 939457
rect 62302 939383 62358 939392
rect 62304 819800 62356 819806
rect 62304 819742 62356 819748
rect 62210 383072 62266 383081
rect 62210 383007 62266 383016
rect 58438 376272 58494 376281
rect 58438 376207 58494 376216
rect 58452 375426 58480 376207
rect 58440 375420 58492 375426
rect 58440 375362 58492 375368
rect 58438 363352 58494 363361
rect 58438 363287 58494 363296
rect 58452 361622 58480 363287
rect 58440 361616 58492 361622
rect 58440 361558 58492 361564
rect 58438 350296 58494 350305
rect 58438 350231 58494 350240
rect 58452 347818 58480 350231
rect 58440 347812 58492 347818
rect 58440 347754 58492 347760
rect 53932 344276 53984 344282
rect 53932 344218 53984 344224
rect 58438 337240 58494 337249
rect 58438 337175 58494 337184
rect 58452 336802 58480 337175
rect 58440 336796 58492 336802
rect 58440 336738 58492 336744
rect 58162 324184 58218 324193
rect 58162 324119 58218 324128
rect 58176 323542 58204 324119
rect 53932 323536 53984 323542
rect 53932 323478 53984 323484
rect 58164 323536 58216 323542
rect 58164 323478 58216 323484
rect 53838 300520 53894 300529
rect 53838 300455 53894 300464
rect 52276 259480 52328 259486
rect 52276 259422 52328 259428
rect 50988 257576 51040 257582
rect 50988 257518 51040 257524
rect 52184 251252 52236 251258
rect 52184 251194 52236 251200
rect 52092 242956 52144 242962
rect 52092 242898 52144 242904
rect 48964 219904 49016 219910
rect 48964 219846 49016 219852
rect 46756 219768 46808 219774
rect 46756 219710 46808 219716
rect 46204 219700 46256 219706
rect 46204 219642 46256 219648
rect 46112 219632 46164 219638
rect 46112 219574 46164 219580
rect 45928 219496 45980 219502
rect 45928 219438 45980 219444
rect 45744 219428 45796 219434
rect 45744 219370 45796 219376
rect 46940 218068 46992 218074
rect 46940 218010 46992 218016
rect 46952 212537 46980 218010
rect 48228 215892 48280 215898
rect 48228 215834 48280 215840
rect 46938 212528 46994 212537
rect 46938 212463 46994 212472
rect 45650 212120 45706 212129
rect 45650 212055 45706 212064
rect 45466 211304 45522 211313
rect 45466 211239 45522 211248
rect 32954 209808 33010 209817
rect 32954 209743 33010 209752
rect 31850 204912 31906 204921
rect 31850 204847 31906 204856
rect 31666 204096 31722 204105
rect 31666 204031 31722 204040
rect 32968 200054 32996 209743
rect 33046 208176 33102 208185
rect 33046 208111 33102 208120
rect 33060 200258 33088 208111
rect 42890 206816 42946 206825
rect 42890 206751 42946 206760
rect 42798 205184 42854 205193
rect 42798 205119 42854 205128
rect 33048 200252 33100 200258
rect 33048 200194 33100 200200
rect 41880 200252 41932 200258
rect 41880 200194 41932 200200
rect 32956 200048 33008 200054
rect 32956 199990 33008 199996
rect 41892 197470 41920 200194
rect 42524 200048 42576 200054
rect 42524 199990 42576 199996
rect 41880 197464 41932 197470
rect 41880 197406 41932 197412
rect 41880 197192 41932 197198
rect 41880 197134 41932 197140
rect 41892 196656 41920 197134
rect 42536 195294 42564 199990
rect 42156 195288 42208 195294
rect 42156 195230 42208 195236
rect 42524 195288 42576 195294
rect 42524 195230 42576 195236
rect 42168 194820 42196 195230
rect 42064 193520 42116 193526
rect 42064 193462 42116 193468
rect 42076 192984 42104 193462
rect 42812 192234 42840 205119
rect 42904 193526 42932 206751
rect 43074 206408 43130 206417
rect 43074 206343 43130 206352
rect 42982 205592 43038 205601
rect 42982 205527 43038 205536
rect 42892 193520 42944 193526
rect 42892 193462 42944 193468
rect 42156 192228 42208 192234
rect 42156 192170 42208 192176
rect 42800 192228 42852 192234
rect 42800 192170 42852 192176
rect 42168 191760 42196 192170
rect 42064 191480 42116 191486
rect 42064 191422 42116 191428
rect 42076 191148 42104 191422
rect 42996 191010 43024 205527
rect 43088 191486 43116 206343
rect 48240 204377 48268 215834
rect 48226 204368 48282 204377
rect 48226 204303 48282 204312
rect 43076 191480 43128 191486
rect 43076 191422 43128 191428
rect 42156 191004 42208 191010
rect 42156 190946 42208 190952
rect 42984 191004 43036 191010
rect 42984 190946 43036 190952
rect 42168 190468 42196 190946
rect 42154 190224 42210 190233
rect 42154 190159 42210 190168
rect 42168 189924 42196 190159
rect 41878 187640 41934 187649
rect 41878 187575 41934 187584
rect 41892 187445 41920 187575
rect 41970 187096 42026 187105
rect 41970 187031 42026 187040
rect 41984 186796 42012 187031
rect 42062 186416 42118 186425
rect 42062 186351 42118 186360
rect 42076 186184 42104 186351
rect 42154 185872 42210 185881
rect 42154 185807 42210 185816
rect 42168 185605 42196 185807
rect 42154 184240 42210 184249
rect 42154 184175 42210 184184
rect 42168 183765 42196 184175
rect 41786 183696 41842 183705
rect 41786 183631 41842 183640
rect 41800 183124 41828 183631
rect 41786 182744 41842 182753
rect 41786 182679 41842 182688
rect 41800 182477 41828 182679
rect 52104 47122 52132 242898
rect 52092 47116 52144 47122
rect 52092 47058 52144 47064
rect 52196 42906 52224 251194
rect 52288 47054 52316 259422
rect 53944 257854 53972 323478
rect 62026 316160 62082 316169
rect 62026 316095 62082 316104
rect 59266 311128 59322 311137
rect 59266 311063 59322 311072
rect 53932 257848 53984 257854
rect 53932 257790 53984 257796
rect 58624 227792 58676 227798
rect 58624 227734 58676 227740
rect 53564 227724 53616 227730
rect 53564 227666 53616 227672
rect 52736 221332 52788 221338
rect 52736 221274 52788 221280
rect 52748 217410 52776 221274
rect 53576 217410 53604 227666
rect 55128 224936 55180 224942
rect 55128 224878 55180 224884
rect 56874 224904 56930 224913
rect 54392 222216 54444 222222
rect 54392 222158 54444 222164
rect 54404 217410 54432 222158
rect 55140 217410 55168 224878
rect 56874 224839 56930 224848
rect 56048 222420 56100 222426
rect 56048 222362 56100 222368
rect 56060 217410 56088 222362
rect 56888 217410 56916 224839
rect 57704 221400 57756 221406
rect 57704 221342 57756 221348
rect 57716 217410 57744 221342
rect 58636 217410 58664 227734
rect 59176 221196 59228 221202
rect 59176 221138 59228 221144
rect 59188 217410 59216 221138
rect 52440 217382 52776 217410
rect 53268 217382 53604 217410
rect 54096 217382 54432 217410
rect 54924 217382 55168 217410
rect 55752 217382 56088 217410
rect 56580 217382 56916 217410
rect 57408 217382 57744 217410
rect 58328 217382 58664 217410
rect 59156 217382 59216 217410
rect 59280 216646 59308 311063
rect 59358 298208 59414 298217
rect 59358 298143 59414 298152
rect 59372 216782 59400 298143
rect 59450 285152 59506 285161
rect 59450 285087 59506 285096
rect 59360 216776 59412 216782
rect 59360 216718 59412 216724
rect 59464 216714 59492 285087
rect 62040 278390 62068 316095
rect 62028 278384 62080 278390
rect 62316 278361 62344 819742
rect 62408 596193 62436 982942
rect 62500 938505 62528 986682
rect 62580 985448 62632 985454
rect 62580 985390 62632 985396
rect 62486 938496 62542 938505
rect 62486 938431 62542 938440
rect 62488 817012 62540 817018
rect 62488 816954 62540 816960
rect 62394 596184 62450 596193
rect 62394 596119 62450 596128
rect 62396 430704 62448 430710
rect 62396 430646 62448 430652
rect 62028 278326 62080 278332
rect 62302 278352 62358 278361
rect 62408 278322 62436 430646
rect 62302 278287 62358 278296
rect 62396 278316 62448 278322
rect 62396 278258 62448 278264
rect 62500 278225 62528 816954
rect 62592 684321 62620 985390
rect 62684 943294 62712 986818
rect 62856 985516 62908 985522
rect 62856 985458 62908 985464
rect 62764 982932 62816 982938
rect 62764 982874 62816 982880
rect 62672 943288 62724 943294
rect 62672 943230 62724 943236
rect 62672 814292 62724 814298
rect 62672 814234 62724 814240
rect 62578 684312 62634 684321
rect 62578 684247 62634 684256
rect 62580 643204 62632 643210
rect 62580 643146 62632 643152
rect 62592 278458 62620 643146
rect 62580 278452 62632 278458
rect 62580 278394 62632 278400
rect 62486 278216 62542 278225
rect 62486 278151 62542 278160
rect 62684 278089 62712 814234
rect 62776 684486 62804 982874
rect 62868 814201 62896 985458
rect 73448 983620 73476 989402
rect 89640 983620 89668 990082
rect 92952 989466 92980 1004634
rect 116032 999932 116084 999938
rect 116032 999874 116084 999880
rect 104348 999864 104400 999870
rect 102782 999832 102838 999841
rect 102782 999767 102784 999776
rect 102836 999767 102838 999776
rect 104346 999832 104348 999841
rect 104400 999832 104402 999841
rect 104346 999767 104402 999776
rect 102784 999738 102836 999744
rect 102322 999696 102378 999705
rect 102322 999631 102324 999640
rect 102376 999631 102378 999640
rect 102324 999602 102376 999608
rect 101954 999560 102010 999569
rect 101954 999495 101956 999504
rect 102008 999495 102010 999504
rect 101956 999466 102008 999472
rect 99288 999456 99340 999462
rect 103152 999456 103204 999462
rect 99288 999398 99340 999404
rect 103150 999424 103152 999433
rect 103204 999424 103206 999433
rect 96528 996464 96580 996470
rect 96526 996432 96528 996441
rect 96580 996432 96582 996441
rect 96526 996367 96582 996376
rect 96528 996124 96580 996130
rect 96528 996066 96580 996072
rect 96436 996056 96488 996062
rect 96436 995998 96488 996004
rect 96448 995897 96476 995998
rect 96434 995888 96490 995897
rect 96434 995823 96490 995832
rect 96540 995353 96568 996066
rect 96526 995344 96582 995353
rect 96526 995279 96582 995288
rect 99300 995217 99328 999398
rect 103150 999359 103206 999368
rect 107658 997248 107714 997257
rect 107658 997183 107660 997192
rect 107712 997183 107714 997192
rect 115938 997248 115994 997257
rect 115938 997183 115940 997192
rect 107660 997154 107712 997160
rect 115992 997183 115994 997192
rect 115940 997154 115992 997160
rect 101128 996464 101180 996470
rect 101126 996432 101128 996441
rect 101180 996432 101182 996441
rect 101126 996367 101182 996376
rect 100298 996160 100354 996169
rect 100298 996095 100300 996104
rect 100352 996095 100354 996104
rect 100758 996160 100814 996169
rect 100758 996095 100814 996104
rect 101494 996160 101550 996169
rect 101494 996095 101550 996104
rect 108486 996160 108542 996169
rect 108486 996095 108542 996104
rect 108854 996160 108910 996169
rect 108854 996095 108856 996104
rect 100300 996066 100352 996072
rect 100772 995858 100800 996095
rect 101508 996062 101536 996095
rect 108500 996062 108528 996095
rect 108908 996095 108910 996104
rect 113272 996124 113324 996130
rect 108856 996066 108908 996072
rect 113272 996066 113324 996072
rect 101496 996056 101548 996062
rect 101496 995998 101548 996004
rect 108488 996056 108540 996062
rect 108488 995998 108540 996004
rect 113180 996056 113232 996062
rect 113180 995998 113232 996004
rect 110418 995888 110474 995897
rect 100760 995852 100812 995858
rect 110418 995823 110474 995832
rect 100760 995794 100812 995800
rect 100206 995616 100262 995625
rect 100206 995551 100262 995560
rect 104162 995616 104218 995625
rect 104162 995551 104218 995560
rect 104346 995616 104402 995625
rect 104346 995551 104402 995560
rect 99286 995208 99342 995217
rect 99286 995143 99342 995152
rect 100220 993857 100248 995551
rect 100206 993848 100262 993857
rect 100206 993783 100262 993792
rect 104176 993682 104204 995551
rect 104360 993721 104388 995551
rect 104346 993712 104402 993721
rect 104164 993676 104216 993682
rect 104346 993647 104402 993656
rect 104164 993618 104216 993624
rect 92940 989460 92992 989466
rect 92940 989402 92992 989408
rect 105820 989460 105872 989466
rect 105820 989402 105872 989408
rect 105832 983620 105860 989402
rect 110432 984162 110460 995823
rect 110786 995752 110842 995761
rect 110786 995687 110842 995696
rect 110602 995616 110658 995625
rect 110602 995551 110658 995560
rect 110616 986814 110644 995551
rect 110604 986808 110656 986814
rect 110604 986750 110656 986756
rect 110800 986746 110828 995687
rect 113192 986882 113220 995998
rect 113284 989466 113312 996066
rect 116044 990894 116072 999874
rect 116032 990888 116084 990894
rect 116032 990830 116084 990836
rect 122104 990820 122156 990826
rect 122104 990762 122156 990768
rect 113272 989460 113324 989466
rect 113272 989402 113324 989408
rect 113180 986876 113232 986882
rect 113180 986818 113232 986824
rect 110788 986740 110840 986746
rect 110788 986682 110840 986688
rect 110420 984156 110472 984162
rect 110420 984098 110472 984104
rect 122116 983620 122144 990762
rect 125520 986950 125548 1004634
rect 125612 996062 125640 1005110
rect 125692 1004828 125744 1004834
rect 125692 1004770 125744 1004776
rect 125704 996198 125732 1004770
rect 125692 996192 125744 996198
rect 125692 996134 125744 996140
rect 125796 996130 125824 1005178
rect 144276 999116 144328 999122
rect 144276 999058 144328 999064
rect 143816 997756 143868 997762
rect 143816 997698 143868 997704
rect 125784 996124 125836 996130
rect 125784 996066 125836 996072
rect 125600 996056 125652 996062
rect 125600 995998 125652 996004
rect 136272 995852 136324 995858
rect 136272 995794 136324 995800
rect 136824 995852 136876 995858
rect 136824 995794 136876 995800
rect 137928 995852 137980 995858
rect 137928 995794 137980 995800
rect 136284 995738 136312 995794
rect 136836 995738 136864 995794
rect 137940 995738 137968 995794
rect 139216 995784 139268 995790
rect 135930 995710 136312 995738
rect 136482 995710 136864 995738
rect 137770 995710 137968 995738
rect 138966 995732 139216 995738
rect 142802 995752 142858 995761
rect 138966 995726 139268 995732
rect 138966 995710 139256 995726
rect 142646 995710 142802 995738
rect 142802 995687 142858 995696
rect 133144 995648 133196 995654
rect 132158 995586 132448 995602
rect 132802 995596 133144 995602
rect 137374 995616 137430 995625
rect 132802 995590 133196 995596
rect 132158 995580 132460 995586
rect 132158 995574 132408 995580
rect 132802 995574 133184 995590
rect 137126 995574 137374 995602
rect 137374 995551 137430 995560
rect 132408 995522 132460 995528
rect 143828 995518 143856 997698
rect 144288 997257 144316 999058
rect 144274 997248 144330 997257
rect 144274 997183 144330 997192
rect 130016 995512 130068 995518
rect 129766 995460 130016 995466
rect 143816 995512 143868 995518
rect 133694 995480 133750 995489
rect 129766 995454 130068 995460
rect 128464 993682 128492 995452
rect 129108 993750 129136 995452
rect 129766 995438 130056 995454
rect 131606 995450 131896 995466
rect 131606 995444 131908 995450
rect 131606 995438 131856 995444
rect 133446 995438 133694 995466
rect 141054 995480 141110 995489
rect 140162 995438 140544 995466
rect 140806 995438 141054 995466
rect 133694 995415 133750 995424
rect 131856 995386 131908 995392
rect 140516 993750 140544 995438
rect 143816 995454 143868 995460
rect 141054 995415 141110 995424
rect 129096 993744 129148 993750
rect 129096 993686 129148 993692
rect 140504 993744 140556 993750
rect 140504 993686 140556 993692
rect 128452 993676 128504 993682
rect 128452 993618 128504 993624
rect 144840 988786 144868 1005382
rect 160282 1005343 160338 1005352
rect 209226 1005408 209282 1005417
rect 356518 1005408 356520 1005417
rect 356572 1005408 356574 1005417
rect 209226 1005343 209228 1005352
rect 209280 1005343 209282 1005352
rect 227720 1005372 227772 1005378
rect 209228 1005314 209280 1005320
rect 227720 1005314 227772 1005320
rect 253296 1005372 253348 1005378
rect 253296 1005314 253348 1005320
rect 280068 1005372 280120 1005378
rect 356518 1005343 356574 1005352
rect 361026 1005408 361082 1005417
rect 361026 1005343 361028 1005352
rect 280068 1005314 280120 1005320
rect 361080 1005343 361082 1005352
rect 361028 1005314 361080 1005320
rect 195336 1005168 195388 1005174
rect 209596 1005168 209648 1005174
rect 195336 1005110 195388 1005116
rect 201498 1005136 201554 1005145
rect 150900 1005032 150952 1005038
rect 150898 1005000 150900 1005009
rect 175188 1005032 175240 1005038
rect 150952 1005000 150954 1005009
rect 150898 1004935 150954 1004944
rect 157798 1005000 157854 1005009
rect 175188 1004974 175240 1004980
rect 157798 1004935 157800 1004944
rect 157852 1004935 157854 1004944
rect 174084 1004964 174136 1004970
rect 157800 1004906 157852 1004912
rect 174084 1004906 174136 1004912
rect 156970 1004864 157026 1004873
rect 156970 1004799 156972 1004808
rect 157024 1004799 157026 1004808
rect 173992 1004828 174044 1004834
rect 156972 1004770 157024 1004776
rect 173992 1004770 174044 1004776
rect 154488 1004760 154540 1004766
rect 149702 1004728 149758 1004737
rect 146024 1004692 146076 1004698
rect 150070 1004728 150126 1004737
rect 149758 1004686 150070 1004714
rect 149702 1004663 149758 1004672
rect 159456 1004760 159508 1004766
rect 154488 1004702 154540 1004708
rect 154946 1004728 155002 1004737
rect 150070 1004663 150126 1004672
rect 146024 1004634 146076 1004640
rect 146036 995450 146064 1004634
rect 148876 996464 148928 996470
rect 148874 996432 148876 996441
rect 154120 996464 154172 996470
rect 148928 996432 148930 996441
rect 146208 996396 146260 996402
rect 148874 996367 148930 996376
rect 151726 996432 151782 996441
rect 151726 996367 151728 996376
rect 146208 996338 146260 996344
rect 151780 996367 151782 996376
rect 154118 996432 154120 996441
rect 154172 996432 154174 996441
rect 154118 996367 154174 996376
rect 151728 996338 151780 996344
rect 146116 996260 146168 996266
rect 146116 996202 146168 996208
rect 146024 995444 146076 995450
rect 146024 995386 146076 995392
rect 146128 993818 146156 996202
rect 146220 995353 146248 996338
rect 153750 996296 153806 996305
rect 153750 996231 153752 996240
rect 153804 996231 153806 996240
rect 153752 996202 153804 996208
rect 150898 996160 150954 996169
rect 150898 996095 150954 996104
rect 151266 996160 151322 996169
rect 151266 996095 151322 996104
rect 152554 996160 152610 996169
rect 152554 996095 152610 996104
rect 152922 996160 152978 996169
rect 152922 996095 152978 996104
rect 153382 996160 153438 996169
rect 153382 996095 153438 996104
rect 150912 995858 150940 996095
rect 151280 995926 151308 996095
rect 151268 995920 151320 995926
rect 151268 995862 151320 995868
rect 150900 995852 150952 995858
rect 150900 995794 150952 995800
rect 152568 995790 152596 996095
rect 152556 995784 152608 995790
rect 152556 995726 152608 995732
rect 152936 995654 152964 996095
rect 152924 995648 152976 995654
rect 152924 995590 152976 995596
rect 153396 995586 153424 996095
rect 153384 995580 153436 995586
rect 153384 995522 153436 995528
rect 146206 995344 146262 995353
rect 146206 995279 146262 995288
rect 146116 993812 146168 993818
rect 146116 993754 146168 993760
rect 151820 993744 151872 993750
rect 151820 993686 151872 993692
rect 151832 989466 151860 993686
rect 151820 989460 151872 989466
rect 151820 989402 151872 989408
rect 138296 988780 138348 988786
rect 138296 988722 138348 988728
rect 144828 988780 144880 988786
rect 144828 988722 144880 988728
rect 125508 986944 125560 986950
rect 125508 986886 125560 986892
rect 138308 983620 138336 988722
rect 154500 983620 154528 1004702
rect 154946 1004663 154948 1004672
rect 155000 1004663 155002 1004672
rect 159454 1004728 159456 1004737
rect 173900 1004760 173952 1004766
rect 159508 1004728 159510 1004737
rect 159454 1004663 159510 1004672
rect 160650 1004728 160706 1004737
rect 173900 1004702 173952 1004708
rect 160650 1004663 160652 1004672
rect 154948 1004634 155000 1004640
rect 160704 1004663 160706 1004672
rect 160652 1004634 160704 1004640
rect 155776 999592 155828 999598
rect 155774 999560 155776 999569
rect 160284 999592 160336 999598
rect 155828 999560 155830 999569
rect 155774 999495 155830 999504
rect 159086 999560 159142 999569
rect 160284 999534 160336 999540
rect 159086 999495 159088 999504
rect 159140 999495 159142 999504
rect 159088 999466 159140 999472
rect 158258 999152 158314 999161
rect 158258 999087 158260 999096
rect 158312 999087 158314 999096
rect 158260 999058 158312 999064
rect 156142 997792 156198 997801
rect 156142 997727 156144 997736
rect 156196 997727 156198 997736
rect 156144 997698 156196 997704
rect 159456 996192 159508 996198
rect 154578 996160 154634 996169
rect 154578 996095 154634 996104
rect 156970 996160 157026 996169
rect 156970 996095 157026 996104
rect 157798 996160 157854 996169
rect 157798 996095 157800 996104
rect 154592 995994 154620 996095
rect 156984 996062 157012 996095
rect 157852 996095 157854 996104
rect 159454 996160 159456 996169
rect 159508 996160 159510 996169
rect 159454 996095 159510 996104
rect 157800 996066 157852 996072
rect 156972 996056 157024 996062
rect 156972 995998 157024 996004
rect 160192 996056 160244 996062
rect 160192 995998 160244 996004
rect 154580 995988 154632 995994
rect 154580 995930 154632 995936
rect 160204 984162 160232 995998
rect 160296 993682 160324 999534
rect 162860 999524 162912 999530
rect 162860 999466 162912 999472
rect 162872 997121 162900 999466
rect 162858 997112 162914 997121
rect 162858 997047 162914 997056
rect 173912 996198 173940 1004702
rect 173900 996192 173952 996198
rect 173900 996134 173952 996140
rect 174004 996130 174032 1004770
rect 173992 996124 174044 996130
rect 173992 996066 174044 996072
rect 174096 996062 174124 1004906
rect 174084 996056 174136 996062
rect 174084 995998 174136 996004
rect 168378 995888 168434 995897
rect 168378 995823 168434 995832
rect 162950 995752 163006 995761
rect 162950 995687 163006 995696
rect 162858 995616 162914 995625
rect 162858 995551 162914 995560
rect 160284 993676 160336 993682
rect 160284 993618 160336 993624
rect 162872 984298 162900 995551
rect 162860 984292 162912 984298
rect 162860 984234 162912 984240
rect 162964 984230 162992 995687
rect 168392 990690 168420 995823
rect 168380 990684 168432 990690
rect 168380 990626 168432 990632
rect 170404 990684 170456 990690
rect 170404 990626 170456 990632
rect 162952 984224 163004 984230
rect 162952 984166 163004 984172
rect 160192 984156 160244 984162
rect 160192 984098 160244 984104
rect 170416 983634 170444 990626
rect 175200 987018 175228 1004974
rect 195152 1004624 195204 1004630
rect 195152 1004566 195204 1004572
rect 195164 997257 195192 1004566
rect 195244 999660 195296 999666
rect 195244 999602 195296 999608
rect 195150 997248 195206 997257
rect 195150 997183 195206 997192
rect 188160 995852 188212 995858
rect 188160 995794 188212 995800
rect 184480 995784 184532 995790
rect 184184 995732 184480 995738
rect 187606 995752 187662 995761
rect 184184 995726 184532 995732
rect 184184 995710 184520 995726
rect 187312 995710 187606 995738
rect 188172 995738 188200 995794
rect 195256 995790 195284 999602
rect 195348 997121 195376 1005110
rect 201498 1005071 201500 1005080
rect 201552 1005071 201554 1005080
rect 202326 1005136 202382 1005145
rect 202326 1005071 202328 1005080
rect 201500 1005042 201552 1005048
rect 202380 1005071 202382 1005080
rect 209594 1005136 209596 1005145
rect 210884 1005168 210936 1005174
rect 209648 1005136 209650 1005145
rect 209594 1005071 209650 1005080
rect 210882 1005136 210884 1005145
rect 210936 1005136 210938 1005145
rect 210882 1005071 210938 1005080
rect 227628 1005100 227680 1005106
rect 202328 1005042 202380 1005048
rect 227628 1005042 227680 1005048
rect 208398 1005000 208454 1005009
rect 208398 1004935 208400 1004944
rect 208452 1004935 208454 1004944
rect 208400 1004906 208452 1004912
rect 195980 1004760 196032 1004766
rect 206376 1004760 206428 1004766
rect 195980 1004702 196032 1004708
rect 205178 1004728 205234 1004737
rect 195704 1004692 195756 1004698
rect 195704 1004634 195756 1004640
rect 195612 999592 195664 999598
rect 195612 999534 195664 999540
rect 195428 999524 195480 999530
rect 195428 999466 195480 999472
rect 195334 997112 195390 997121
rect 195334 997047 195390 997056
rect 194324 995784 194376 995790
rect 187864 995710 188200 995738
rect 190348 995722 190684 995738
rect 194028 995732 194324 995738
rect 194028 995726 194376 995732
rect 195244 995784 195296 995790
rect 195244 995726 195296 995732
rect 190348 995716 190696 995722
rect 190348 995710 190644 995716
rect 187606 995687 187662 995696
rect 194028 995710 194364 995726
rect 195440 995722 195468 999466
rect 195520 999456 195572 999462
rect 195520 999398 195572 999404
rect 195428 995716 195480 995722
rect 190644 995658 190696 995664
rect 195428 995658 195480 995664
rect 195532 995654 195560 999398
rect 189448 995648 189500 995654
rect 184676 995586 184828 995602
rect 184664 995580 184828 995586
rect 184716 995574 184828 995580
rect 189152 995596 189448 995602
rect 195520 995648 195572 995654
rect 192482 995616 192538 995625
rect 189152 995590 189500 995596
rect 189152 995574 189488 995590
rect 192188 995574 192482 995602
rect 195520 995590 195572 995596
rect 192482 995551 192538 995560
rect 184664 995522 184716 995528
rect 195624 995518 195652 999534
rect 188804 995512 188856 995518
rect 179860 995438 180196 995466
rect 180168 993750 180196 995438
rect 180490 995314 180518 995452
rect 181148 995438 181484 995466
rect 182988 995438 183324 995466
rect 183540 995450 183876 995466
rect 188508 995460 188804 995466
rect 195612 995512 195664 995518
rect 188508 995454 188856 995460
rect 183540 995444 183888 995450
rect 183540 995438 183836 995444
rect 180478 995308 180530 995314
rect 180478 995250 180530 995256
rect 180156 993744 180208 993750
rect 180156 993686 180208 993692
rect 181456 993682 181484 995438
rect 183296 995382 183324 995438
rect 188508 995438 188844 995454
rect 191544 995438 191880 995466
rect 195612 995454 195664 995460
rect 183836 995386 183888 995392
rect 183284 995376 183336 995382
rect 183284 995318 183336 995324
rect 191852 993721 191880 995438
rect 195716 995314 195744 1004634
rect 195992 995382 196020 1004702
rect 205178 1004663 205180 1004672
rect 205232 1004663 205234 1004672
rect 205914 1004728 205970 1004737
rect 205914 1004663 205970 1004672
rect 206374 1004728 206376 1004737
rect 206428 1004728 206430 1004737
rect 206374 1004663 206430 1004672
rect 218058 1004728 218114 1004737
rect 218058 1004663 218114 1004672
rect 205180 1004634 205232 1004640
rect 205928 1004630 205956 1004663
rect 205916 1004624 205968 1004630
rect 205916 1004566 205968 1004572
rect 205546 999696 205602 999705
rect 205546 999631 205548 999640
rect 205600 999631 205602 999640
rect 205548 999602 205600 999608
rect 203524 999592 203576 999598
rect 203522 999560 203524 999569
rect 203576 999560 203578 999569
rect 203522 999495 203578 999504
rect 203890 999560 203946 999569
rect 203890 999495 203892 999504
rect 203944 999495 203946 999504
rect 203892 999466 203944 999472
rect 202328 999456 202380 999462
rect 202326 999424 202328 999433
rect 202380 999424 202382 999433
rect 198372 999388 198424 999394
rect 202326 999359 202382 999368
rect 204718 999424 204774 999433
rect 204718 999359 204720 999368
rect 198372 999330 198424 999336
rect 204772 999359 204774 999368
rect 204720 999330 204772 999336
rect 198384 995450 198412 999330
rect 198464 999320 198516 999326
rect 204352 999320 204404 999326
rect 198464 999262 198516 999268
rect 202694 999288 202750 999297
rect 198476 995926 198504 999262
rect 198648 999252 198700 999258
rect 202694 999223 202696 999232
rect 198648 999194 198700 999200
rect 202748 999223 202750 999232
rect 204350 999288 204352 999297
rect 204404 999288 204406 999297
rect 204350 999223 204406 999232
rect 202696 999194 202748 999200
rect 198556 999184 198608 999190
rect 198556 999126 198608 999132
rect 198464 995920 198516 995926
rect 198464 995862 198516 995868
rect 198568 995586 198596 999126
rect 198660 995858 198688 999194
rect 203064 999184 203116 999190
rect 203062 999152 203064 999161
rect 203116 999152 203118 999161
rect 218072 999134 218100 1004663
rect 218072 999106 219112 999134
rect 203062 999087 203118 999096
rect 210422 997248 210478 997257
rect 210422 997183 210424 997192
rect 210476 997183 210478 997192
rect 215298 997248 215354 997257
rect 215298 997183 215300 997192
rect 210424 997154 210476 997160
rect 215352 997183 215354 997192
rect 215300 997154 215352 997160
rect 211252 996260 211304 996266
rect 211252 996202 211304 996208
rect 208768 996192 208820 996198
rect 208766 996160 208768 996169
rect 211264 996169 211292 996202
rect 212816 996192 212868 996198
rect 208820 996160 208822 996169
rect 204168 996124 204220 996130
rect 208766 996095 208822 996104
rect 209594 996160 209650 996169
rect 209594 996095 209650 996104
rect 211250 996160 211306 996169
rect 211250 996095 211306 996104
rect 211618 996160 211674 996169
rect 212816 996134 212868 996140
rect 211618 996095 211620 996104
rect 204168 996066 204220 996072
rect 198648 995852 198700 995858
rect 198648 995794 198700 995800
rect 198556 995580 198608 995586
rect 198556 995522 198608 995528
rect 198372 995444 198424 995450
rect 198372 995386 198424 995392
rect 195980 995376 196032 995382
rect 195980 995318 196032 995324
rect 195704 995308 195756 995314
rect 195704 995250 195756 995256
rect 191838 993712 191894 993721
rect 181444 993676 181496 993682
rect 191838 993647 191894 993656
rect 181444 993618 181496 993624
rect 204180 990690 204208 996066
rect 209608 996062 209636 996095
rect 209596 996056 209648 996062
rect 209596 995998 209648 996004
rect 211264 995994 211292 996095
rect 211672 996095 211674 996104
rect 211620 996066 211672 996072
rect 212632 996056 212684 996062
rect 212632 995998 212684 996004
rect 211252 995988 211304 995994
rect 211252 995930 211304 995936
rect 207018 995888 207074 995897
rect 207018 995823 207074 995832
rect 207032 993750 207060 995823
rect 207754 995616 207810 995625
rect 207754 995551 207810 995560
rect 207020 993744 207072 993750
rect 207020 993686 207072 993692
rect 207768 993682 207796 995551
rect 207756 993676 207808 993682
rect 207756 993618 207808 993624
rect 203156 990684 203208 990690
rect 203156 990626 203208 990632
rect 204168 990684 204220 990690
rect 204168 990626 204220 990632
rect 186964 989460 187016 989466
rect 186964 989402 187016 989408
rect 175188 987012 175240 987018
rect 175188 986954 175240 986960
rect 170416 983606 170798 983634
rect 186976 983620 187004 989402
rect 203168 983620 203196 990626
rect 212644 984570 212672 995998
rect 212828 987086 212856 996134
rect 215484 995988 215536 995994
rect 215484 995930 215536 995936
rect 215496 987154 215524 995930
rect 216586 995888 216642 995897
rect 216586 995823 216642 995832
rect 216600 989466 216628 995823
rect 216588 989460 216640 989466
rect 216588 989402 216640 989408
rect 215484 987148 215536 987154
rect 215484 987090 215536 987096
rect 212816 987080 212868 987086
rect 212816 987022 212868 987028
rect 212632 984564 212684 984570
rect 212632 984506 212684 984512
rect 219084 983634 219112 999106
rect 227640 987222 227668 1005042
rect 227732 996062 227760 1005314
rect 227904 1005168 227956 1005174
rect 227904 1005110 227956 1005116
rect 227812 1004964 227864 1004970
rect 227812 1004906 227864 1004912
rect 227824 996130 227852 1004906
rect 227916 996198 227944 1005110
rect 253308 1005038 253336 1005314
rect 259828 1005304 259880 1005310
rect 259826 1005272 259828 1005281
rect 259880 1005272 259882 1005281
rect 259826 1005207 259882 1005216
rect 260194 1005272 260250 1005281
rect 260194 1005207 260196 1005216
rect 260248 1005207 260250 1005216
rect 265072 1005236 265124 1005242
rect 260196 1005178 260248 1005184
rect 265072 1005178 265124 1005184
rect 263048 1005168 263100 1005174
rect 261022 1005136 261078 1005145
rect 261022 1005071 261024 1005080
rect 261076 1005071 261078 1005080
rect 263046 1005136 263048 1005145
rect 264336 1005168 264388 1005174
rect 263100 1005136 263102 1005145
rect 263046 1005071 263102 1005080
rect 264334 1005136 264336 1005145
rect 264388 1005136 264390 1005145
rect 264334 1005071 264390 1005080
rect 261024 1005042 261076 1005048
rect 252836 1005032 252888 1005038
rect 252834 1005000 252836 1005009
rect 253296 1005032 253348 1005038
rect 252888 1005000 252890 1005009
rect 252834 1004935 252890 1004944
rect 253294 1005000 253296 1005009
rect 260656 1005032 260708 1005038
rect 253348 1005000 253350 1005009
rect 253294 1004935 253350 1004944
rect 260654 1005000 260656 1005009
rect 260708 1005000 260710 1005009
rect 260654 1004935 260710 1004944
rect 262678 1005000 262734 1005009
rect 262678 1004935 262680 1004944
rect 262732 1004935 262734 1004944
rect 264334 1005000 264390 1005009
rect 264334 1004935 264336 1004944
rect 262680 1004906 262732 1004912
rect 264388 1004935 264390 1004944
rect 264336 1004906 264388 1004912
rect 261852 1004896 261904 1004902
rect 261850 1004864 261852 1004873
rect 261904 1004864 261906 1004873
rect 261850 1004799 261906 1004808
rect 262220 1004760 262272 1004766
rect 252466 1004728 252522 1004737
rect 252834 1004728 252890 1004737
rect 252522 1004686 252834 1004714
rect 252466 1004663 252522 1004672
rect 252834 1004663 252890 1004672
rect 261482 1004728 261538 1004737
rect 261482 1004663 261484 1004672
rect 261536 1004663 261538 1004672
rect 262218 1004728 262220 1004737
rect 262272 1004728 262274 1004737
rect 262218 1004663 262274 1004672
rect 263506 1004728 263562 1004737
rect 263874 1004728 263930 1004737
rect 263562 1004686 263874 1004714
rect 263506 1004663 263562 1004672
rect 263874 1004663 263930 1004672
rect 261484 1004634 261536 1004640
rect 258630 999968 258686 999977
rect 246764 999932 246816 999938
rect 258630 999903 258632 999912
rect 246764 999874 246816 999880
rect 258684 999903 258686 999912
rect 258632 999874 258684 999880
rect 246580 999864 246632 999870
rect 246580 999806 246632 999812
rect 246592 999274 246620 999806
rect 246672 999796 246724 999802
rect 246672 999738 246724 999744
rect 246500 999246 246620 999274
rect 227904 996192 227956 996198
rect 227904 996134 227956 996140
rect 227812 996124 227864 996130
rect 227812 996066 227864 996072
rect 227720 996056 227772 996062
rect 227720 995998 227772 996004
rect 246500 995926 246528 999246
rect 246580 999116 246632 999122
rect 246580 999058 246632 999064
rect 246592 997257 246620 999058
rect 246578 997248 246634 997257
rect 246578 997183 246634 997192
rect 246488 995920 246540 995926
rect 246488 995862 246540 995868
rect 239036 995852 239088 995858
rect 239036 995794 239088 995800
rect 239588 995852 239640 995858
rect 239588 995794 239640 995800
rect 234526 995752 234582 995761
rect 234416 995710 234526 995738
rect 239048 995738 239076 995794
rect 239600 995738 239628 995794
rect 246684 995790 246712 999738
rect 245568 995784 245620 995790
rect 240046 995752 240102 995761
rect 238740 995710 239076 995738
rect 239292 995710 239628 995738
rect 239936 995710 240046 995738
rect 234526 995687 234582 995696
rect 243616 995722 243952 995738
rect 245456 995732 245568 995738
rect 245456 995726 245620 995732
rect 246672 995784 246724 995790
rect 246672 995726 246724 995732
rect 243616 995716 243964 995722
rect 243616 995710 243912 995716
rect 240046 995687 240102 995696
rect 245456 995710 245608 995726
rect 246776 995722 246804 999874
rect 257344 999864 257396 999870
rect 256974 999832 257030 999841
rect 256974 999767 256976 999776
rect 257028 999767 257030 999776
rect 257342 999832 257344 999841
rect 257396 999832 257398 999841
rect 257342 999767 257398 999776
rect 256976 999738 257028 999744
rect 246948 999728 247000 999734
rect 257804 999728 257856 999734
rect 246948 999670 247000 999676
rect 257802 999696 257804 999705
rect 257856 999696 257858 999705
rect 246960 996033 246988 999670
rect 257802 999631 257858 999640
rect 256514 999288 256570 999297
rect 253848 999252 253900 999258
rect 256514 999223 256516 999232
rect 253848 999194 253900 999200
rect 256568 999223 256570 999232
rect 256516 999194 256568 999200
rect 253662 996160 253718 996169
rect 253662 996095 253718 996104
rect 246946 996024 247002 996033
rect 246946 995959 247002 995968
rect 246764 995716 246816 995722
rect 243912 995658 243964 995664
rect 246764 995658 246816 995664
rect 253676 995654 253704 996095
rect 240876 995648 240928 995654
rect 240580 995596 240876 995602
rect 253664 995648 253716 995654
rect 242070 995616 242126 995625
rect 240580 995590 240928 995596
rect 240580 995574 240916 995590
rect 241776 995574 242070 995602
rect 253664 995590 253716 995596
rect 242070 995551 242126 995560
rect 235906 995480 235962 995489
rect 231288 995438 231624 995466
rect 231932 995438 232268 995466
rect 232576 995438 232912 995466
rect 231596 993682 231624 995438
rect 232240 994129 232268 995438
rect 232226 994120 232282 994129
rect 232226 994055 232282 994064
rect 232884 993993 232912 995438
rect 234954 995217 234982 995452
rect 235612 995438 235906 995466
rect 235906 995415 235962 995424
rect 236242 995353 236270 995452
rect 242972 995438 243308 995466
rect 236228 995344 236284 995353
rect 236228 995279 236284 995288
rect 234940 995208 234996 995217
rect 234940 995143 234996 995152
rect 232870 993984 232926 993993
rect 232870 993919 232926 993928
rect 243280 993857 243308 995438
rect 253860 994129 253888 999194
rect 258540 999184 258592 999190
rect 258538 999152 258540 999161
rect 262220 999184 262272 999190
rect 258592 999152 258594 999161
rect 262220 999126 262272 999132
rect 258538 999087 258594 999096
rect 254122 996160 254178 996169
rect 254122 996095 254178 996104
rect 254490 996160 254546 996169
rect 254490 996095 254546 996104
rect 254136 995858 254164 996095
rect 254124 995852 254176 995858
rect 254124 995794 254176 995800
rect 254504 995353 254532 996095
rect 254490 995344 254546 995353
rect 254490 995279 254546 995288
rect 253846 994120 253902 994129
rect 253846 994055 253902 994064
rect 243266 993848 243322 993857
rect 243266 993783 243322 993792
rect 248326 993712 248382 993721
rect 231584 993676 231636 993682
rect 262232 993682 262260 999126
rect 265084 996130 265112 1005178
rect 269210 1005136 269266 1005145
rect 265256 1005100 265308 1005106
rect 269210 1005071 269266 1005080
rect 265256 1005042 265308 1005048
rect 265164 1004692 265216 1004698
rect 265164 1004634 265216 1004640
rect 265176 999122 265204 1004634
rect 265164 999116 265216 999122
rect 265164 999058 265216 999064
rect 265072 996124 265124 996130
rect 265072 996066 265124 996072
rect 265268 996062 265296 1005042
rect 267830 1005000 267886 1005009
rect 267830 1004935 267886 1004944
rect 266268 1004896 266320 1004902
rect 266268 1004838 266320 1004844
rect 266280 997257 266308 1004838
rect 267738 1004728 267794 1004737
rect 267738 1004663 267794 1004672
rect 266266 997248 266322 997257
rect 266266 997183 266322 997192
rect 267648 996124 267700 996130
rect 267648 996066 267700 996072
rect 265256 996056 265308 996062
rect 265256 995998 265308 996004
rect 267556 996056 267608 996062
rect 267556 995998 267608 996004
rect 248326 993647 248382 993656
rect 262220 993676 262272 993682
rect 231584 993618 231636 993624
rect 235632 989460 235684 989466
rect 235632 989402 235684 989408
rect 227628 987216 227680 987222
rect 227628 987158 227680 987164
rect 219084 983606 219466 983634
rect 235644 983620 235672 989402
rect 248340 988174 248368 993647
rect 262220 993618 262272 993624
rect 248328 988168 248380 988174
rect 248328 988110 248380 988116
rect 251824 988168 251876 988174
rect 251824 988110 251876 988116
rect 251836 983620 251864 988110
rect 267568 987290 267596 995998
rect 267660 987426 267688 996066
rect 267648 987420 267700 987426
rect 267648 987362 267700 987368
rect 267556 987284 267608 987290
rect 267556 987226 267608 987232
rect 267752 983634 267780 1004663
rect 267844 996198 267872 1004935
rect 269026 1004864 269082 1004873
rect 269026 1004799 269082 1004808
rect 267832 996192 267884 996198
rect 267832 996134 267884 996140
rect 269040 989466 269068 1004799
rect 269224 989534 269252 1005071
rect 270408 996192 270460 996198
rect 270408 996134 270460 996140
rect 269212 989528 269264 989534
rect 269212 989470 269264 989476
rect 269028 989460 269080 989466
rect 269028 989402 269080 989408
rect 270420 987494 270448 996134
rect 280080 987562 280108 1005314
rect 280252 1005304 280304 1005310
rect 280252 1005246 280304 1005252
rect 360198 1005272 360254 1005281
rect 280160 1004964 280212 1004970
rect 280160 1004906 280212 1004912
rect 280172 996198 280200 1004906
rect 280160 996192 280212 996198
rect 280160 996134 280212 996140
rect 280264 996062 280292 1005246
rect 360198 1005207 360200 1005216
rect 360252 1005207 360254 1005216
rect 360200 1005178 360252 1005184
rect 358176 1005032 358228 1005038
rect 350262 1005000 350318 1005009
rect 350262 1004935 350318 1004944
rect 353666 1005000 353722 1005009
rect 353666 1004935 353722 1004944
rect 358174 1005000 358176 1005009
rect 358228 1005000 358230 1005009
rect 358174 1004935 358230 1004944
rect 280344 1004760 280396 1004766
rect 280344 1004702 280396 1004708
rect 304078 1004728 304134 1004737
rect 280356 996130 280384 1004702
rect 304446 1004728 304502 1004737
rect 304134 1004686 304446 1004714
rect 304078 1004663 304134 1004672
rect 304446 1004663 304502 1004672
rect 315118 1004728 315174 1004737
rect 315118 1004663 315120 1004672
rect 315172 1004663 315174 1004672
rect 321466 1004728 321522 1004737
rect 321466 1004663 321522 1004672
rect 331220 1004692 331272 1004698
rect 315120 1004634 315172 1004640
rect 312176 999864 312228 999870
rect 311438 999832 311494 999841
rect 311438 999767 311440 999776
rect 311492 999767 311494 999776
rect 312174 999832 312176 999841
rect 318892 999864 318944 999870
rect 312228 999832 312230 999841
rect 318892 999806 318944 999812
rect 312174 999767 312230 999776
rect 315948 999796 316000 999802
rect 311440 999738 311492 999744
rect 315948 999738 316000 999744
rect 313832 999728 313884 999734
rect 310150 999696 310206 999705
rect 310150 999631 310152 999640
rect 310204 999631 310206 999640
rect 313830 999696 313832 999705
rect 313884 999696 313886 999705
rect 313830 999631 313886 999640
rect 314936 999660 314988 999666
rect 310152 999602 310204 999608
rect 314936 999602 314988 999608
rect 313004 999592 313056 999598
rect 313002 999560 313004 999569
rect 313056 999560 313058 999569
rect 313002 999495 313058 999504
rect 314658 999560 314714 999569
rect 314658 999495 314660 999504
rect 314712 999495 314714 999504
rect 314660 999466 314712 999472
rect 309784 999456 309836 999462
rect 309782 999424 309784 999433
rect 314844 999456 314896 999462
rect 309836 999424 309838 999433
rect 309782 999359 309838 999368
rect 312634 999424 312690 999433
rect 314844 999398 314896 999404
rect 312634 999359 312636 999368
rect 312688 999359 312690 999368
rect 312636 999330 312688 999336
rect 310980 999320 311032 999326
rect 310978 999288 310980 999297
rect 311032 999288 311034 999297
rect 310978 999223 311034 999232
rect 311806 999288 311862 999297
rect 311806 999223 311808 999232
rect 311860 999223 311862 999232
rect 311808 999194 311860 999200
rect 314292 999184 314344 999190
rect 314290 999152 314292 999161
rect 314344 999152 314346 999161
rect 298744 999116 298796 999122
rect 314290 999087 314346 999096
rect 298744 999058 298796 999064
rect 298756 997257 298784 999058
rect 298742 997248 298798 997257
rect 298742 997183 298798 997192
rect 301780 996328 301832 996334
rect 308128 996328 308180 996334
rect 301780 996270 301832 996276
rect 308126 996296 308128 996305
rect 308180 996296 308182 996305
rect 300216 996260 300268 996266
rect 300216 996202 300268 996208
rect 280344 996124 280396 996130
rect 280344 996066 280396 996072
rect 280252 996056 280304 996062
rect 280252 995998 280304 996004
rect 286784 995852 286836 995858
rect 286784 995794 286836 995800
rect 293592 995852 293644 995858
rect 293592 995794 293644 995800
rect 295064 995852 295116 995858
rect 295064 995794 295116 995800
rect 286796 995738 286824 995794
rect 288070 995752 288126 995761
rect 286534 995710 286824 995738
rect 287822 995710 288070 995738
rect 292486 995752 292542 995761
rect 291502 995722 291792 995738
rect 291502 995716 291804 995722
rect 291502 995710 291752 995716
rect 288070 995687 288126 995696
rect 292146 995710 292486 995738
rect 293604 995738 293632 995794
rect 293342 995710 293632 995738
rect 295076 995738 295104 995794
rect 295076 995710 295182 995738
rect 292486 995687 292542 995696
rect 291752 995658 291804 995664
rect 287520 995648 287572 995654
rect 287178 995596 287520 995602
rect 300228 995625 300256 996202
rect 300766 995888 300822 995897
rect 300766 995823 300822 995832
rect 290646 995616 290702 995625
rect 287178 995590 287572 995596
rect 287178 995574 287560 995590
rect 290306 995574 290646 995602
rect 290646 995551 290702 995560
rect 300214 995616 300270 995625
rect 300214 995551 300270 995560
rect 291106 995480 291162 995489
rect 282840 993682 282868 995452
rect 283484 993886 283512 995452
rect 283472 993880 283524 993886
rect 283472 993822 283524 993828
rect 284128 993750 284156 995452
rect 285968 993818 285996 995452
rect 290858 995438 291106 995466
rect 297270 995480 297326 995489
rect 291106 995415 291162 995424
rect 285956 993812 286008 993818
rect 285956 993754 286008 993760
rect 284116 993744 284168 993750
rect 294524 993721 294552 995452
rect 297022 995438 297270 995466
rect 297270 995415 297326 995424
rect 284116 993686 284168 993692
rect 294510 993712 294566 993721
rect 282828 993676 282880 993682
rect 294510 993647 294566 993656
rect 282828 993618 282880 993624
rect 300492 989528 300544 989534
rect 300492 989470 300544 989476
rect 284300 989460 284352 989466
rect 284300 989402 284352 989408
rect 280068 987556 280120 987562
rect 280068 987498 280120 987504
rect 270408 987488 270460 987494
rect 270408 987430 270460 987436
rect 267752 983606 268134 983634
rect 284312 983620 284340 989402
rect 300504 983620 300532 989470
rect 300780 984774 300808 995823
rect 301792 993886 301820 996270
rect 308126 996231 308182 996240
rect 308954 996296 309010 996305
rect 308954 996231 308956 996240
rect 309008 996231 309010 996240
rect 308956 996202 309008 996208
rect 305274 996160 305330 996169
rect 305274 996095 305330 996104
rect 305734 996160 305790 996169
rect 305734 996095 305790 996104
rect 306470 996160 306526 996169
rect 306470 996095 306526 996104
rect 306930 996160 306986 996169
rect 306930 996095 306986 996104
rect 307298 996160 307354 996169
rect 307298 996095 307354 996104
rect 307758 996160 307814 996169
rect 307758 996095 307814 996104
rect 310150 996160 310206 996169
rect 310150 996095 310206 996104
rect 305288 995625 305316 996095
rect 305274 995616 305330 995625
rect 305274 995551 305330 995560
rect 305748 995353 305776 996095
rect 306484 995722 306512 996095
rect 306944 995926 306972 996095
rect 306932 995920 306984 995926
rect 306932 995862 306984 995868
rect 306472 995716 306524 995722
rect 306472 995658 306524 995664
rect 307312 995654 307340 996095
rect 307772 995994 307800 996095
rect 307760 995988 307812 995994
rect 307760 995930 307812 995936
rect 310164 995858 310192 996095
rect 310152 995852 310204 995858
rect 310152 995794 310204 995800
rect 307300 995648 307352 995654
rect 307300 995590 307352 995596
rect 305734 995344 305790 995353
rect 305734 995279 305790 995288
rect 303528 994772 303580 994778
rect 303528 994714 303580 994720
rect 301780 993880 301832 993886
rect 301780 993822 301832 993828
rect 303540 989466 303568 994714
rect 314856 993818 314884 999398
rect 314844 993812 314896 993818
rect 314844 993754 314896 993760
rect 314948 993682 314976 999602
rect 315028 999320 315080 999326
rect 315028 999262 315080 999268
rect 315040 993750 315068 999262
rect 315120 999252 315172 999258
rect 315120 999194 315172 999200
rect 315132 996062 315160 999194
rect 315120 996056 315172 996062
rect 315120 995998 315172 996004
rect 315028 993744 315080 993750
rect 315028 993686 315080 993692
rect 314936 993676 314988 993682
rect 314936 993618 314988 993624
rect 303528 989460 303580 989466
rect 303528 989402 303580 989408
rect 315132 987630 315160 995998
rect 315120 987624 315172 987630
rect 315120 987566 315172 987572
rect 315960 984842 315988 999738
rect 318708 999728 318760 999734
rect 318708 999670 318760 999676
rect 317604 999592 317656 999598
rect 317604 999534 317656 999540
rect 317420 999388 317472 999394
rect 317420 999330 317472 999336
rect 317432 996198 317460 999330
rect 317512 999184 317564 999190
rect 317512 999126 317564 999132
rect 317420 996192 317472 996198
rect 317420 996134 317472 996140
rect 316774 993848 316830 993857
rect 316774 993783 316830 993792
rect 315948 984836 316000 984842
rect 315948 984778 316000 984784
rect 300768 984768 300820 984774
rect 300768 984710 300820 984716
rect 316788 983620 316816 993783
rect 317432 984910 317460 996134
rect 317524 996130 317552 999126
rect 317616 999122 317644 999534
rect 317604 999116 317656 999122
rect 317604 999058 317656 999064
rect 317512 996124 317564 996130
rect 317512 996066 317564 996072
rect 317524 987766 317552 996066
rect 317512 987760 317564 987766
rect 317512 987702 317564 987708
rect 318720 987698 318748 999670
rect 318904 987834 318932 999806
rect 319076 999524 319128 999530
rect 319076 999466 319128 999472
rect 319088 989534 319116 999466
rect 321480 989602 321508 1004663
rect 331220 1004634 331272 1004640
rect 331232 990690 331260 1004634
rect 331220 990684 331272 990690
rect 331220 990626 331272 990632
rect 332692 990684 332744 990690
rect 332692 990626 332744 990632
rect 321468 989596 321520 989602
rect 321468 989538 321520 989544
rect 319076 989528 319128 989534
rect 319076 989470 319128 989476
rect 318892 987828 318944 987834
rect 318892 987770 318944 987776
rect 318708 987692 318760 987698
rect 318708 987634 318760 987640
rect 317420 984904 317472 984910
rect 317420 984846 317472 984852
rect 332704 983634 332732 990626
rect 349160 989596 349212 989602
rect 349160 989538 349212 989544
rect 332704 983606 332994 983634
rect 349172 983620 349200 989538
rect 350276 985182 350304 1004935
rect 353680 995897 353708 1004935
rect 358544 1004760 358596 1004766
rect 354494 1004728 354550 1004737
rect 354862 1004728 354918 1004737
rect 354550 1004686 354862 1004714
rect 354494 1004663 354550 1004672
rect 354862 1004663 354918 1004672
rect 358542 1004728 358544 1004737
rect 358596 1004728 358598 1004737
rect 358542 1004663 358598 1004672
rect 359738 1004728 359794 1004737
rect 359738 1004663 359740 1004672
rect 359792 1004663 359794 1004672
rect 369860 1004692 369912 1004698
rect 359740 1004634 359792 1004640
rect 369860 1004634 369912 1004640
rect 360566 1000784 360622 1000793
rect 360566 1000719 360568 1000728
rect 360620 1000719 360622 1000728
rect 360568 1000690 360620 1000696
rect 361396 1000680 361448 1000686
rect 361394 1000648 361396 1000657
rect 361448 1000648 361450 1000657
rect 369872 1000618 369900 1004634
rect 373184 1001094 373212 1005586
rect 378048 1005576 378100 1005582
rect 378048 1005518 378100 1005524
rect 376668 1005440 376720 1005446
rect 376668 1005382 376720 1005388
rect 376680 1001162 376708 1005382
rect 377956 1005372 378008 1005378
rect 377956 1005314 378008 1005320
rect 376668 1001156 376720 1001162
rect 376668 1001098 376720 1001104
rect 373172 1001088 373224 1001094
rect 373172 1001030 373224 1001036
rect 361394 1000583 361450 1000592
rect 369860 1000612 369912 1000618
rect 369860 1000554 369912 1000560
rect 358912 1000544 358964 1000550
rect 358910 1000512 358912 1000521
rect 358964 1000512 358966 1000521
rect 358910 1000447 358966 1000456
rect 357346 999288 357402 999297
rect 357346 999223 357348 999232
rect 357400 999223 357402 999232
rect 364892 999252 364944 999258
rect 357348 999194 357400 999200
rect 364892 999194 364944 999200
rect 357716 999184 357768 999190
rect 357714 999152 357716 999161
rect 357768 999152 357770 999161
rect 357714 999087 357770 999096
rect 364904 998510 364932 999194
rect 365076 999184 365128 999190
rect 365076 999126 365128 999132
rect 364892 998504 364944 998510
rect 364892 998446 364944 998452
rect 365088 997830 365116 999126
rect 377968 999002 377996 1005314
rect 378060 999190 378088 1005518
rect 425152 1005440 425204 1005446
rect 425150 1005408 425152 1005417
rect 425204 1005408 425206 1005417
rect 425150 1005343 425206 1005352
rect 428370 1005408 428426 1005417
rect 428370 1005343 428372 1005352
rect 428424 1005343 428426 1005352
rect 428372 1005314 428424 1005320
rect 380808 1005236 380860 1005242
rect 380808 1005178 380860 1005184
rect 380820 1001994 380848 1005178
rect 427544 1005168 427596 1005174
rect 427542 1005136 427544 1005145
rect 427596 1005136 427598 1005145
rect 427542 1005071 427598 1005080
rect 428830 1005136 428886 1005145
rect 428830 1005071 428832 1005080
rect 428884 1005071 428886 1005080
rect 428832 1005042 428884 1005048
rect 383292 1005032 383344 1005038
rect 426808 1005032 426860 1005038
rect 383292 1004974 383344 1004980
rect 425518 1005000 425574 1005009
rect 381728 1004692 381780 1004698
rect 381728 1004634 381780 1004640
rect 380820 1001966 380940 1001994
rect 378324 1001156 378376 1001162
rect 378324 1001098 378376 1001104
rect 378048 999184 378100 999190
rect 378048 999126 378100 999132
rect 377968 998974 378180 999002
rect 374552 998504 374604 998510
rect 374552 998446 374604 998452
rect 365076 997824 365128 997830
rect 365076 997766 365128 997772
rect 374460 997824 374512 997830
rect 374460 997766 374512 997772
rect 363418 997248 363474 997257
rect 363418 997183 363420 997192
rect 363472 997183 363474 997192
rect 367098 997248 367154 997257
rect 367098 997183 367100 997192
rect 363420 997154 363472 997160
rect 367152 997183 367154 997192
rect 367100 997154 367152 997160
rect 365442 996296 365498 996305
rect 365442 996231 365444 996240
rect 365496 996231 365498 996240
rect 371148 996260 371200 996266
rect 365444 996202 365496 996208
rect 371148 996202 371200 996208
rect 364248 996192 364300 996198
rect 362590 996160 362646 996169
rect 362590 996095 362646 996104
rect 364246 996160 364248 996169
rect 367284 996192 367336 996198
rect 364300 996160 364302 996169
rect 364246 996095 364302 996104
rect 364706 996160 364762 996169
rect 364706 996095 364708 996104
rect 362604 995994 362632 996095
rect 364760 996095 364762 996104
rect 365074 996160 365130 996169
rect 367284 996134 367336 996140
rect 365074 996095 365130 996104
rect 364708 996066 364760 996072
rect 365088 996062 365116 996095
rect 365076 996056 365128 996062
rect 365076 995998 365128 996004
rect 362592 995988 362644 995994
rect 362592 995930 362644 995936
rect 353666 995888 353722 995897
rect 353666 995823 353722 995832
rect 367098 995888 367154 995897
rect 367098 995823 367154 995832
rect 359186 995616 359242 995625
rect 359186 995551 359242 995560
rect 359200 993682 359228 995551
rect 366178 993712 366234 993721
rect 359188 993676 359240 993682
rect 366178 993647 366234 993656
rect 359188 993618 359240 993624
rect 366192 989738 366220 993647
rect 366180 989732 366232 989738
rect 366180 989674 366232 989680
rect 365444 989528 365496 989534
rect 365444 989470 365496 989476
rect 350264 985176 350316 985182
rect 350264 985118 350316 985124
rect 365456 983620 365484 989470
rect 367112 985114 367140 995823
rect 367190 995752 367246 995761
rect 367190 995687 367246 995696
rect 367204 988038 367232 995687
rect 367296 993478 367324 996134
rect 369860 996124 369912 996130
rect 369860 996066 369912 996072
rect 367376 995988 367428 995994
rect 367376 995930 367428 995936
rect 367388 993546 367416 995930
rect 367466 995616 367522 995625
rect 367466 995551 367522 995560
rect 367376 993540 367428 993546
rect 367376 993482 367428 993488
rect 367284 993472 367336 993478
rect 367284 993414 367336 993420
rect 367480 992594 367508 995551
rect 368572 993540 368624 993546
rect 368572 993482 368624 993488
rect 368388 993472 368440 993478
rect 368388 993414 368440 993420
rect 367468 992588 367520 992594
rect 367468 992530 367520 992536
rect 367192 988032 367244 988038
rect 367192 987974 367244 987980
rect 367100 985108 367152 985114
rect 367100 985050 367152 985056
rect 368400 984978 368428 993414
rect 368584 985046 368612 993482
rect 368756 993472 368808 993478
rect 368756 993414 368808 993420
rect 368768 992594 368796 993414
rect 368756 992588 368808 992594
rect 368756 992530 368808 992536
rect 368768 987970 368796 992530
rect 368756 987964 368808 987970
rect 368756 987906 368808 987912
rect 369872 987902 369900 996066
rect 371160 989670 371188 996202
rect 371514 996160 371570 996169
rect 371514 996095 371570 996104
rect 371332 996056 371384 996062
rect 371332 995998 371384 996004
rect 371148 989664 371200 989670
rect 371148 989606 371200 989612
rect 371344 989534 371372 995998
rect 371528 989602 371556 996095
rect 374472 993721 374500 997766
rect 374564 993750 374592 998446
rect 378152 993857 378180 998974
rect 378336 993886 378364 1001098
rect 380912 1000346 380940 1001966
rect 381268 1001088 381320 1001094
rect 381268 1001030 381320 1001036
rect 380900 1000340 380952 1000346
rect 380900 1000282 380952 1000288
rect 381280 995450 381308 1001030
rect 381740 996441 381768 1004634
rect 383200 999184 383252 999190
rect 383200 999126 383252 999132
rect 381726 996432 381782 996441
rect 381726 996367 381782 996376
rect 383212 995926 383240 999126
rect 383200 995920 383252 995926
rect 383200 995862 383252 995868
rect 383304 995518 383332 1004974
rect 425518 1004935 425520 1004944
rect 425572 1004935 425574 1004944
rect 426806 1005000 426808 1005009
rect 426860 1005000 426862 1005009
rect 426806 1004935 426862 1004944
rect 425520 1004906 425572 1004912
rect 427176 1004896 427228 1004902
rect 423494 1004864 423550 1004873
rect 423494 1004799 423496 1004808
rect 423548 1004799 423550 1004808
rect 427174 1004864 427176 1004873
rect 427228 1004864 427230 1004873
rect 427174 1004799 427230 1004808
rect 423496 1004770 423548 1004776
rect 422312 1004737 422340 1004763
rect 424692 1004760 424744 1004766
rect 422298 1004728 422354 1004737
rect 419448 1004692 419500 1004698
rect 422666 1004728 422722 1004737
rect 422354 1004686 422666 1004714
rect 422298 1004663 422300 1004672
rect 419448 1004634 419500 1004640
rect 422352 1004663 422354 1004672
rect 422666 1004663 422722 1004672
rect 424690 1004728 424692 1004737
rect 424744 1004728 424746 1004737
rect 424690 1004663 424746 1004672
rect 422300 1004634 422352 1004640
rect 383568 1000748 383620 1000754
rect 383568 1000690 383620 1000696
rect 383384 1000680 383436 1000686
rect 383384 1000622 383436 1000628
rect 383580 1000634 383608 1000690
rect 383396 995654 383424 1000622
rect 383476 1000612 383528 1000618
rect 383580 1000606 383792 1000634
rect 383476 1000554 383528 1000560
rect 383488 995994 383516 1000554
rect 383568 1000544 383620 1000550
rect 383620 1000492 383700 1000498
rect 383568 1000486 383700 1000492
rect 383580 1000470 383700 1000486
rect 383568 1000340 383620 1000346
rect 383568 1000282 383620 1000288
rect 383476 995988 383528 995994
rect 383476 995930 383528 995936
rect 383384 995648 383436 995654
rect 383384 995590 383436 995596
rect 383580 995586 383608 1000282
rect 383672 995790 383700 1000470
rect 383660 995784 383712 995790
rect 383660 995726 383712 995732
rect 383764 995722 383792 1000606
rect 400036 999184 400088 999190
rect 400036 999126 400088 999132
rect 399944 999116 399996 999122
rect 399944 999058 399996 999064
rect 399956 997257 399984 999058
rect 399942 997248 399998 997257
rect 399942 997183 399998 997192
rect 400048 995858 400076 999126
rect 391940 995852 391992 995858
rect 391940 995794 391992 995800
rect 396632 995852 396684 995858
rect 396632 995794 396684 995800
rect 400036 995852 400088 995858
rect 400036 995794 400088 995800
rect 384948 995784 385000 995790
rect 384408 995722 384698 995738
rect 389364 995784 389416 995790
rect 388166 995752 388222 995761
rect 385000 995732 385342 995738
rect 384948 995726 385342 995732
rect 383752 995716 383804 995722
rect 383752 995658 383804 995664
rect 384396 995716 384698 995722
rect 384448 995710 384698 995716
rect 384960 995710 385342 995726
rect 388222 995710 388378 995738
rect 391952 995738 391980 995794
rect 396644 995738 396672 995794
rect 389416 995732 389666 995738
rect 389364 995726 389666 995732
rect 389376 995710 389666 995726
rect 391952 995710 392150 995738
rect 396382 995710 396672 995738
rect 388166 995687 388222 995696
rect 384396 995658 384448 995664
rect 385684 995648 385736 995654
rect 385736 995596 385986 995602
rect 385684 995590 385986 995596
rect 383568 995580 383620 995586
rect 385696 995574 385986 995590
rect 387536 995586 387826 995602
rect 387524 995580 387826 995586
rect 383568 995522 383620 995528
rect 387576 995574 387826 995580
rect 387524 995522 387576 995528
rect 383292 995512 383344 995518
rect 383292 995454 383344 995460
rect 388628 995512 388680 995518
rect 393596 995512 393648 995518
rect 388680 995460 389022 995466
rect 388628 995454 389022 995460
rect 393648 995460 393990 995466
rect 393596 995454 393990 995460
rect 381268 995444 381320 995450
rect 388640 995438 389022 995454
rect 381268 995386 381320 995392
rect 392688 993886 392716 995452
rect 378324 993880 378376 993886
rect 378138 993848 378194 993857
rect 378324 993822 378376 993828
rect 392676 993880 392728 993886
rect 392676 993822 392728 993828
rect 378138 993783 378194 993792
rect 393332 993750 393360 995452
rect 393608 995438 393990 995454
rect 374552 993744 374604 993750
rect 374458 993712 374514 993721
rect 374552 993686 374604 993692
rect 393320 993744 393372 993750
rect 395172 993721 395200 995452
rect 397012 993857 397040 995452
rect 396998 993848 397054 993857
rect 396998 993783 397054 993792
rect 393320 993686 393372 993692
rect 395158 993712 395214 993721
rect 374458 993647 374514 993656
rect 398852 993682 398880 995452
rect 395158 993647 395214 993656
rect 398840 993676 398892 993682
rect 398840 993618 398892 993624
rect 381636 989732 381688 989738
rect 381636 989674 381688 989680
rect 371516 989596 371568 989602
rect 371516 989538 371568 989544
rect 371332 989528 371384 989534
rect 371332 989470 371384 989476
rect 369860 987896 369912 987902
rect 369860 987838 369912 987844
rect 368572 985040 368624 985046
rect 368572 984982 368624 984988
rect 368388 984972 368440 984978
rect 368388 984914 368440 984920
rect 381648 983620 381676 989674
rect 397828 989664 397880 989670
rect 397828 989606 397880 989612
rect 397840 983620 397868 989606
rect 414112 989596 414164 989602
rect 414112 989538 414164 989544
rect 414124 983620 414152 989538
rect 419460 984978 419488 1004634
rect 440252 1001978 440280 1005790
rect 440436 1002046 440464 1005858
rect 453948 1005372 454000 1005378
rect 453948 1005314 454000 1005320
rect 440424 1002040 440476 1002046
rect 440424 1001982 440476 1001988
rect 440240 1001972 440292 1001978
rect 440240 1001914 440292 1001920
rect 447140 1001904 447192 1001910
rect 447140 1001846 447192 1001852
rect 447324 1001904 447376 1001910
rect 447324 1001846 447376 1001852
rect 428002 1000648 428058 1000657
rect 428002 1000583 428004 1000592
rect 428056 1000583 428058 1000592
rect 428004 1000554 428056 1000560
rect 426348 1000544 426400 1000550
rect 426346 1000512 426348 1000521
rect 426400 1000512 426402 1000521
rect 426346 1000447 426402 1000456
rect 434628 999864 434680 999870
rect 430854 999832 430910 999841
rect 434628 999806 434680 999812
rect 430854 999767 430856 999776
rect 430908 999767 430910 999776
rect 430856 999738 430908 999744
rect 431684 999728 431736 999734
rect 429198 999696 429254 999705
rect 429198 999631 429200 999640
rect 429252 999631 429254 999640
rect 431682 999696 431684 999705
rect 431736 999696 431738 999705
rect 431682 999631 431738 999640
rect 429200 999602 429252 999608
rect 430028 999592 430080 999598
rect 430026 999560 430028 999569
rect 430080 999560 430082 999569
rect 430026 999495 430082 999504
rect 431222 999560 431278 999569
rect 431222 999495 431224 999504
rect 431276 999495 431278 999504
rect 431224 999466 431276 999472
rect 429660 999456 429712 999462
rect 429658 999424 429660 999433
rect 433432 999456 433484 999462
rect 429712 999424 429714 999433
rect 429658 999359 429714 999368
rect 432510 999424 432566 999433
rect 433432 999398 433484 999404
rect 432510 999359 432512 999368
rect 432564 999359 432566 999368
rect 432512 999330 432564 999336
rect 432880 999320 432932 999326
rect 432050 999288 432106 999297
rect 432050 999223 432052 999232
rect 432104 999223 432106 999232
rect 432878 999288 432880 999297
rect 432932 999288 432934 999297
rect 432878 999223 432934 999232
rect 432052 999194 432104 999200
rect 430396 999184 430448 999190
rect 430394 999152 430396 999161
rect 433340 999184 433392 999190
rect 430448 999152 430450 999161
rect 433340 999126 433392 999132
rect 430394 999087 430450 999096
rect 433352 993546 433380 999126
rect 433340 993540 433392 993546
rect 433340 993482 433392 993488
rect 433444 993478 433472 999398
rect 433524 993608 433576 993614
rect 433524 993550 433576 993556
rect 433432 993472 433484 993478
rect 433432 993414 433484 993420
rect 430304 989528 430356 989534
rect 430304 989470 430356 989476
rect 419448 984972 419500 984978
rect 419448 984914 419500 984920
rect 430316 983620 430344 989470
rect 433536 987358 433564 993550
rect 433616 993540 433668 993546
rect 433616 993482 433668 993488
rect 433524 987352 433576 987358
rect 433524 987294 433576 987300
rect 433628 984706 433656 993482
rect 434640 989738 434668 999806
rect 438124 999796 438176 999802
rect 438124 999738 438176 999744
rect 437940 999728 437992 999734
rect 437940 999670 437992 999676
rect 434720 999660 434772 999666
rect 434720 999602 434772 999608
rect 434732 993614 434760 999602
rect 434812 999592 434864 999598
rect 434812 999534 434864 999540
rect 434720 993608 434772 993614
rect 434720 993550 434772 993556
rect 434824 993546 434852 999534
rect 436192 999524 436244 999530
rect 436192 999466 436244 999472
rect 436100 999252 436152 999258
rect 436100 999194 436152 999200
rect 434812 993540 434864 993546
rect 434812 993482 434864 993488
rect 436112 993410 436140 999194
rect 436204 999122 436232 999466
rect 437388 999388 437440 999394
rect 437388 999330 437440 999336
rect 436192 999116 436244 999122
rect 436192 999058 436244 999064
rect 436192 993472 436244 993478
rect 436192 993414 436244 993420
rect 436100 993404 436152 993410
rect 436100 993346 436152 993352
rect 434628 989732 434680 989738
rect 434628 989674 434680 989680
rect 433616 984700 433668 984706
rect 433616 984642 433668 984648
rect 436204 984638 436232 993414
rect 437400 989534 437428 999330
rect 437572 999320 437624 999326
rect 437572 999262 437624 999268
rect 437584 989670 437612 999262
rect 437754 999152 437810 999161
rect 437754 999087 437810 999096
rect 437572 989664 437624 989670
rect 437572 989606 437624 989612
rect 437768 989602 437796 999087
rect 437952 993478 437980 999670
rect 438136 997121 438164 999738
rect 438122 997112 438178 997121
rect 438122 997047 438178 997056
rect 447152 995761 447180 1001846
rect 447138 995752 447194 995761
rect 447138 995687 447194 995696
rect 447336 993721 447364 1001846
rect 453960 999122 453988 1005314
rect 455604 1005032 455656 1005038
rect 455604 1004974 455656 1004980
rect 455420 1004964 455472 1004970
rect 455420 1004906 455472 1004912
rect 455432 1003406 455460 1004906
rect 455512 1004896 455564 1004902
rect 455512 1004838 455564 1004844
rect 455420 1003400 455472 1003406
rect 455420 1003342 455472 1003348
rect 455524 1003338 455552 1004838
rect 455512 1003332 455564 1003338
rect 455512 1003274 455564 1003280
rect 455616 1003270 455644 1004974
rect 458928 1004698 458956 1005994
rect 504548 1005712 504600 1005718
rect 504546 1005680 504548 1005689
rect 519728 1005712 519780 1005718
rect 504600 1005680 504602 1005689
rect 504546 1005615 504602 1005624
rect 505006 1005680 505062 1005689
rect 519728 1005654 519780 1005660
rect 505006 1005615 505008 1005624
rect 505060 1005615 505062 1005624
rect 517428 1005644 517480 1005650
rect 505008 1005586 505060 1005592
rect 517428 1005586 517480 1005592
rect 505376 1005576 505428 1005582
rect 502982 1005544 503038 1005553
rect 502982 1005479 502984 1005488
rect 503036 1005479 503038 1005488
rect 505374 1005544 505376 1005553
rect 505428 1005544 505430 1005553
rect 505374 1005479 505430 1005488
rect 502984 1005450 503036 1005456
rect 467932 1005440 467984 1005446
rect 467932 1005382 467984 1005388
rect 505834 1005408 505890 1005417
rect 460848 1005168 460900 1005174
rect 460848 1005110 460900 1005116
rect 458916 1004692 458968 1004698
rect 458916 1004634 458968 1004640
rect 455604 1003264 455656 1003270
rect 455604 1003206 455656 1003212
rect 460860 1001858 460888 1005110
rect 465264 1005100 465316 1005106
rect 465264 1005042 465316 1005048
rect 464252 1003400 464304 1003406
rect 464252 1003342 464304 1003348
rect 460860 1001830 461072 1001858
rect 453948 999116 454000 999122
rect 453948 999058 454000 999064
rect 461044 996441 461072 1001830
rect 464264 1001774 464292 1003342
rect 464252 1001768 464304 1001774
rect 464252 1001710 464304 1001716
rect 465276 999190 465304 1005042
rect 467748 1004828 467800 1004834
rect 467748 1004770 467800 1004776
rect 466460 1003264 466512 1003270
rect 466460 1003206 466512 1003212
rect 466472 1001910 466500 1003206
rect 466460 1001904 466512 1001910
rect 466460 1001846 466512 1001852
rect 465264 999184 465316 999190
rect 465264 999126 465316 999132
rect 462596 999116 462648 999122
rect 462596 999058 462648 999064
rect 461030 996432 461086 996441
rect 461030 996367 461086 996376
rect 447322 993712 447378 993721
rect 462608 993682 462636 999058
rect 467760 998102 467788 1004770
rect 467840 1004760 467892 1004766
rect 467840 1004702 467892 1004708
rect 467852 998374 467880 1004702
rect 467840 998368 467892 998374
rect 467840 998310 467892 998316
rect 467944 998238 467972 1005382
rect 505834 1005343 505836 1005352
rect 505888 1005343 505890 1005352
rect 517060 1005372 517112 1005378
rect 505836 1005314 505888 1005320
rect 517060 1005314 517112 1005320
rect 502522 1005136 502578 1005145
rect 502522 1005071 502524 1005080
rect 502576 1005071 502578 1005080
rect 502524 1005042 502576 1005048
rect 504180 1005032 504232 1005038
rect 504178 1005000 504180 1005009
rect 504232 1005000 504234 1005009
rect 504178 1004935 504234 1004944
rect 499316 1004737 499344 1004763
rect 501696 1004760 501748 1004766
rect 499302 1004728 499358 1004737
rect 472348 1004692 472400 1004698
rect 472348 1004634 472400 1004640
rect 496728 1004692 496780 1004698
rect 499670 1004728 499726 1004737
rect 499358 1004686 499670 1004714
rect 499302 1004663 499304 1004672
rect 496728 1004634 496780 1004640
rect 499356 1004663 499358 1004672
rect 499670 1004663 499726 1004672
rect 501694 1004728 501696 1004737
rect 509148 1004760 509200 1004766
rect 501748 1004728 501750 1004737
rect 501694 1004663 501750 1004672
rect 502154 1004728 502210 1004737
rect 509148 1004702 509200 1004708
rect 502154 1004663 502156 1004672
rect 499304 1004634 499356 1004640
rect 502208 1004663 502210 1004672
rect 502156 1004634 502208 1004640
rect 469128 1003332 469180 1003338
rect 469128 1003274 469180 1003280
rect 469140 999134 469168 1003274
rect 469772 1001904 469824 1001910
rect 469772 1001846 469824 1001852
rect 469140 999106 469444 999134
rect 469220 998368 469272 998374
rect 469220 998310 469272 998316
rect 467932 998232 467984 998238
rect 467932 998174 467984 998180
rect 467748 998096 467800 998102
rect 467748 998038 467800 998044
rect 469232 995654 469260 998310
rect 469312 998096 469364 998102
rect 469312 998038 469364 998044
rect 469220 995648 469272 995654
rect 469220 995590 469272 995596
rect 469324 995586 469352 998038
rect 469312 995580 469364 995586
rect 469312 995522 469364 995528
rect 469416 995353 469444 999106
rect 469402 995344 469458 995353
rect 469402 995279 469458 995288
rect 469784 993818 469812 1001846
rect 471704 1001768 471756 1001774
rect 471704 1001710 471756 1001716
rect 471060 998232 471112 998238
rect 471060 998174 471112 998180
rect 469772 993812 469824 993818
rect 469772 993754 469824 993760
rect 471072 993750 471100 998174
rect 471716 995625 471744 1001710
rect 472360 995722 472388 1004634
rect 472624 1000612 472676 1000618
rect 472624 1000554 472676 1000560
rect 472532 1000544 472584 1000550
rect 472532 1000486 472584 1000492
rect 472440 999184 472492 999190
rect 472440 999126 472492 999132
rect 472452 995926 472480 999126
rect 472440 995920 472492 995926
rect 472440 995862 472492 995868
rect 472544 995858 472572 1000486
rect 472532 995852 472584 995858
rect 472532 995794 472584 995800
rect 472636 995790 472664 1000554
rect 488908 999184 488960 999190
rect 488908 999126 488960 999132
rect 488920 995858 488948 999126
rect 489460 999116 489512 999122
rect 489460 999058 489512 999064
rect 489472 997121 489500 999058
rect 489458 997112 489514 997121
rect 489458 997047 489514 997056
rect 474004 995852 474056 995858
rect 474004 995794 474056 995800
rect 474740 995852 474792 995858
rect 474740 995794 474792 995800
rect 485688 995852 485740 995858
rect 485688 995794 485740 995800
rect 488908 995852 488960 995858
rect 488908 995794 488960 995800
rect 472624 995784 472676 995790
rect 472624 995726 472676 995732
rect 473268 995784 473320 995790
rect 474016 995738 474044 995794
rect 474752 995738 474780 995794
rect 481454 995752 481510 995761
rect 473320 995732 473662 995738
rect 473268 995726 473662 995732
rect 472348 995716 472400 995722
rect 473280 995710 473662 995726
rect 474016 995710 474306 995738
rect 474752 995710 474950 995738
rect 476960 995722 477342 995738
rect 476948 995716 477342 995722
rect 472348 995658 472400 995664
rect 477000 995710 477342 995716
rect 485700 995738 485728 995794
rect 481510 995710 481666 995738
rect 485346 995710 485728 995738
rect 481454 995687 481510 995696
rect 476948 995658 477000 995664
rect 481916 995648 481968 995654
rect 471702 995616 471758 995625
rect 471702 995551 471758 995560
rect 477682 995616 477738 995625
rect 477738 995574 477986 995602
rect 481968 995596 482310 995602
rect 481916 995590 482310 995596
rect 481928 995574 482310 995590
rect 482664 995586 482954 995602
rect 482652 995580 482954 995586
rect 477682 995551 477738 995560
rect 482704 995574 482954 995580
rect 482652 995522 482704 995528
rect 476486 995480 476542 995489
rect 476542 995438 476790 995466
rect 476486 995415 476542 995424
rect 471060 993744 471112 993750
rect 478616 993721 478644 995452
rect 481100 995353 481128 995452
rect 481086 995344 481142 995353
rect 481086 995279 481142 995288
rect 484136 993750 484164 995452
rect 484124 993744 484176 993750
rect 471060 993686 471112 993692
rect 478602 993712 478658 993721
rect 447322 993647 447378 993656
rect 462596 993676 462648 993682
rect 484124 993686 484176 993692
rect 485976 993682 486004 995452
rect 487816 993818 487844 995452
rect 487804 993812 487856 993818
rect 487804 993754 487856 993760
rect 478602 993647 478658 993656
rect 485964 993676 486016 993682
rect 462596 993618 462648 993624
rect 485964 993618 486016 993624
rect 437940 993472 437992 993478
rect 437940 993414 437992 993420
rect 446496 989732 446548 989738
rect 446496 989674 446548 989680
rect 437756 989596 437808 989602
rect 437756 989538 437808 989544
rect 437388 989528 437440 989534
rect 437388 989470 437440 989476
rect 436192 984632 436244 984638
rect 436192 984574 436244 984580
rect 446508 983620 446536 989674
rect 462780 989664 462832 989670
rect 462780 989606 462832 989612
rect 462792 983620 462820 989606
rect 478972 989596 479024 989602
rect 478972 989538 479024 989544
rect 478984 983620 479012 989538
rect 495164 989528 495216 989534
rect 495164 989470 495216 989476
rect 495176 983620 495204 989470
rect 496740 984638 496768 1004634
rect 503352 1000000 503404 1000006
rect 503350 999968 503352 999977
rect 503404 999968 503406 999977
rect 503350 999903 503406 999912
rect 508686 999832 508742 999841
rect 508686 999767 508688 999776
rect 508740 999767 508742 999776
rect 508688 999738 508740 999744
rect 506204 999728 506256 999734
rect 506202 999696 506204 999705
rect 506256 999696 506258 999705
rect 506202 999631 506258 999640
rect 507030 999696 507086 999705
rect 507030 999631 507032 999640
rect 507084 999631 507086 999640
rect 507032 999602 507084 999608
rect 508228 999592 508280 999598
rect 507858 999560 507914 999569
rect 507858 999495 507860 999504
rect 507912 999495 507914 999504
rect 508226 999560 508228 999569
rect 508280 999560 508282 999569
rect 508226 999495 508282 999504
rect 507860 999466 507912 999472
rect 506572 999456 506624 999462
rect 500498 999424 500554 999433
rect 500498 999359 500500 999368
rect 500552 999359 500554 999368
rect 506570 999424 506572 999433
rect 506624 999424 506626 999433
rect 509054 999424 509110 999433
rect 506570 999359 506626 999368
rect 508780 999388 508832 999394
rect 500500 999330 500552 999336
rect 509054 999359 509056 999368
rect 508780 999330 508832 999336
rect 509108 999359 509110 999368
rect 509056 999330 509108 999336
rect 500866 999288 500922 999297
rect 500866 999223 500868 999232
rect 500920 999223 500922 999232
rect 507398 999288 507454 999297
rect 507398 999223 507400 999232
rect 500868 999194 500920 999200
rect 507452 999223 507454 999232
rect 507400 999194 507452 999200
rect 505652 999184 505704 999190
rect 505652 999126 505704 999132
rect 501326 997792 501382 997801
rect 501326 997727 501328 997736
rect 501380 997727 501382 997736
rect 501328 997698 501380 997704
rect 503626 995616 503682 995625
rect 503626 995551 503682 995560
rect 503640 993682 503668 995551
rect 503628 993676 503680 993682
rect 503628 993618 503680 993624
rect 505664 988310 505692 999126
rect 508792 999054 508820 999330
rect 508780 999048 508832 999054
rect 508780 998990 508832 998996
rect 509160 998986 509188 1004702
rect 509240 1004692 509292 1004698
rect 509240 1004634 509292 1004640
rect 509148 998980 509200 998986
rect 509148 998922 509200 998928
rect 509252 998918 509280 1004634
rect 517072 1001910 517100 1005314
rect 517440 1004630 517468 1005586
rect 518808 1005576 518860 1005582
rect 518808 1005518 518860 1005524
rect 517428 1004624 517480 1004630
rect 517428 1004566 517480 1004572
rect 517060 1001904 517112 1001910
rect 517060 1001846 517112 1001852
rect 516048 1000000 516100 1000006
rect 516046 999968 516048 999977
rect 516100 999968 516102 999977
rect 516046 999903 516102 999912
rect 515220 999796 515272 999802
rect 515220 999738 515272 999744
rect 511908 999728 511960 999734
rect 511908 999670 511960 999676
rect 510896 999456 510948 999462
rect 510896 999398 510948 999404
rect 509516 999320 509568 999326
rect 509514 999288 509516 999297
rect 509568 999288 509570 999297
rect 509514 999223 509570 999232
rect 510712 999252 510764 999258
rect 510712 999194 510764 999200
rect 509516 999184 509568 999190
rect 509884 999184 509936 999190
rect 509516 999126 509568 999132
rect 509882 999152 509884 999161
rect 509936 999152 509938 999161
rect 509240 998912 509292 998918
rect 509240 998854 509292 998860
rect 509528 998850 509556 999126
rect 509882 999087 509938 999096
rect 509516 998844 509568 998850
rect 509516 998786 509568 998792
rect 510724 993546 510752 999194
rect 510908 993614 510936 999398
rect 510896 993608 510948 993614
rect 510896 993550 510948 993556
rect 510988 993608 511040 993614
rect 510988 993550 511040 993556
rect 510712 993540 510764 993546
rect 510712 993482 510764 993488
rect 510804 993540 510856 993546
rect 510804 993482 510856 993488
rect 505652 988304 505704 988310
rect 505652 988246 505704 988252
rect 496728 984632 496780 984638
rect 496728 984574 496780 984580
rect 510816 984434 510844 993482
rect 511000 984502 511028 993550
rect 511920 993546 511948 999670
rect 512092 999660 512144 999666
rect 512092 999602 512144 999608
rect 512104 993614 512132 999602
rect 513472 999592 513524 999598
rect 513472 999534 513524 999540
rect 512276 999524 512328 999530
rect 512276 999466 512328 999472
rect 512288 996198 512316 999466
rect 513484 999122 513512 999534
rect 513656 999388 513708 999394
rect 513656 999330 513708 999336
rect 513472 999116 513524 999122
rect 513472 999058 513524 999064
rect 512276 996192 512328 996198
rect 512276 996134 512328 996140
rect 512092 993608 512144 993614
rect 512092 993550 512144 993556
rect 511908 993540 511960 993546
rect 511908 993482 511960 993488
rect 513668 993478 513696 999330
rect 514852 999320 514904 999326
rect 514852 999262 514904 999268
rect 514668 999184 514720 999190
rect 514668 999126 514720 999132
rect 513656 993472 513708 993478
rect 513656 993414 513708 993420
rect 513748 993472 513800 993478
rect 513748 993414 513800 993420
rect 511448 988304 511500 988310
rect 511448 988246 511500 988252
rect 510988 984496 511040 984502
rect 510988 984438 511040 984444
rect 510804 984428 510856 984434
rect 510804 984370 510856 984376
rect 511460 983620 511488 988246
rect 513760 984366 513788 993414
rect 514680 989670 514708 999126
rect 514668 989664 514720 989670
rect 514668 989606 514720 989612
rect 514864 989534 514892 999262
rect 515034 999152 515090 999161
rect 515034 999087 515090 999096
rect 515048 989602 515076 999087
rect 515232 993478 515260 999738
rect 518820 999134 518848 1005518
rect 519084 1005032 519136 1005038
rect 519084 1004974 519136 1004980
rect 519096 999161 519124 1004974
rect 519740 1001910 519768 1005654
rect 523040 1005508 523092 1005514
rect 523040 1005450 523092 1005456
rect 519544 1001904 519596 1001910
rect 519544 1001846 519596 1001852
rect 519728 1001904 519780 1001910
rect 519728 1001846 519780 1001852
rect 519082 999152 519138 999161
rect 518820 999106 518940 999134
rect 518912 998238 518940 999106
rect 519082 999087 519138 999096
rect 518900 998232 518952 998238
rect 518900 998174 518952 998180
rect 519556 996441 519584 1001846
rect 521292 999048 521344 999054
rect 521292 998990 521344 998996
rect 520556 998912 520608 998918
rect 520556 998854 520608 998860
rect 519542 996432 519598 996441
rect 519542 996367 519598 996376
rect 520568 993818 520596 998854
rect 521304 995353 521332 998990
rect 521384 998980 521436 998986
rect 521384 998922 521436 998928
rect 521396 995586 521424 998922
rect 521476 998844 521528 998850
rect 521476 998786 521528 998792
rect 521488 995654 521516 998786
rect 521660 998232 521712 998238
rect 521660 998174 521712 998180
rect 521568 997756 521620 997762
rect 521568 997698 521620 997704
rect 521476 995648 521528 995654
rect 521580 995625 521608 997698
rect 521476 995590 521528 995596
rect 521566 995616 521622 995625
rect 521384 995580 521436 995586
rect 521566 995551 521622 995560
rect 521384 995522 521436 995528
rect 521290 995344 521346 995353
rect 521290 995279 521346 995288
rect 521672 995217 521700 998174
rect 523052 995926 523080 1005450
rect 523224 1005100 523276 1005106
rect 523224 1005042 523276 1005048
rect 523040 995920 523092 995926
rect 523040 995862 523092 995868
rect 523236 995722 523264 1005042
rect 546314 1005000 546370 1005009
rect 546314 1004935 546370 1004944
rect 549442 1005000 549498 1005009
rect 549442 1004935 549498 1004944
rect 552754 1005000 552810 1005009
rect 552754 1004935 552756 1004944
rect 523960 1004624 524012 1004630
rect 523960 1004566 524012 1004572
rect 523868 1001904 523920 1001910
rect 523868 1001846 523920 1001852
rect 523774 999152 523830 999161
rect 523774 999087 523830 999096
rect 523788 996577 523816 999087
rect 523774 996568 523830 996577
rect 523774 996503 523830 996512
rect 523880 995761 523908 1001846
rect 523972 995858 524000 1004566
rect 524050 999968 524106 999977
rect 524050 999903 524106 999912
rect 523960 995852 524012 995858
rect 523960 995794 524012 995800
rect 524064 995790 524092 999903
rect 540336 999252 540388 999258
rect 540336 999194 540388 999200
rect 540348 995858 540376 999194
rect 524788 995852 524840 995858
rect 524788 995794 524840 995800
rect 528468 995852 528520 995858
rect 528468 995794 528520 995800
rect 537024 995852 537076 995858
rect 537024 995794 537076 995800
rect 540336 995852 540388 995858
rect 540336 995794 540388 995800
rect 524052 995784 524104 995790
rect 523866 995752 523922 995761
rect 523224 995716 523276 995722
rect 524052 995726 524104 995732
rect 524800 995738 524828 995794
rect 525340 995784 525392 995790
rect 524800 995710 525090 995738
rect 527914 995752 527970 995761
rect 525392 995732 525734 995738
rect 525340 995726 525734 995732
rect 525352 995710 525734 995726
rect 523866 995687 523922 995696
rect 528480 995738 528508 995794
rect 532238 995752 532294 995761
rect 527970 995710 528218 995738
rect 528480 995710 528770 995738
rect 529032 995722 529414 995738
rect 529020 995716 529414 995722
rect 527914 995687 527970 995696
rect 523224 995658 523276 995664
rect 529072 995710 529414 995716
rect 537036 995738 537064 995794
rect 532294 995710 532542 995738
rect 536774 995710 537064 995738
rect 532238 995687 532294 995696
rect 529020 995658 529072 995664
rect 532700 995648 532752 995654
rect 530122 995616 530178 995625
rect 530058 995574 530122 995602
rect 532752 995596 533094 995602
rect 532700 995590 533094 995596
rect 532712 995574 533094 995590
rect 533448 995586 533738 995602
rect 533436 995580 533738 995586
rect 530122 995551 530178 995560
rect 533488 995574 533738 995580
rect 533436 995522 533488 995528
rect 526166 995480 526222 995489
rect 526222 995438 526378 995466
rect 534000 995438 534382 995466
rect 526166 995415 526222 995424
rect 534000 995353 534028 995438
rect 533986 995344 534042 995353
rect 533986 995279 534042 995288
rect 521658 995208 521714 995217
rect 521658 995143 521714 995152
rect 535564 993818 535592 995452
rect 537404 995353 537432 995452
rect 537390 995344 537446 995353
rect 537390 995279 537446 995288
rect 520556 993812 520608 993818
rect 520556 993754 520608 993760
rect 535552 993812 535604 993818
rect 535552 993754 535604 993760
rect 539244 993682 539272 995452
rect 539232 993676 539284 993682
rect 539232 993618 539284 993624
rect 515220 993472 515272 993478
rect 515220 993414 515272 993420
rect 527640 989664 527692 989670
rect 527640 989606 527692 989612
rect 515036 989596 515088 989602
rect 515036 989538 515088 989544
rect 514852 989528 514904 989534
rect 514852 989470 514904 989476
rect 513748 984360 513800 984366
rect 513748 984302 513800 984308
rect 527652 983620 527680 989606
rect 543832 989596 543884 989602
rect 543832 989538 543884 989544
rect 543844 983620 543872 989538
rect 546328 984366 546356 1004935
rect 549456 995897 549484 1004935
rect 552808 1004935 552810 1004944
rect 568580 1004964 568632 1004970
rect 552756 1004906 552808 1004912
rect 568580 1004906 568632 1004912
rect 553122 1004864 553178 1004873
rect 553122 1004799 553124 1004808
rect 553176 1004799 553178 1004808
rect 557448 1004828 557500 1004834
rect 553124 1004770 553176 1004776
rect 557448 1004770 557500 1004776
rect 551928 1004760 551980 1004766
rect 550270 1004728 550326 1004737
rect 550638 1004728 550694 1004737
rect 550326 1004686 550638 1004714
rect 550270 1004663 550326 1004672
rect 550638 1004663 550694 1004672
rect 551926 1004728 551928 1004737
rect 551980 1004728 551982 1004737
rect 551926 1004663 551982 1004672
rect 554318 1004728 554374 1004737
rect 554318 1004663 554320 1004672
rect 554372 1004663 554374 1004672
rect 554320 1004634 554372 1004640
rect 557460 1004154 557488 1004770
rect 558736 1004760 558788 1004766
rect 558736 1004702 558788 1004708
rect 561310 1004728 561366 1004737
rect 557448 1004148 557500 1004154
rect 557448 1004090 557500 1004096
rect 553952 1003944 554004 1003950
rect 553950 1003912 553952 1003921
rect 554004 1003912 554006 1003921
rect 553950 1003847 554006 1003856
rect 555514 1003368 555570 1003377
rect 555514 1003303 555516 1003312
rect 555568 1003303 555570 1003312
rect 555516 1003274 555568 1003280
rect 554780 1003264 554832 1003270
rect 554778 1003232 554780 1003241
rect 554832 1003232 554834 1003241
rect 554778 1003167 554834 1003176
rect 558748 1001910 558776 1004702
rect 561310 1004663 561312 1004672
rect 561364 1004663 561366 1004672
rect 567290 1004728 567346 1004737
rect 567290 1004663 567346 1004672
rect 567476 1004692 567528 1004698
rect 561312 1004634 561364 1004640
rect 558736 1001904 558788 1001910
rect 558736 1001846 558788 1001852
rect 566556 1000068 566608 1000074
rect 566556 1000010 566608 1000016
rect 560850 999832 560906 999841
rect 560850 999767 560852 999776
rect 560904 999767 560906 999776
rect 560852 999738 560904 999744
rect 560482 999696 560538 999705
rect 560482 999631 560484 999640
rect 560536 999631 560538 999640
rect 565820 999660 565872 999666
rect 560484 999602 560536 999608
rect 565820 999602 565872 999608
rect 552296 999184 552348 999190
rect 552294 999152 552296 999161
rect 558920 999184 558972 999190
rect 552348 999152 552350 999161
rect 558920 999126 558972 999132
rect 552294 999087 552350 999096
rect 558932 997966 558960 999126
rect 558920 997960 558972 997966
rect 558920 997902 558972 997908
rect 553490 997792 553546 997801
rect 553490 997727 553492 997736
rect 553544 997727 553546 997736
rect 553492 997698 553544 997704
rect 556344 997688 556396 997694
rect 556342 997656 556344 997665
rect 556396 997656 556398 997665
rect 556342 997591 556398 997600
rect 557170 997520 557226 997529
rect 557170 997455 557172 997464
rect 557224 997455 557226 997464
rect 557172 997426 557224 997432
rect 559288 996192 559340 996198
rect 558458 996160 558514 996169
rect 558458 996095 558460 996104
rect 558512 996095 558514 996104
rect 559286 996160 559288 996169
rect 559340 996160 559342 996169
rect 559286 996095 559342 996104
rect 564440 996124 564492 996130
rect 558460 996066 558512 996072
rect 564440 996066 564492 996072
rect 549442 995888 549498 995897
rect 549442 995823 549498 995832
rect 557722 995752 557778 995761
rect 557722 995687 557778 995696
rect 558550 995752 558606 995761
rect 558550 995687 558606 995696
rect 564346 995752 564402 995761
rect 564346 995687 564402 995696
rect 555054 995616 555110 995625
rect 555054 995551 555110 995560
rect 555068 993682 555096 995551
rect 555056 993676 555108 993682
rect 555056 993618 555108 993624
rect 557736 993546 557764 995687
rect 558564 993614 558592 995687
rect 561678 995616 561734 995625
rect 561678 995551 561734 995560
rect 561494 995480 561550 995489
rect 561494 995415 561550 995424
rect 561310 995344 561366 995353
rect 561310 995279 561366 995288
rect 561324 993857 561352 995279
rect 561310 993848 561366 993857
rect 561310 993783 561366 993792
rect 561508 993721 561536 995415
rect 561494 993712 561550 993721
rect 561494 993647 561550 993656
rect 558552 993608 558604 993614
rect 558552 993550 558604 993556
rect 557724 993540 557776 993546
rect 557724 993482 557776 993488
rect 560116 989528 560168 989534
rect 560116 989470 560168 989476
rect 546316 984360 546368 984366
rect 546316 984302 546368 984308
rect 560128 983620 560156 989470
rect 561692 985697 561720 995551
rect 561678 985688 561734 985697
rect 561678 985623 561734 985632
rect 561692 984094 561720 985623
rect 564360 984094 564388 995687
rect 564452 985833 564480 996066
rect 564714 995888 564770 995897
rect 564714 995823 564770 995832
rect 564438 985824 564494 985833
rect 564438 985759 564494 985768
rect 561680 984088 561732 984094
rect 561680 984030 561732 984036
rect 564348 984088 564400 984094
rect 564348 984030 564400 984036
rect 564452 983958 564480 985759
rect 564728 985590 564756 995823
rect 565832 993478 565860 999602
rect 566568 995994 566596 1000010
rect 567108 999796 567160 999802
rect 567108 999738 567160 999744
rect 566556 995988 566608 995994
rect 566556 995930 566608 995936
rect 565820 993472 565872 993478
rect 565820 993414 565872 993420
rect 567120 989534 567148 999738
rect 567304 989602 567332 1004663
rect 567476 1004634 567528 1004640
rect 567488 989670 567516 1004634
rect 568592 1001842 568620 1004906
rect 571340 1004624 571392 1004630
rect 571340 1004566 571392 1004572
rect 570144 1004148 570196 1004154
rect 570144 1004090 570196 1004096
rect 569960 1003264 570012 1003270
rect 569960 1003206 570012 1003212
rect 569868 1001904 569920 1001910
rect 569868 1001846 569920 1001852
rect 568580 1001836 568632 1001842
rect 568580 1001778 568632 1001784
rect 568672 997960 568724 997966
rect 568672 997902 568724 997908
rect 568580 997756 568632 997762
rect 568580 997698 568632 997704
rect 568592 994129 568620 997698
rect 568684 994265 568712 997902
rect 569880 997762 569908 1001846
rect 569868 997756 569920 997762
rect 569868 997698 569920 997704
rect 569972 997558 570000 1003206
rect 569960 997552 570012 997558
rect 569960 997494 570012 997500
rect 568670 994256 568726 994265
rect 568670 994191 568726 994200
rect 568578 994120 568634 994129
rect 568578 994055 568634 994064
rect 570156 993993 570184 1004090
rect 571352 997626 571380 1004566
rect 571432 1003944 571484 1003950
rect 571432 1003886 571484 1003892
rect 571340 997620 571392 997626
rect 571340 997562 571392 997568
rect 571444 997422 571472 1003886
rect 574008 1003332 574060 1003338
rect 574008 1003274 574060 1003280
rect 572628 1001836 572680 1001842
rect 572628 1001778 572680 1001784
rect 571432 997416 571484 997422
rect 571432 997358 571484 997364
rect 572640 997354 572668 1001778
rect 574020 999002 574048 1003274
rect 590660 999524 590712 999530
rect 590660 999466 590712 999472
rect 625804 999524 625856 999530
rect 625804 999466 625856 999472
rect 574020 998974 574140 999002
rect 572628 997348 572680 997354
rect 572628 997290 572680 997296
rect 570142 993984 570198 993993
rect 570142 993919 570198 993928
rect 574112 993750 574140 998974
rect 590672 997422 590700 999466
rect 610072 999456 610124 999462
rect 610072 999398 610124 999404
rect 625712 999456 625764 999462
rect 625712 999398 625764 999404
rect 625816 999410 625844 999466
rect 609980 999388 610032 999394
rect 609980 999330 610032 999336
rect 601608 999320 601660 999326
rect 601608 999262 601660 999268
rect 593420 999252 593472 999258
rect 593420 999194 593472 999200
rect 590660 997416 590712 997422
rect 590660 997358 590712 997364
rect 593432 997354 593460 999194
rect 601620 997694 601648 999262
rect 601608 997688 601660 997694
rect 601608 997630 601660 997636
rect 609992 997626 610020 999330
rect 609980 997620 610032 997626
rect 609980 997562 610032 997568
rect 610084 997558 610112 999398
rect 625620 999388 625672 999394
rect 625620 999330 625672 999336
rect 625528 999252 625580 999258
rect 625528 999194 625580 999200
rect 623780 997756 623832 997762
rect 623780 997698 623832 997704
rect 610072 997552 610124 997558
rect 610072 997494 610124 997500
rect 620928 997484 620980 997490
rect 620928 997426 620980 997432
rect 593420 997348 593472 997354
rect 593420 997290 593472 997296
rect 576308 995988 576360 995994
rect 576308 995930 576360 995936
rect 574100 993744 574152 993750
rect 574100 993686 574152 993692
rect 567476 989664 567528 989670
rect 567476 989606 567528 989612
rect 567292 989596 567344 989602
rect 567292 989538 567344 989544
rect 567108 989528 567160 989534
rect 567108 989470 567160 989476
rect 564532 985584 564584 985590
rect 564532 985526 564584 985532
rect 564716 985584 564768 985590
rect 564716 985526 564768 985532
rect 564544 984026 564572 985526
rect 564532 984020 564584 984026
rect 564532 983962 564584 983968
rect 564440 983952 564492 983958
rect 564440 983894 564492 983900
rect 576320 983620 576348 995930
rect 620940 995790 620968 997426
rect 620928 995784 620980 995790
rect 620928 995726 620980 995732
rect 623792 995654 623820 997698
rect 625540 996062 625568 999194
rect 625528 996056 625580 996062
rect 625528 995998 625580 996004
rect 625632 995994 625660 999330
rect 625620 995988 625672 995994
rect 625620 995930 625672 995936
rect 625724 995926 625752 999398
rect 625816 999382 625936 999410
rect 625804 999320 625856 999326
rect 625804 999262 625856 999268
rect 625712 995920 625764 995926
rect 625712 995862 625764 995868
rect 625816 995858 625844 999262
rect 625804 995852 625856 995858
rect 625804 995794 625856 995800
rect 625908 995722 625936 999382
rect 626540 995852 626592 995858
rect 626540 995794 626592 995800
rect 627184 995852 627236 995858
rect 627184 995794 627236 995800
rect 630220 995852 630272 995858
rect 630220 995794 630272 995800
rect 631508 995852 631560 995858
rect 631508 995794 631560 995800
rect 626552 995738 626580 995794
rect 627196 995738 627224 995794
rect 627828 995784 627880 995790
rect 625896 995716 625948 995722
rect 626552 995710 626888 995738
rect 627196 995710 627532 995738
rect 630232 995738 630260 995794
rect 631520 995738 631548 995794
rect 627880 995732 628176 995738
rect 627828 995726 628176 995732
rect 627840 995710 628176 995726
rect 630232 995710 630568 995738
rect 630876 995722 631212 995738
rect 630864 995716 631212 995722
rect 625896 995658 625948 995664
rect 630916 995710 631212 995716
rect 631520 995710 631856 995738
rect 630864 995658 630916 995664
rect 623780 995648 623832 995654
rect 623780 995590 623832 995596
rect 635832 995648 635884 995654
rect 635884 995596 636180 995602
rect 635832 995590 636180 995596
rect 635844 995574 636180 995590
rect 629680 995438 630016 995466
rect 634004 995438 634340 995466
rect 634832 995438 634892 995466
rect 635200 995438 635536 995466
rect 637040 995438 637376 995466
rect 629680 993857 629708 995438
rect 629666 993848 629722 993857
rect 629666 993783 629722 993792
rect 634004 993750 634032 995438
rect 634832 994265 634860 995438
rect 634818 994256 634874 994265
rect 634818 994191 634874 994200
rect 635200 993993 635228 995438
rect 637040 994129 637068 995438
rect 638558 995217 638586 995452
rect 638880 995438 639216 995466
rect 640720 995438 641056 995466
rect 638544 995208 638600 995217
rect 638544 995143 638600 995152
rect 637026 994120 637082 994129
rect 637026 994055 637082 994064
rect 635186 993984 635242 993993
rect 635186 993919 635242 993928
rect 633992 993744 634044 993750
rect 638880 993721 638908 995438
rect 633992 993686 634044 993692
rect 638866 993712 638922 993721
rect 640720 993682 640748 995438
rect 641166 995208 641222 995217
rect 641166 995143 641222 995152
rect 638866 993647 638922 993656
rect 640708 993676 640760 993682
rect 640708 993618 640760 993624
rect 592500 989664 592552 989670
rect 592500 989606 592552 989612
rect 592512 983620 592540 989606
rect 608784 989596 608836 989602
rect 608784 989538 608836 989544
rect 608796 983620 608824 989538
rect 624976 989528 625028 989534
rect 624976 989470 625028 989476
rect 624988 983620 625016 989470
rect 641180 983620 641208 995143
rect 666560 989460 666612 989466
rect 666560 989402 666612 989408
rect 651380 987556 651432 987562
rect 651380 987498 651432 987504
rect 649908 984088 649960 984094
rect 649908 984030 649960 984036
rect 649920 935678 649948 984030
rect 649908 935672 649960 935678
rect 649908 935614 649960 935620
rect 62854 814192 62910 814201
rect 62854 814127 62910 814136
rect 62856 772880 62908 772886
rect 62856 772822 62908 772828
rect 62764 684480 62816 684486
rect 62764 684422 62816 684428
rect 62762 427952 62818 427961
rect 62762 427887 62818 427896
rect 62776 278254 62804 427887
rect 62764 278248 62816 278254
rect 62764 278190 62816 278196
rect 62670 278080 62726 278089
rect 62670 278015 62726 278024
rect 62868 277953 62896 772822
rect 63222 729872 63278 729881
rect 63222 729807 63278 729816
rect 63040 728748 63092 728754
rect 63040 728690 63092 728696
rect 62948 427848 63000 427854
rect 62948 427790 63000 427796
rect 62960 278186 62988 427790
rect 62948 278180 63000 278186
rect 62948 278122 63000 278128
rect 62854 277944 62910 277953
rect 62854 277879 62910 277888
rect 63052 277817 63080 728690
rect 63132 386436 63184 386442
rect 63132 386378 63184 386384
rect 63144 278050 63172 386378
rect 63132 278044 63184 278050
rect 63132 277986 63184 277992
rect 63038 277808 63094 277817
rect 63038 277743 63094 277752
rect 63236 277681 63264 729807
rect 63314 383888 63370 383897
rect 63314 383823 63370 383832
rect 63328 278118 63356 383823
rect 63316 278112 63368 278118
rect 63316 278054 63368 278060
rect 63222 277672 63278 277681
rect 63222 277607 63278 277616
rect 65904 271862 65932 277780
rect 67008 271930 67036 277780
rect 66996 271924 67048 271930
rect 66996 271866 67048 271872
rect 65892 271856 65944 271862
rect 65892 271798 65944 271804
rect 68204 266354 68232 277780
rect 69400 269113 69428 277780
rect 70596 271833 70624 277780
rect 70582 271824 70638 271833
rect 70582 271759 70638 271768
rect 71792 269210 71820 277780
rect 71780 269204 71832 269210
rect 71780 269146 71832 269152
rect 69386 269104 69442 269113
rect 69386 269039 69442 269048
rect 72988 266490 73016 277780
rect 74092 269482 74120 277780
rect 75288 271998 75316 277780
rect 75276 271992 75328 271998
rect 76484 271969 76512 277780
rect 75276 271934 75328 271940
rect 76470 271960 76526 271969
rect 76470 271895 76526 271904
rect 74080 269476 74132 269482
rect 74080 269418 74132 269424
rect 77680 269249 77708 277780
rect 78876 269385 78904 277780
rect 80072 269414 80100 277780
rect 80060 269408 80112 269414
rect 78862 269376 78918 269385
rect 80060 269350 80112 269356
rect 78862 269311 78918 269320
rect 81268 269278 81296 277780
rect 82372 269346 82400 277780
rect 83568 272105 83596 277780
rect 83554 272096 83610 272105
rect 83554 272031 83610 272040
rect 84764 269521 84792 277780
rect 85960 272241 85988 277780
rect 85946 272232 86002 272241
rect 85946 272167 86002 272176
rect 87156 269793 87184 277780
rect 87142 269784 87198 269793
rect 87142 269719 87198 269728
rect 84750 269512 84806 269521
rect 84750 269447 84806 269456
rect 82360 269340 82412 269346
rect 82360 269282 82412 269288
rect 81256 269272 81308 269278
rect 77666 269240 77722 269249
rect 81256 269214 81308 269220
rect 77666 269175 77722 269184
rect 88352 267986 88380 277780
rect 89548 272066 89576 277780
rect 89536 272060 89588 272066
rect 89536 272002 89588 272008
rect 90652 269657 90680 277780
rect 91848 272377 91876 277780
rect 91834 272368 91890 272377
rect 91834 272303 91890 272312
rect 93044 272202 93072 277780
rect 93032 272196 93084 272202
rect 93032 272138 93084 272144
rect 90638 269648 90694 269657
rect 90638 269583 90694 269592
rect 94240 269550 94268 277780
rect 95436 269686 95464 277780
rect 96632 269929 96660 277780
rect 97736 272785 97764 277780
rect 97722 272776 97778 272785
rect 97722 272711 97778 272720
rect 98932 272513 98960 277780
rect 100128 272649 100156 277780
rect 100114 272640 100170 272649
rect 100114 272575 100170 272584
rect 98918 272504 98974 272513
rect 98918 272439 98974 272448
rect 101324 270065 101352 277780
rect 101310 270056 101366 270065
rect 101310 269991 101366 270000
rect 96618 269920 96674 269929
rect 96618 269855 96674 269864
rect 95424 269680 95476 269686
rect 95424 269622 95476 269628
rect 102520 269618 102548 277780
rect 103716 270201 103744 277780
rect 104912 272134 104940 277780
rect 106016 272921 106044 277780
rect 107212 273057 107240 277780
rect 107198 273048 107254 273057
rect 107198 272983 107254 272992
rect 106002 272912 106058 272921
rect 106002 272847 106058 272856
rect 104900 272128 104952 272134
rect 104900 272070 104952 272076
rect 108408 270337 108436 277780
rect 108394 270328 108450 270337
rect 108394 270263 108450 270272
rect 103702 270192 103758 270201
rect 103702 270127 103758 270136
rect 109604 269754 109632 277780
rect 110800 269822 110828 277780
rect 111996 273193 112024 277780
rect 111982 273184 112038 273193
rect 111982 273119 112038 273128
rect 110788 269816 110840 269822
rect 110788 269758 110840 269764
rect 109592 269748 109644 269754
rect 109592 269690 109644 269696
rect 102508 269612 102560 269618
rect 102508 269554 102560 269560
rect 94228 269544 94280 269550
rect 94228 269486 94280 269492
rect 88340 267980 88392 267986
rect 88340 267922 88392 267928
rect 72976 266484 73028 266490
rect 72976 266426 73028 266432
rect 113192 266422 113220 277780
rect 114296 269890 114324 277780
rect 115492 271697 115520 277780
rect 115478 271688 115534 271697
rect 115478 271623 115534 271632
rect 114284 269884 114336 269890
rect 114284 269826 114336 269832
rect 116688 266558 116716 277780
rect 117884 272270 117912 277780
rect 117872 272264 117924 272270
rect 117872 272206 117924 272212
rect 119080 269958 119108 277780
rect 120276 271794 120304 277780
rect 120264 271788 120316 271794
rect 120264 271730 120316 271736
rect 121380 270473 121408 277780
rect 122576 271561 122604 277780
rect 122562 271552 122618 271561
rect 122562 271487 122618 271496
rect 121366 270464 121422 270473
rect 121366 270399 121422 270408
rect 119068 269952 119120 269958
rect 119068 269894 119120 269900
rect 123772 266626 123800 277780
rect 124968 272406 124996 277780
rect 124956 272400 125008 272406
rect 124956 272342 125008 272348
rect 126164 270026 126192 277780
rect 126152 270020 126204 270026
rect 126152 269962 126204 269968
rect 127360 268841 127388 277780
rect 128556 268977 128584 277780
rect 129660 272338 129688 277780
rect 129648 272332 129700 272338
rect 129648 272274 129700 272280
rect 130856 271726 130884 277780
rect 132052 272474 132080 277780
rect 132040 272468 132092 272474
rect 132040 272410 132092 272416
rect 130844 271720 130896 271726
rect 130844 271662 130896 271668
rect 133248 270230 133276 277780
rect 133236 270224 133288 270230
rect 133236 270166 133288 270172
rect 134444 270094 134472 277780
rect 135640 270162 135668 277780
rect 136836 272542 136864 277780
rect 137940 272610 137968 277780
rect 139136 272678 139164 277780
rect 139124 272672 139176 272678
rect 139124 272614 139176 272620
rect 137928 272604 137980 272610
rect 137928 272546 137980 272552
rect 136824 272536 136876 272542
rect 136824 272478 136876 272484
rect 140332 270298 140360 277780
rect 141528 270366 141556 277780
rect 141516 270360 141568 270366
rect 141516 270302 141568 270308
rect 140320 270292 140372 270298
rect 140320 270234 140372 270240
rect 135628 270156 135680 270162
rect 135628 270098 135680 270104
rect 134432 270088 134484 270094
rect 134432 270030 134484 270036
rect 128542 268968 128598 268977
rect 128542 268903 128598 268912
rect 127346 268832 127402 268841
rect 127346 268767 127402 268776
rect 142724 268705 142752 277780
rect 143920 272882 143948 277780
rect 143908 272876 143960 272882
rect 143908 272818 143960 272824
rect 145024 272814 145052 277780
rect 145012 272808 145064 272814
rect 145012 272750 145064 272756
rect 146220 272746 146248 277780
rect 146208 272740 146260 272746
rect 146208 272682 146260 272688
rect 147416 270434 147444 277780
rect 148612 273086 148640 277780
rect 148600 273080 148652 273086
rect 148600 273022 148652 273028
rect 149808 273018 149836 277780
rect 149796 273012 149848 273018
rect 149796 272954 149848 272960
rect 151004 272950 151032 277780
rect 150992 272944 151044 272950
rect 150992 272886 151044 272892
rect 152200 270502 152228 277780
rect 152188 270496 152240 270502
rect 152188 270438 152240 270444
rect 147404 270428 147456 270434
rect 147404 270370 147456 270376
rect 142710 268696 142766 268705
rect 142710 268631 142766 268640
rect 153304 268569 153332 277780
rect 154500 269074 154528 277780
rect 155696 273154 155724 277780
rect 155684 273148 155736 273154
rect 155684 273090 155736 273096
rect 156892 271794 156920 277780
rect 156788 271788 156840 271794
rect 156788 271730 156840 271736
rect 156880 271788 156932 271794
rect 156880 271730 156932 271736
rect 154488 269068 154540 269074
rect 154488 269010 154540 269016
rect 153290 268560 153346 268569
rect 156800 268530 156828 271730
rect 158088 271522 158116 277780
rect 158076 271516 158128 271522
rect 158076 271458 158128 271464
rect 159284 269006 159312 277780
rect 159272 269000 159324 269006
rect 159272 268942 159324 268948
rect 160480 268938 160508 277780
rect 160468 268932 160520 268938
rect 160468 268874 160520 268880
rect 161584 268870 161612 277780
rect 162780 271318 162808 277780
rect 163976 271590 164004 277780
rect 165172 271658 165200 277780
rect 165160 271652 165212 271658
rect 165160 271594 165212 271600
rect 163964 271584 164016 271590
rect 163964 271526 164016 271532
rect 162768 271312 162820 271318
rect 162768 271254 162820 271260
rect 161572 268864 161624 268870
rect 161572 268806 161624 268812
rect 166368 268802 166396 277780
rect 166356 268796 166408 268802
rect 166356 268738 166408 268744
rect 167564 268734 167592 277780
rect 167552 268728 167604 268734
rect 167552 268670 167604 268676
rect 168668 268598 168696 277780
rect 169864 271114 169892 277780
rect 171060 271454 171088 277780
rect 171048 271448 171100 271454
rect 171048 271390 171100 271396
rect 172256 271386 172284 277780
rect 172244 271380 172296 271386
rect 172244 271322 172296 271328
rect 169852 271108 169904 271114
rect 169852 271050 169904 271056
rect 173452 268666 173480 277780
rect 173440 268660 173492 268666
rect 173440 268602 173492 268608
rect 168656 268592 168708 268598
rect 168656 268534 168708 268540
rect 153290 268495 153346 268504
rect 156788 268524 156840 268530
rect 156788 268466 156840 268472
rect 174648 268462 174676 277780
rect 175844 270842 175872 277780
rect 176948 271046 176976 277780
rect 177856 273148 177908 273154
rect 177856 273090 177908 273096
rect 177868 271794 177896 273090
rect 178144 272066 178172 277780
rect 178040 272060 178092 272066
rect 178040 272002 178092 272008
rect 178132 272060 178184 272066
rect 178132 272002 178184 272008
rect 177856 271788 177908 271794
rect 177856 271730 177908 271736
rect 177948 271788 178000 271794
rect 177948 271730 178000 271736
rect 177960 271522 177988 271730
rect 177948 271516 178000 271522
rect 177948 271458 178000 271464
rect 178052 271250 178080 272002
rect 178132 271516 178184 271522
rect 178132 271458 178184 271464
rect 178144 271318 178172 271458
rect 178132 271312 178184 271318
rect 178132 271254 178184 271260
rect 178040 271244 178092 271250
rect 178040 271186 178092 271192
rect 179340 271182 179368 277780
rect 180064 271380 180116 271386
rect 180064 271322 180116 271328
rect 179328 271176 179380 271182
rect 179328 271118 179380 271124
rect 180076 271114 180104 271322
rect 180064 271108 180116 271114
rect 180064 271050 180116 271056
rect 176936 271040 176988 271046
rect 176936 270982 176988 270988
rect 175832 270836 175884 270842
rect 175832 270778 175884 270784
rect 179328 270836 179380 270842
rect 179328 270778 179380 270784
rect 174636 268456 174688 268462
rect 174636 268398 174688 268404
rect 179340 268394 179368 270778
rect 179328 268388 179380 268394
rect 179328 268330 179380 268336
rect 180536 268258 180564 277780
rect 181732 268326 181760 277780
rect 182928 271114 182956 277780
rect 182916 271108 182968 271114
rect 182916 271050 182968 271056
rect 181720 268320 181772 268326
rect 181720 268262 181772 268268
rect 180524 268252 180576 268258
rect 180524 268194 180576 268200
rect 184124 268190 184152 277780
rect 184940 272196 184992 272202
rect 184940 272138 184992 272144
rect 184952 268433 184980 272138
rect 185228 270978 185256 277780
rect 185216 270972 185268 270978
rect 185216 270914 185268 270920
rect 186424 270910 186452 277780
rect 186412 270904 186464 270910
rect 186412 270846 186464 270852
rect 187620 270774 187648 277780
rect 188816 272202 188844 277780
rect 188804 272196 188856 272202
rect 188804 272138 188856 272144
rect 189264 271244 189316 271250
rect 189264 271186 189316 271192
rect 187608 270768 187660 270774
rect 187608 270710 187660 270716
rect 184938 268424 184994 268433
rect 184938 268359 184994 268368
rect 184112 268184 184164 268190
rect 184112 268126 184164 268132
rect 189276 268054 189304 271186
rect 190012 270842 190040 277780
rect 190000 270836 190052 270842
rect 190000 270778 190052 270784
rect 191208 270706 191236 277780
rect 192116 271856 192168 271862
rect 192116 271798 192168 271804
rect 191196 270700 191248 270706
rect 191196 270642 191248 270648
rect 189264 268048 189316 268054
rect 189264 267990 189316 267996
rect 123760 266620 123812 266626
rect 123760 266562 123812 266568
rect 116676 266552 116728 266558
rect 116676 266494 116728 266500
rect 113180 266416 113232 266422
rect 113180 266358 113232 266364
rect 68192 266348 68244 266354
rect 68192 266290 68244 266296
rect 192128 264330 192156 271798
rect 192312 270570 192340 277780
rect 192484 271924 192536 271930
rect 192484 271866 192536 271872
rect 192300 270564 192352 270570
rect 192300 270506 192352 270512
rect 192496 264330 192524 271866
rect 193508 269142 193536 277780
rect 194138 271824 194194 271833
rect 194138 271759 194194 271768
rect 194506 271824 194562 271833
rect 194506 271759 194508 271768
rect 193496 269136 193548 269142
rect 193496 269078 193548 269084
rect 193678 269104 193734 269113
rect 193678 269039 193734 269048
rect 193220 266348 193272 266354
rect 193220 266290 193272 266296
rect 192128 264302 192418 264330
rect 192496 264302 192786 264330
rect 193232 264316 193260 266290
rect 193692 264316 193720 269039
rect 194152 264316 194180 271759
rect 194560 271759 194562 271768
rect 194508 271730 194560 271736
rect 194704 271726 194732 277780
rect 195428 271992 195480 271998
rect 195428 271934 195480 271940
rect 194692 271720 194744 271726
rect 194692 271662 194744 271668
rect 194600 269204 194652 269210
rect 194600 269146 194652 269152
rect 194612 264316 194640 269146
rect 195060 266484 195112 266490
rect 195060 266426 195112 266432
rect 195072 264316 195100 266426
rect 195440 264316 195468 271934
rect 195900 269634 195928 277780
rect 197110 277766 197400 277794
rect 197268 272060 197320 272066
rect 197268 272002 197320 272008
rect 196346 271960 196402 271969
rect 196346 271895 196402 271904
rect 195808 269606 195928 269634
rect 195808 269210 195836 269606
rect 195888 269476 195940 269482
rect 195888 269418 195940 269424
rect 195796 269204 195848 269210
rect 195796 269146 195848 269152
rect 195900 264316 195928 269418
rect 196360 264316 196388 271895
rect 197176 271856 197228 271862
rect 197176 271798 197228 271804
rect 196806 269240 196862 269249
rect 196806 269175 196862 269184
rect 196820 264316 196848 269175
rect 197188 268122 197216 271798
rect 197280 271250 197308 272002
rect 197268 271244 197320 271250
rect 197268 271186 197320 271192
rect 197372 269414 197400 277766
rect 198292 271862 198320 277780
rect 199106 272096 199162 272105
rect 199488 272066 199516 277780
rect 199934 272232 199990 272241
rect 199934 272167 199990 272176
rect 199106 272031 199162 272040
rect 199476 272060 199528 272066
rect 198280 271856 198332 271862
rect 198280 271798 198332 271804
rect 198648 270564 198700 270570
rect 198648 270506 198700 270512
rect 198660 269482 198688 270506
rect 199014 269512 199070 269521
rect 198648 269476 198700 269482
rect 199014 269447 199070 269456
rect 198648 269418 198700 269424
rect 197268 269408 197320 269414
rect 197268 269350 197320 269356
rect 197360 269408 197412 269414
rect 197360 269350 197412 269356
rect 197726 269376 197782 269385
rect 197176 268116 197228 268122
rect 197176 268058 197228 268064
rect 197280 264316 197308 269350
rect 197726 269311 197782 269320
rect 198556 269340 198608 269346
rect 197740 264316 197768 269311
rect 198556 269282 198608 269288
rect 198096 269272 198148 269278
rect 198096 269214 198148 269220
rect 198108 264316 198136 269214
rect 198568 264316 198596 269282
rect 199028 264316 199056 269447
rect 199120 264330 199148 272031
rect 199476 272002 199528 272008
rect 199120 264302 199502 264330
rect 199948 264316 199976 272167
rect 200394 269784 200450 269793
rect 200394 269719 200450 269728
rect 200408 264316 200436 269719
rect 200592 269278 200620 277780
rect 201314 272776 201370 272785
rect 201314 272711 201370 272720
rect 200580 269272 200632 269278
rect 200580 269214 200632 269220
rect 201328 268054 201356 272711
rect 201788 271998 201816 277780
rect 202142 272368 202198 272377
rect 202142 272303 202198 272312
rect 201776 271992 201828 271998
rect 201776 271934 201828 271940
rect 201682 269648 201738 269657
rect 201682 269583 201738 269592
rect 200764 268048 200816 268054
rect 200764 267990 200816 267996
rect 201316 268048 201368 268054
rect 201316 267990 201368 267996
rect 200776 264316 200804 267990
rect 201224 267980 201276 267986
rect 201224 267922 201276 267928
rect 201236 264316 201264 267922
rect 201696 264316 201724 269583
rect 202156 264316 202184 272303
rect 202788 272128 202840 272134
rect 202788 272070 202840 272076
rect 202512 270224 202564 270230
rect 202512 270166 202564 270172
rect 202604 270224 202656 270230
rect 202604 270166 202656 270172
rect 202524 267850 202552 270166
rect 202616 270026 202644 270166
rect 202604 270020 202656 270026
rect 202604 269962 202656 269968
rect 202604 269544 202656 269550
rect 202604 269486 202656 269492
rect 202512 267844 202564 267850
rect 202512 267786 202564 267792
rect 202616 264316 202644 269486
rect 202800 267782 202828 272070
rect 202984 269822 203012 277780
rect 203430 273048 203486 273057
rect 203430 272983 203486 272992
rect 202972 269816 203024 269822
rect 202972 269758 203024 269764
rect 203062 268424 203118 268433
rect 203062 268359 203118 268368
rect 202788 267776 202840 267782
rect 202788 267718 202840 267724
rect 203076 264316 203104 268359
rect 203444 268161 203472 272983
rect 203524 269680 203576 269686
rect 203524 269622 203576 269628
rect 203430 268152 203486 268161
rect 203430 268087 203486 268096
rect 203536 264316 203564 269622
rect 204180 269550 204208 277780
rect 204810 272504 204866 272513
rect 204810 272439 204866 272448
rect 204350 269920 204406 269929
rect 204350 269855 204406 269864
rect 204168 269544 204220 269550
rect 204168 269486 204220 269492
rect 203892 268048 203944 268054
rect 203892 267990 203944 267996
rect 203904 264316 203932 267990
rect 204364 264316 204392 269855
rect 204824 264316 204852 272439
rect 205376 272134 205404 277780
rect 205730 272640 205786 272649
rect 205730 272575 205786 272584
rect 205364 272128 205416 272134
rect 205364 272070 205416 272076
rect 205270 270056 205326 270065
rect 205270 269991 205326 270000
rect 205284 264316 205312 269991
rect 205744 264316 205772 272575
rect 206572 269686 206600 277780
rect 207478 272912 207534 272921
rect 207478 272847 207534 272856
rect 206652 272264 206704 272270
rect 206652 272206 206704 272212
rect 206560 269680 206612 269686
rect 206560 269622 206612 269628
rect 206192 269612 206244 269618
rect 206192 269554 206244 269560
rect 206204 264316 206232 269554
rect 206664 267782 206692 272206
rect 207018 270192 207074 270201
rect 207018 270127 207074 270136
rect 206560 267776 206612 267782
rect 206560 267718 206612 267724
rect 206652 267776 206704 267782
rect 206652 267718 206704 267724
rect 206572 264316 206600 267718
rect 207032 264316 207060 270127
rect 207492 264316 207520 272847
rect 207768 269754 207796 277780
rect 208886 277766 209176 277794
rect 208490 271824 208546 271833
rect 208490 271759 208546 271768
rect 208504 271726 208532 271759
rect 208492 271720 208544 271726
rect 208492 271662 208544 271668
rect 208032 270496 208084 270502
rect 208032 270438 208084 270444
rect 207938 270328 207994 270337
rect 207938 270263 207994 270272
rect 207756 269748 207808 269754
rect 207756 269690 207808 269696
rect 207952 264316 207980 270263
rect 208044 267918 208072 270438
rect 208124 270428 208176 270434
rect 208124 270370 208176 270376
rect 208136 268054 208164 270370
rect 208400 269816 208452 269822
rect 208400 269758 208452 269764
rect 208412 269482 208440 269758
rect 209148 269618 209176 277766
rect 209226 273184 209282 273193
rect 209226 273119 209282 273128
rect 208860 269612 208912 269618
rect 208860 269554 208912 269560
rect 209136 269612 209188 269618
rect 209136 269554 209188 269560
rect 208400 269476 208452 269482
rect 208400 269418 208452 269424
rect 208398 268152 208454 268161
rect 208398 268087 208454 268096
rect 208124 268048 208176 268054
rect 208124 267990 208176 267996
rect 208032 267912 208084 267918
rect 208032 267854 208084 267860
rect 208412 264316 208440 268087
rect 208872 264316 208900 269554
rect 209240 264316 209268 273119
rect 210068 269890 210096 277780
rect 210606 271688 210662 271697
rect 210606 271623 210662 271632
rect 209688 269884 209740 269890
rect 209688 269826 209740 269832
rect 210056 269884 210108 269890
rect 210056 269826 210108 269832
rect 209700 264316 209728 269826
rect 210148 266416 210200 266422
rect 210148 266358 210200 266364
rect 210160 264316 210188 266358
rect 210620 264316 210648 271623
rect 211068 269952 211120 269958
rect 211068 269894 211120 269900
rect 211080 264316 211108 269894
rect 211264 267986 211292 277780
rect 211896 270020 211948 270026
rect 211896 269962 211948 269968
rect 211252 267980 211304 267986
rect 211252 267922 211304 267928
rect 211528 266552 211580 266558
rect 211528 266494 211580 266500
rect 211540 264316 211568 266494
rect 211908 264316 211936 269962
rect 212460 269822 212488 277780
rect 213274 271552 213330 271561
rect 213274 271487 213330 271496
rect 212448 269816 212500 269822
rect 212448 269758 212500 269764
rect 212816 268524 212868 268530
rect 212816 268466 212868 268472
rect 212356 267776 212408 267782
rect 212356 267718 212408 267724
rect 212368 264316 212396 267718
rect 212828 264316 212856 268466
rect 213288 264316 213316 271487
rect 213656 268530 213684 277780
rect 213734 270464 213790 270473
rect 213734 270399 213790 270408
rect 213644 268524 213696 268530
rect 213644 268466 213696 268472
rect 213748 264316 213776 270399
rect 214656 270224 214708 270230
rect 214656 270166 214708 270172
rect 214196 266620 214248 266626
rect 214196 266562 214248 266568
rect 214208 264316 214236 266562
rect 214668 264316 214696 270166
rect 214852 269958 214880 277780
rect 215024 272400 215076 272406
rect 215024 272342 215076 272348
rect 214840 269952 214892 269958
rect 214840 269894 214892 269900
rect 215036 264316 215064 272342
rect 215668 272332 215720 272338
rect 215668 272274 215720 272280
rect 215482 268832 215538 268841
rect 215482 268767 215538 268776
rect 215496 264316 215524 268767
rect 215680 264330 215708 272274
rect 215956 270026 215984 277780
rect 217152 270230 217180 277780
rect 217692 272468 217744 272474
rect 217692 272410 217744 272416
rect 217140 270224 217192 270230
rect 217140 270166 217192 270172
rect 215944 270020 215996 270026
rect 215944 269962 215996 269968
rect 216402 268968 216458 268977
rect 216402 268903 216458 268912
rect 215680 264302 215970 264330
rect 216416 264316 216444 268903
rect 216864 268116 216916 268122
rect 216864 268058 216916 268064
rect 216876 264316 216904 268058
rect 217324 267844 217376 267850
rect 217324 267786 217376 267792
rect 217336 264316 217364 267786
rect 217704 264316 217732 272410
rect 218152 270156 218204 270162
rect 218152 270098 218204 270104
rect 218164 264316 218192 270098
rect 218348 268122 218376 277780
rect 219164 272604 219216 272610
rect 219164 272546 219216 272552
rect 218612 272536 218664 272542
rect 218612 272478 218664 272484
rect 218336 268116 218388 268122
rect 218336 268058 218388 268064
rect 218624 264316 218652 272478
rect 219072 270360 219124 270366
rect 219072 270302 219124 270308
rect 219084 264316 219112 270302
rect 219176 264330 219204 272546
rect 219544 270298 219572 277780
rect 220360 272672 220412 272678
rect 220360 272614 220412 272620
rect 219992 270428 220044 270434
rect 219992 270370 220044 270376
rect 219532 270292 219584 270298
rect 219532 270234 219584 270240
rect 219176 264302 219558 264330
rect 220004 264316 220032 270370
rect 220372 264316 220400 272614
rect 220740 270094 220768 277780
rect 221280 272876 221332 272882
rect 221280 272818 221332 272824
rect 220820 270496 220872 270502
rect 220820 270438 220872 270444
rect 220728 270088 220780 270094
rect 220728 270030 220780 270036
rect 220832 264316 220860 270438
rect 221292 264316 221320 272818
rect 221936 270434 221964 277780
rect 222200 272808 222252 272814
rect 222200 272750 222252 272756
rect 221924 270428 221976 270434
rect 221924 270370 221976 270376
rect 221738 268696 221794 268705
rect 221738 268631 221794 268640
rect 221752 264316 221780 268631
rect 222212 264316 222240 272750
rect 223028 272740 223080 272746
rect 223028 272682 223080 272688
rect 222660 268048 222712 268054
rect 222660 267990 222712 267996
rect 222672 264316 222700 267990
rect 223040 264316 223068 272682
rect 223132 270162 223160 277780
rect 223488 273080 223540 273086
rect 223488 273022 223540 273028
rect 223120 270156 223172 270162
rect 223120 270098 223172 270104
rect 223500 264316 223528 273022
rect 223948 272944 224000 272950
rect 223948 272886 224000 272892
rect 223764 268864 223816 268870
rect 223764 268806 223816 268812
rect 223580 268660 223632 268666
rect 223580 268602 223632 268608
rect 223592 268410 223620 268602
rect 223592 268382 223712 268410
rect 223684 268326 223712 268382
rect 223580 268320 223632 268326
rect 223580 268262 223632 268268
rect 223672 268320 223724 268326
rect 223672 268262 223724 268268
rect 223592 268122 223620 268262
rect 223580 268116 223632 268122
rect 223580 268058 223632 268064
rect 223776 267850 223804 268806
rect 223764 267844 223816 267850
rect 223764 267786 223816 267792
rect 223960 264316 223988 272886
rect 224236 270366 224264 277780
rect 224408 273012 224460 273018
rect 224408 272954 224460 272960
rect 224224 270360 224276 270366
rect 224224 270302 224276 270308
rect 224132 269680 224184 269686
rect 224132 269622 224184 269628
rect 224144 269006 224172 269622
rect 224040 269000 224092 269006
rect 224040 268942 224092 268948
rect 224132 269000 224184 269006
rect 224132 268942 224184 268948
rect 224052 268802 224080 268942
rect 224040 268796 224092 268802
rect 224040 268738 224092 268744
rect 224420 264316 224448 272954
rect 225432 270502 225460 277780
rect 226156 273216 226208 273222
rect 226156 273158 226208 273164
rect 225420 270496 225472 270502
rect 225420 270438 225472 270444
rect 225328 269068 225380 269074
rect 225328 269010 225380 269016
rect 224868 267912 224920 267918
rect 224868 267854 224920 267860
rect 224880 264316 224908 267854
rect 225340 264316 225368 269010
rect 225786 268560 225842 268569
rect 225786 268495 225842 268504
rect 225800 264316 225828 268495
rect 226168 264316 226196 273158
rect 226340 271720 226392 271726
rect 226340 271662 226392 271668
rect 226352 264330 226380 271662
rect 226628 270570 226656 277780
rect 227076 273148 227128 273154
rect 227076 273090 227128 273096
rect 226616 270564 226668 270570
rect 226616 270506 226668 270512
rect 226352 264302 226642 264330
rect 227088 264316 227116 273090
rect 227628 271040 227680 271046
rect 227628 270982 227680 270988
rect 227536 268796 227588 268802
rect 227536 268738 227588 268744
rect 227548 264316 227576 268738
rect 227640 267782 227668 270982
rect 227824 270638 227852 277780
rect 229020 271726 229048 277780
rect 230216 272542 230244 277780
rect 230204 272536 230256 272542
rect 230204 272478 230256 272484
rect 229008 271720 229060 271726
rect 229008 271662 229060 271668
rect 231412 271658 231440 277780
rect 232516 272746 232544 277780
rect 232504 272740 232556 272746
rect 232504 272682 232556 272688
rect 233712 272610 233740 277780
rect 234908 272814 234936 277780
rect 236104 272882 236132 277780
rect 236092 272876 236144 272882
rect 236092 272818 236144 272824
rect 234896 272808 234948 272814
rect 234896 272750 234948 272756
rect 237300 272678 237328 277780
rect 237288 272672 237340 272678
rect 237288 272614 237340 272620
rect 233700 272604 233752 272610
rect 233700 272546 233752 272552
rect 238496 272202 238524 277780
rect 239600 272950 239628 277780
rect 239588 272944 239640 272950
rect 239588 272886 239640 272892
rect 234620 272196 234672 272202
rect 234620 272138 234672 272144
rect 238484 272196 238536 272202
rect 238484 272138 238536 272144
rect 229284 271652 229336 271658
rect 229284 271594 229336 271600
rect 231400 271652 231452 271658
rect 231400 271594 231452 271600
rect 228824 271516 228876 271522
rect 228824 271458 228876 271464
rect 227812 270632 227864 270638
rect 227812 270574 227864 270580
rect 228456 268864 228508 268870
rect 228456 268806 228508 268812
rect 227996 267844 228048 267850
rect 227996 267786 228048 267792
rect 227628 267776 227680 267782
rect 227628 267718 227680 267724
rect 228008 264316 228036 267786
rect 228468 264316 228496 268806
rect 228836 264316 228864 271458
rect 229100 270700 229152 270706
rect 229100 270642 229152 270648
rect 229112 268870 229140 270642
rect 229100 268864 229152 268870
rect 229100 268806 229152 268812
rect 229296 264316 229324 271594
rect 229744 271584 229796 271590
rect 229744 271526 229796 271532
rect 229756 264316 229784 271526
rect 232412 271448 232464 271454
rect 232412 271390 232464 271396
rect 231492 271380 231544 271386
rect 231492 271322 231544 271328
rect 230756 270768 230808 270774
rect 230756 270710 230808 270716
rect 230204 268728 230256 268734
rect 230204 268670 230256 268676
rect 230216 264316 230244 268670
rect 230768 268598 230796 270710
rect 231124 268660 231176 268666
rect 231124 268602 231176 268608
rect 230664 268592 230716 268598
rect 230664 268534 230716 268540
rect 230756 268592 230808 268598
rect 230756 268534 230808 268540
rect 230676 264316 230704 268534
rect 231136 264316 231164 268602
rect 231504 264316 231532 271322
rect 231768 271312 231820 271318
rect 231768 271254 231820 271260
rect 231780 267764 231808 271254
rect 231860 270836 231912 270842
rect 231860 270778 231912 270784
rect 231872 268938 231900 270778
rect 231860 268932 231912 268938
rect 231860 268874 231912 268880
rect 231780 267736 231900 267764
rect 231872 264330 231900 267736
rect 231872 264302 231978 264330
rect 232424 264316 232452 271390
rect 232688 271244 232740 271250
rect 232688 271186 232740 271192
rect 232700 267850 232728 271186
rect 234528 271176 234580 271182
rect 234528 271118 234580 271124
rect 232964 271108 233016 271114
rect 232964 271050 233016 271056
rect 232976 268326 233004 271050
rect 233424 270904 233476 270910
rect 233424 270846 233476 270852
rect 233436 268394 233464 270846
rect 233792 268456 233844 268462
rect 233792 268398 233844 268404
rect 233332 268388 233384 268394
rect 233332 268330 233384 268336
rect 233424 268388 233476 268394
rect 233424 268330 233476 268336
rect 232872 268320 232924 268326
rect 232872 268262 232924 268268
rect 232964 268320 233016 268326
rect 232964 268262 233016 268268
rect 232688 267844 232740 267850
rect 232688 267786 232740 267792
rect 232884 264316 232912 268262
rect 233344 264316 233372 268330
rect 233804 264316 233832 268398
rect 234160 267776 234212 267782
rect 234540 267764 234568 271118
rect 234632 269686 234660 272138
rect 240140 272128 240192 272134
rect 240140 272070 240192 272076
rect 234712 270972 234764 270978
rect 234712 270914 234764 270920
rect 234620 269680 234672 269686
rect 234620 269622 234672 269628
rect 234724 267782 234752 270914
rect 239128 269680 239180 269686
rect 239128 269622 239180 269628
rect 238668 268932 238720 268938
rect 238668 268874 238720 268880
rect 236644 268592 236696 268598
rect 236644 268534 236696 268540
rect 236000 268320 236052 268326
rect 236000 268262 236052 268268
rect 235540 268252 235592 268258
rect 235540 268194 235592 268200
rect 235080 267844 235132 267850
rect 235080 267786 235132 267792
rect 234712 267776 234764 267782
rect 234540 267736 234660 267764
rect 234160 267718 234212 267724
rect 234172 264316 234200 267718
rect 234632 264316 234660 267736
rect 234712 267718 234764 267724
rect 235092 264316 235120 267786
rect 235552 264316 235580 268194
rect 236012 264316 236040 268262
rect 236460 268116 236512 268122
rect 236460 268058 236512 268064
rect 236472 264316 236500 268058
rect 236656 268054 236684 268534
rect 237288 268388 237340 268394
rect 237288 268330 237340 268336
rect 236920 268184 236972 268190
rect 236920 268126 236972 268132
rect 236644 268048 236696 268054
rect 236644 267990 236696 267996
rect 236932 264316 236960 268126
rect 237300 264316 237328 268330
rect 238208 268048 238260 268054
rect 238208 267990 238260 267996
rect 237748 267776 237800 267782
rect 237748 267718 237800 267724
rect 237760 264316 237788 267718
rect 238220 264316 238248 267990
rect 238680 264316 238708 268874
rect 239140 264316 239168 269622
rect 239956 269408 240008 269414
rect 239956 269350 240008 269356
rect 239588 268864 239640 268870
rect 239588 268806 239640 268812
rect 239600 264316 239628 268806
rect 239968 264316 239996 269350
rect 240152 268598 240180 272070
rect 240796 271794 240824 277780
rect 241992 273018 242020 277780
rect 243188 273086 243216 277780
rect 243176 273080 243228 273086
rect 243176 273022 243228 273028
rect 241980 273012 242032 273018
rect 241980 272954 242032 272960
rect 242624 272060 242676 272066
rect 242624 272002 242676 272008
rect 242256 271924 242308 271930
rect 242256 271866 242308 271872
rect 240876 271856 240928 271862
rect 240876 271798 240928 271804
rect 240784 271788 240836 271794
rect 240784 271730 240836 271736
rect 240416 269136 240468 269142
rect 240416 269078 240468 269084
rect 240140 268592 240192 268598
rect 240140 268534 240192 268540
rect 240428 264316 240456 269078
rect 240888 264316 240916 271798
rect 241796 269340 241848 269346
rect 241796 269282 241848 269288
rect 241336 269204 241388 269210
rect 241336 269146 241388 269152
rect 241348 264316 241376 269146
rect 241808 264316 241836 269282
rect 242268 264316 242296 271866
rect 242636 264316 242664 272002
rect 243544 271992 243596 271998
rect 243544 271934 243596 271940
rect 243084 269272 243136 269278
rect 243084 269214 243136 269220
rect 243096 264316 243124 269214
rect 243556 264316 243584 271934
rect 244384 271930 244412 277780
rect 244372 271924 244424 271930
rect 244372 271866 244424 271872
rect 245580 271862 245608 277780
rect 245568 271856 245620 271862
rect 245568 271798 245620 271804
rect 246776 271046 246804 277780
rect 247880 271182 247908 277780
rect 249076 271590 249104 277780
rect 249064 271584 249116 271590
rect 249064 271526 249116 271532
rect 247868 271176 247920 271182
rect 247868 271118 247920 271124
rect 246764 271040 246816 271046
rect 246764 270982 246816 270988
rect 250272 270978 250300 277780
rect 251468 271250 251496 277780
rect 252664 271522 252692 277780
rect 253756 271720 253808 271726
rect 253756 271662 253808 271668
rect 252652 271516 252704 271522
rect 252652 271458 252704 271464
rect 251456 271244 251508 271250
rect 251456 271186 251508 271192
rect 250260 270972 250312 270978
rect 250260 270914 250312 270920
rect 253388 270632 253440 270638
rect 253388 270574 253440 270580
rect 252928 270564 252980 270570
rect 252928 270506 252980 270512
rect 252468 270496 252520 270502
rect 252468 270438 252520 270444
rect 251088 270428 251140 270434
rect 251088 270370 251140 270376
rect 250260 270292 250312 270298
rect 250260 270234 250312 270240
rect 249340 270224 249392 270230
rect 249340 270166 249392 270172
rect 248880 270020 248932 270026
rect 248880 269962 248932 269968
rect 248420 269952 248472 269958
rect 248420 269894 248472 269900
rect 246672 269884 246724 269890
rect 246672 269826 246724 269832
rect 245752 269748 245804 269754
rect 245752 269690 245804 269696
rect 244464 269544 244516 269550
rect 244464 269486 244516 269492
rect 244004 269476 244056 269482
rect 244004 269418 244056 269424
rect 244016 264316 244044 269418
rect 244476 264316 244504 269486
rect 245292 269000 245344 269006
rect 245292 268942 245344 268948
rect 244924 268592 244976 268598
rect 244924 268534 244976 268540
rect 244936 264316 244964 268534
rect 245304 264316 245332 268942
rect 245764 264316 245792 269690
rect 246212 269612 246264 269618
rect 246212 269554 246264 269560
rect 246224 264316 246252 269554
rect 246684 264316 246712 269826
rect 247592 269816 247644 269822
rect 247592 269758 247644 269764
rect 247132 267980 247184 267986
rect 247132 267922 247184 267928
rect 247144 264316 247172 267922
rect 247604 264316 247632 269758
rect 248052 268524 248104 268530
rect 248052 268466 248104 268472
rect 248064 264316 248092 268466
rect 248432 264316 248460 269894
rect 248892 264316 248920 269962
rect 249352 264316 249380 270166
rect 249800 268116 249852 268122
rect 249800 268058 249852 268064
rect 249812 264316 249840 268058
rect 250272 264316 250300 270234
rect 250720 270088 250772 270094
rect 250720 270030 250772 270036
rect 250732 264316 250760 270030
rect 251100 264316 251128 270370
rect 252008 270360 252060 270366
rect 252008 270302 252060 270308
rect 251548 270156 251600 270162
rect 251548 270098 251600 270104
rect 251560 264316 251588 270098
rect 252020 264316 252048 270302
rect 252480 264316 252508 270438
rect 252940 264316 252968 270506
rect 253400 264316 253428 270574
rect 253768 264316 253796 271662
rect 253860 271114 253888 277780
rect 254216 272536 254268 272542
rect 254216 272478 254268 272484
rect 253848 271108 253900 271114
rect 253848 271050 253900 271056
rect 254228 264316 254256 272478
rect 254676 271652 254728 271658
rect 254676 271594 254728 271600
rect 254688 264316 254716 271594
rect 255056 271318 255084 277780
rect 256056 272808 256108 272814
rect 256056 272750 256108 272756
rect 255136 272740 255188 272746
rect 255136 272682 255188 272688
rect 255044 271312 255096 271318
rect 255044 271254 255096 271260
rect 255148 264316 255176 272682
rect 255596 272604 255648 272610
rect 255596 272546 255648 272552
rect 255608 264316 255636 272546
rect 256068 264316 256096 272750
rect 256160 271386 256188 277780
rect 256424 272876 256476 272882
rect 256424 272818 256476 272824
rect 256148 271380 256200 271386
rect 256148 271322 256200 271328
rect 256436 264316 256464 272818
rect 257160 272672 257212 272678
rect 257160 272614 257212 272620
rect 257172 264330 257200 272614
rect 257252 272196 257304 272202
rect 257252 272138 257304 272144
rect 257264 270586 257292 272138
rect 257356 270706 257384 277780
rect 257804 272944 257856 272950
rect 257804 272886 257856 272892
rect 257344 270700 257396 270706
rect 257344 270642 257396 270648
rect 257264 270558 257384 270586
rect 256910 264302 257200 264330
rect 257356 264316 257384 270558
rect 257816 264316 257844 272886
rect 258264 271788 258316 271794
rect 258264 271730 258316 271736
rect 258276 264316 258304 271730
rect 258552 271454 258580 277780
rect 259184 273080 259236 273086
rect 259184 273022 259236 273028
rect 258724 273012 258776 273018
rect 258724 272954 258776 272960
rect 258540 271448 258592 271454
rect 258540 271390 258592 271396
rect 258736 264316 258764 272954
rect 259196 264316 259224 273022
rect 259552 271924 259604 271930
rect 259552 271866 259604 271872
rect 259564 264316 259592 271866
rect 259748 270842 259776 277780
rect 260944 273086 260972 277780
rect 260932 273080 260984 273086
rect 260932 273022 260984 273028
rect 260012 271856 260064 271862
rect 260012 271798 260064 271804
rect 259736 270836 259788 270842
rect 259736 270778 259788 270784
rect 260024 264316 260052 271798
rect 262140 271794 262168 277780
rect 263244 273222 263272 277780
rect 263232 273216 263284 273222
rect 263232 273158 263284 273164
rect 264440 273154 264468 277780
rect 264428 273148 264480 273154
rect 264428 273090 264480 273096
rect 262128 271788 262180 271794
rect 262128 271730 262180 271736
rect 261392 271584 261444 271590
rect 261392 271526 261444 271532
rect 260932 271176 260984 271182
rect 260932 271118 260984 271124
rect 260472 271040 260524 271046
rect 260472 270982 260524 270988
rect 260484 264316 260512 270982
rect 260944 264316 260972 271118
rect 261404 264316 261432 271526
rect 262864 271516 262916 271522
rect 262864 271458 262916 271464
rect 262220 271244 262272 271250
rect 262220 271186 262272 271192
rect 261852 270972 261904 270978
rect 261852 270914 261904 270920
rect 261864 264316 261892 270914
rect 262232 264316 262260 271186
rect 262876 264330 262904 271458
rect 264888 271448 264940 271454
rect 264888 271390 264940 271396
rect 264060 271380 264112 271386
rect 264060 271322 264112 271328
rect 263600 271312 263652 271318
rect 263600 271254 263652 271260
rect 263140 271108 263192 271114
rect 263140 271050 263192 271056
rect 262706 264302 262904 264330
rect 263152 264316 263180 271050
rect 263612 264316 263640 271254
rect 264072 264316 264100 271322
rect 264520 270700 264572 270706
rect 264520 270642 264572 270648
rect 264532 264316 264560 270642
rect 264900 264316 264928 271390
rect 265440 270836 265492 270842
rect 265440 270778 265492 270784
rect 265452 264330 265480 270778
rect 265636 270502 265664 277780
rect 266728 273216 266780 273222
rect 266728 273158 266780 273164
rect 265808 273080 265860 273086
rect 265808 273022 265860 273028
rect 265624 270496 265676 270502
rect 265624 270438 265676 270444
rect 265374 264302 265480 264330
rect 265820 264316 265848 273022
rect 266268 271788 266320 271794
rect 266268 271730 266320 271736
rect 266280 264316 266308 271730
rect 266740 264316 266768 273158
rect 266832 271250 266860 277780
rect 268042 277766 268516 277794
rect 267188 273148 267240 273154
rect 267188 273090 267240 273096
rect 266820 271244 266872 271250
rect 266820 271186 266872 271192
rect 267200 264316 267228 273090
rect 268016 271244 268068 271250
rect 268016 271186 268068 271192
rect 267556 270496 267608 270502
rect 267556 270438 267608 270444
rect 267568 264316 267596 270438
rect 268028 264316 268056 271186
rect 268488 264316 268516 277766
rect 268948 277766 269238 277794
rect 268948 264316 268976 277766
rect 269856 270496 269908 270502
rect 269856 270438 269908 270444
rect 269396 269136 269448 269142
rect 269396 269078 269448 269084
rect 269408 264316 269436 269078
rect 269868 264316 269896 270438
rect 270316 270428 270368 270434
rect 270316 270370 270368 270376
rect 270328 264316 270356 270370
rect 270420 269142 270448 277780
rect 271524 270502 271552 277780
rect 271512 270496 271564 270502
rect 271512 270438 271564 270444
rect 272064 270496 272116 270502
rect 272064 270438 272116 270444
rect 271144 270360 271196 270366
rect 271144 270302 271196 270308
rect 270408 269136 270460 269142
rect 270408 269078 270460 269084
rect 270684 268252 270736 268258
rect 270684 268194 270736 268200
rect 270696 264316 270724 268194
rect 271156 264316 271184 270302
rect 271604 268048 271656 268054
rect 271604 267990 271656 267996
rect 271616 264316 271644 267990
rect 272076 264316 272104 270438
rect 272720 270434 272748 277780
rect 272708 270428 272760 270434
rect 272708 270370 272760 270376
rect 273720 270428 273772 270434
rect 273720 270370 273772 270376
rect 272984 268864 273036 268870
rect 272984 268806 273036 268812
rect 272524 268456 272576 268462
rect 272524 268398 272576 268404
rect 272536 264316 272564 268398
rect 272996 264316 273024 268806
rect 273732 264330 273760 270370
rect 273812 268728 273864 268734
rect 273812 268670 273864 268676
rect 273378 264302 273760 264330
rect 273824 264316 273852 268670
rect 273916 268258 273944 277780
rect 275112 270366 275140 277780
rect 275100 270360 275152 270366
rect 275100 270302 275152 270308
rect 274272 270292 274324 270298
rect 274272 270234 274324 270240
rect 273904 268252 273956 268258
rect 273904 268194 273956 268200
rect 274284 264316 274312 270234
rect 274732 269884 274784 269890
rect 274732 269826 274784 269832
rect 274744 264316 274772 269826
rect 275192 268320 275244 268326
rect 275192 268262 275244 268268
rect 275204 264316 275232 268262
rect 275652 268252 275704 268258
rect 275652 268194 275704 268200
rect 275664 264316 275692 268194
rect 276308 268054 276336 277780
rect 277504 270502 277532 277780
rect 277492 270496 277544 270502
rect 277492 270438 277544 270444
rect 277400 270360 277452 270366
rect 277400 270302 277452 270308
rect 276940 269340 276992 269346
rect 276940 269282 276992 269288
rect 276296 268048 276348 268054
rect 276296 267990 276348 267996
rect 276388 268048 276440 268054
rect 276388 267990 276440 267996
rect 276400 264330 276428 267990
rect 276480 267912 276532 267918
rect 276480 267854 276532 267860
rect 276046 264302 276428 264330
rect 276492 264316 276520 267854
rect 276952 264316 276980 269282
rect 277412 264316 277440 270302
rect 277860 270224 277912 270230
rect 277860 270166 277912 270172
rect 277872 264316 277900 270166
rect 278596 270156 278648 270162
rect 278596 270098 278648 270104
rect 278320 270088 278372 270094
rect 278320 270030 278372 270036
rect 278332 264316 278360 270030
rect 278608 264330 278636 270098
rect 278700 268462 278728 277780
rect 279148 270020 279200 270026
rect 279148 269962 279200 269968
rect 278688 268456 278740 268462
rect 278688 268398 278740 268404
rect 278608 264302 278714 264330
rect 279160 264316 279188 269962
rect 279608 269952 279660 269958
rect 279608 269894 279660 269900
rect 279620 264316 279648 269894
rect 279804 268870 279832 277780
rect 281000 270434 281028 277780
rect 280988 270428 281040 270434
rect 280988 270370 281040 270376
rect 280528 269816 280580 269822
rect 280528 269758 280580 269764
rect 280068 269748 280120 269754
rect 280068 269690 280120 269696
rect 279792 268864 279844 268870
rect 279792 268806 279844 268812
rect 280080 264316 280108 269690
rect 280540 264316 280568 269758
rect 281816 269680 281868 269686
rect 281816 269622 281868 269628
rect 281448 269612 281500 269618
rect 281448 269554 281500 269560
rect 280988 269544 281040 269550
rect 280988 269486 281040 269492
rect 281000 264316 281028 269486
rect 281460 264316 281488 269554
rect 281828 264316 281856 269622
rect 282196 268734 282224 277780
rect 283392 270298 283420 277780
rect 284208 272060 284260 272066
rect 284208 272002 284260 272008
rect 283380 270292 283432 270298
rect 283380 270234 283432 270240
rect 283472 270292 283524 270298
rect 283472 270234 283524 270240
rect 282736 269476 282788 269482
rect 282736 269418 282788 269424
rect 282276 269408 282328 269414
rect 282276 269350 282328 269356
rect 282184 268728 282236 268734
rect 282184 268670 282236 268676
rect 282288 264316 282316 269350
rect 282748 264316 282776 269418
rect 283484 269346 283512 270234
rect 283472 269340 283524 269346
rect 283472 269282 283524 269288
rect 283656 269340 283708 269346
rect 283656 269282 283708 269288
rect 283196 269272 283248 269278
rect 283196 269214 283248 269220
rect 283208 264316 283236 269214
rect 283668 264316 283696 269282
rect 284220 264330 284248 272002
rect 284588 269890 284616 277780
rect 285404 271992 285456 271998
rect 285404 271934 285456 271940
rect 284576 269884 284628 269890
rect 284576 269826 284628 269832
rect 284944 269204 284996 269210
rect 284944 269146 284996 269152
rect 284484 269136 284536 269142
rect 284484 269078 284536 269084
rect 284142 264302 284248 264330
rect 284496 264316 284524 269078
rect 284956 264316 284984 269146
rect 285416 264316 285444 271934
rect 285784 268326 285812 277780
rect 286600 271380 286652 271386
rect 286600 271322 286652 271328
rect 285864 271040 285916 271046
rect 285864 270982 285916 270988
rect 285772 268320 285824 268326
rect 285772 268262 285824 268268
rect 285876 264316 285904 270982
rect 286612 264330 286640 271322
rect 286692 271176 286744 271182
rect 286692 271118 286744 271124
rect 286350 264302 286640 264330
rect 286704 264330 286732 271118
rect 286888 268258 286916 277780
rect 287612 271312 287664 271318
rect 287612 271254 287664 271260
rect 287152 271244 287204 271250
rect 287152 271186 287204 271192
rect 286876 268252 286928 268258
rect 286876 268194 286928 268200
rect 286704 264302 286810 264330
rect 287164 264316 287192 271186
rect 287624 264316 287652 271254
rect 288084 268054 288112 277780
rect 288992 271516 289044 271522
rect 288992 271458 289044 271464
rect 288532 271448 288584 271454
rect 288532 271390 288584 271396
rect 288164 271108 288216 271114
rect 288164 271050 288216 271056
rect 288072 268048 288124 268054
rect 288072 267990 288124 267996
rect 288176 264330 288204 271050
rect 288098 264302 288204 264330
rect 288544 264316 288572 271390
rect 289004 264316 289032 271458
rect 289280 267918 289308 277780
rect 290280 271924 290332 271930
rect 290280 271866 290332 271872
rect 289360 271856 289412 271862
rect 289360 271798 289412 271804
rect 289268 267912 289320 267918
rect 289268 267854 289320 267860
rect 289372 264330 289400 271798
rect 289820 271652 289872 271658
rect 289820 271594 289872 271600
rect 289372 264302 289478 264330
rect 289832 264316 289860 271594
rect 290292 264316 290320 271866
rect 290476 270298 290504 277780
rect 290740 271720 290792 271726
rect 290740 271662 290792 271668
rect 290464 270292 290516 270298
rect 290464 270234 290516 270240
rect 290752 264316 290780 271662
rect 291200 271584 291252 271590
rect 291200 271526 291252 271532
rect 291212 264316 291240 271526
rect 291672 270366 291700 277780
rect 292028 273216 292080 273222
rect 292028 273158 292080 273164
rect 291660 270360 291712 270366
rect 291660 270302 291712 270308
rect 292040 264330 292068 273158
rect 292580 273148 292632 273154
rect 292580 273090 292632 273096
rect 292488 271788 292540 271794
rect 292488 271730 292540 271736
rect 292500 264330 292528 271730
rect 291686 264302 292068 264330
rect 292146 264302 292528 264330
rect 292592 264316 292620 273090
rect 292868 270230 292896 277780
rect 293868 273080 293920 273086
rect 293868 273022 293920 273028
rect 293408 273012 293460 273018
rect 293408 272954 293460 272960
rect 292856 270224 292908 270230
rect 292856 270166 292908 270172
rect 292948 269068 293000 269074
rect 292948 269010 293000 269016
rect 292960 264316 292988 269010
rect 293420 264316 293448 272954
rect 293880 264316 293908 273022
rect 294064 270094 294092 277780
rect 294880 272740 294932 272746
rect 294880 272682 294932 272688
rect 294788 272332 294840 272338
rect 294788 272274 294840 272280
rect 294328 270428 294380 270434
rect 294328 270370 294380 270376
rect 294052 270088 294104 270094
rect 294052 270030 294104 270036
rect 294340 264316 294368 270370
rect 294800 264316 294828 272274
rect 294892 264330 294920 272682
rect 295168 270162 295196 277780
rect 296076 272536 296128 272542
rect 296076 272478 296128 272484
rect 295156 270156 295208 270162
rect 295156 270098 295208 270104
rect 295616 269000 295668 269006
rect 295616 268942 295668 268948
rect 294892 264302 295274 264330
rect 295628 264316 295656 268942
rect 296088 264316 296116 272478
rect 296364 270026 296392 277780
rect 296996 270360 297048 270366
rect 296996 270302 297048 270308
rect 296536 270224 296588 270230
rect 296536 270166 296588 270172
rect 296352 270020 296404 270026
rect 296352 269962 296404 269968
rect 296548 264316 296576 270166
rect 297008 264316 297036 270302
rect 297456 270292 297508 270298
rect 297456 270234 297508 270240
rect 297468 264316 297496 270234
rect 297560 269958 297588 277780
rect 298284 270156 298336 270162
rect 298284 270098 298336 270104
rect 297548 269952 297600 269958
rect 297548 269894 297600 269900
rect 297916 267980 297968 267986
rect 297916 267922 297968 267928
rect 297928 264316 297956 267922
rect 298296 264316 298324 270098
rect 298756 269754 298784 277780
rect 299204 270088 299256 270094
rect 299204 270030 299256 270036
rect 298744 269748 298796 269754
rect 298744 269690 298796 269696
rect 298744 268048 298796 268054
rect 298744 267990 298796 267996
rect 298756 264316 298784 267990
rect 299216 264316 299244 270030
rect 299952 269822 299980 277780
rect 300768 272808 300820 272814
rect 300768 272750 300820 272756
rect 300676 272604 300728 272610
rect 300676 272546 300728 272552
rect 299940 269816 299992 269822
rect 299940 269758 299992 269764
rect 299664 267164 299716 267170
rect 299664 267106 299716 267112
rect 299676 264316 299704 267106
rect 300688 264974 300716 272546
rect 300504 264946 300716 264974
rect 300504 264330 300532 264946
rect 300780 264330 300808 272750
rect 301148 269550 301176 277780
rect 301412 272672 301464 272678
rect 301412 272614 301464 272620
rect 301136 269544 301188 269550
rect 301136 269486 301188 269492
rect 300952 267096 301004 267102
rect 300952 267038 301004 267044
rect 300150 264302 300532 264330
rect 300610 264302 300808 264330
rect 300964 264316 300992 267038
rect 301424 264316 301452 272614
rect 301872 272468 301924 272474
rect 301872 272410 301924 272416
rect 301884 264316 301912 272410
rect 302344 269618 302372 277780
rect 303344 272400 303396 272406
rect 303344 272342 303396 272348
rect 302792 272264 302844 272270
rect 302792 272206 302844 272212
rect 302332 269612 302384 269618
rect 302332 269554 302384 269560
rect 302332 267028 302384 267034
rect 302332 266970 302384 266976
rect 302344 264316 302372 266970
rect 302804 264316 302832 272206
rect 303356 264330 303384 272342
rect 303448 269686 303476 277780
rect 304080 270496 304132 270502
rect 304080 270438 304132 270444
rect 303436 269680 303488 269686
rect 303436 269622 303488 269628
rect 303712 266960 303764 266966
rect 303712 266902 303764 266908
rect 303278 264302 303384 264330
rect 303724 264316 303752 266902
rect 304092 264316 304120 270438
rect 304644 269414 304672 277780
rect 304908 272944 304960 272950
rect 304908 272886 304960 272892
rect 304632 269408 304684 269414
rect 304632 269350 304684 269356
rect 304920 267986 304948 272886
rect 305460 269952 305512 269958
rect 305460 269894 305512 269900
rect 304908 267980 304960 267986
rect 304908 267922 304960 267928
rect 304540 267844 304592 267850
rect 304540 267786 304592 267792
rect 304552 264316 304580 267786
rect 305000 266892 305052 266898
rect 305000 266834 305052 266840
rect 305012 264316 305040 266834
rect 305472 264316 305500 269894
rect 305840 269482 305868 277780
rect 306288 272196 306340 272202
rect 306288 272138 306340 272144
rect 305828 269476 305880 269482
rect 305828 269418 305880 269424
rect 306300 264330 306328 272138
rect 306748 269884 306800 269890
rect 306748 269826 306800 269832
rect 306380 266824 306432 266830
rect 306380 266766 306432 266772
rect 305946 264302 306328 264330
rect 306392 264316 306420 266766
rect 306760 264316 306788 269826
rect 307036 269278 307064 277780
rect 307852 272876 307904 272882
rect 307852 272818 307904 272824
rect 307208 269816 307260 269822
rect 307208 269758 307260 269764
rect 307024 269272 307076 269278
rect 307024 269214 307076 269220
rect 307220 264316 307248 269758
rect 307864 268054 307892 272818
rect 308128 269748 308180 269754
rect 308128 269690 308180 269696
rect 307852 268048 307904 268054
rect 307852 267990 307904 267996
rect 307668 266756 307720 266762
rect 307668 266698 307720 266704
rect 307680 264316 307708 266698
rect 308140 264316 308168 269690
rect 308232 269346 308260 277780
rect 308956 272128 309008 272134
rect 308956 272070 309008 272076
rect 308220 269340 308272 269346
rect 308220 269282 308272 269288
rect 308968 264330 308996 272070
rect 309428 272066 309456 277780
rect 309416 272060 309468 272066
rect 309416 272002 309468 272008
rect 310532 269142 310560 277780
rect 311624 272060 311676 272066
rect 311624 272002 311676 272008
rect 310796 269612 310848 269618
rect 310796 269554 310848 269560
rect 310520 269136 310572 269142
rect 310520 269078 310572 269084
rect 309876 268932 309928 268938
rect 309876 268874 309928 268880
rect 309416 268388 309468 268394
rect 309416 268330 309468 268336
rect 309048 266688 309100 266694
rect 309048 266630 309100 266636
rect 308614 264302 308996 264330
rect 309060 264316 309088 266630
rect 309428 264316 309456 268330
rect 309888 264316 309916 268874
rect 310336 266620 310388 266626
rect 310336 266562 310388 266568
rect 310348 264316 310376 266562
rect 310808 264316 310836 269554
rect 311636 264330 311664 272002
rect 311728 269210 311756 277780
rect 312924 271998 312952 277780
rect 312912 271992 312964 271998
rect 312912 271934 312964 271940
rect 314120 271046 314148 277780
rect 314292 271992 314344 271998
rect 314292 271934 314344 271940
rect 314108 271040 314160 271046
rect 314108 270982 314160 270988
rect 312084 269544 312136 269550
rect 312084 269486 312136 269492
rect 311716 269204 311768 269210
rect 311716 269146 311768 269152
rect 311716 266552 311768 266558
rect 311716 266494 311768 266500
rect 311282 264302 311664 264330
rect 311728 264316 311756 266494
rect 312096 264316 312124 269486
rect 313464 269476 313516 269482
rect 313464 269418 313516 269424
rect 312544 268320 312596 268326
rect 312544 268262 312596 268268
rect 312556 264316 312584 268262
rect 313004 266484 313056 266490
rect 313004 266426 313056 266432
rect 313016 264316 313044 266426
rect 313476 264316 313504 269418
rect 314304 264330 314332 271934
rect 315316 271386 315344 277780
rect 315304 271380 315356 271386
rect 315304 271322 315356 271328
rect 316512 271182 316540 277780
rect 317708 271250 317736 277780
rect 318812 271318 318840 277780
rect 318892 274848 318944 274854
rect 318892 274790 318944 274796
rect 318800 271312 318852 271318
rect 318800 271254 318852 271260
rect 317696 271244 317748 271250
rect 317696 271186 317748 271192
rect 316500 271176 316552 271182
rect 316500 271118 316552 271124
rect 314844 269408 314896 269414
rect 314844 269350 314896 269356
rect 314384 265260 314436 265266
rect 314384 265202 314436 265208
rect 313950 264302 314332 264330
rect 314396 264316 314424 265202
rect 314856 264316 314884 269350
rect 315212 269340 315264 269346
rect 315212 269282 315264 269288
rect 315224 264316 315252 269282
rect 317880 269272 317932 269278
rect 317880 269214 317932 269220
rect 316132 268252 316184 268258
rect 316132 268194 316184 268200
rect 315672 266416 315724 266422
rect 315672 266358 315724 266364
rect 315684 264316 315712 266358
rect 316144 264316 316172 268194
rect 316592 268184 316644 268190
rect 316592 268126 316644 268132
rect 316604 264316 316632 268126
rect 317052 266348 317104 266354
rect 317052 266290 317104 266296
rect 317064 264316 317092 266290
rect 317512 265804 317564 265810
rect 317512 265746 317564 265752
rect 317524 264316 317552 265746
rect 317892 264316 317920 269214
rect 318340 265328 318392 265334
rect 318340 265270 318392 265276
rect 318352 264316 318380 265270
rect 318904 264330 318932 274790
rect 320008 271114 320036 277780
rect 320180 274780 320232 274786
rect 320180 274722 320232 274728
rect 319996 271108 320048 271114
rect 319996 271050 320048 271056
rect 319260 268048 319312 268054
rect 319260 267990 319312 267996
rect 318826 264302 318932 264330
rect 319272 264316 319300 267990
rect 319720 265192 319772 265198
rect 319720 265134 319772 265140
rect 319732 264316 319760 265134
rect 320192 264316 320220 274722
rect 321008 274712 321060 274718
rect 321008 274654 321060 274660
rect 320548 269204 320600 269210
rect 320548 269146 320600 269152
rect 320560 264316 320588 269146
rect 321020 264316 321048 274654
rect 321204 271454 321232 277780
rect 322400 271522 322428 277780
rect 322756 274644 322808 274650
rect 322756 274586 322808 274592
rect 322388 271516 322440 271522
rect 322388 271458 322440 271464
rect 321192 271448 321244 271454
rect 321192 271390 321244 271396
rect 321928 267980 321980 267986
rect 321928 267922 321980 267928
rect 321468 265396 321520 265402
rect 321468 265338 321520 265344
rect 321480 264316 321508 265338
rect 321940 264316 321968 267922
rect 322768 264330 322796 274586
rect 323596 271862 323624 277780
rect 323676 273624 323728 273630
rect 323676 273566 323728 273572
rect 323584 271856 323636 271862
rect 323584 271798 323636 271804
rect 323216 269136 323268 269142
rect 323216 269078 323268 269084
rect 322848 265464 322900 265470
rect 322848 265406 322900 265412
rect 322414 264302 322796 264330
rect 322860 264316 322888 265406
rect 323228 264316 323256 269078
rect 323688 264316 323716 273566
rect 324792 271658 324820 277780
rect 325424 273760 325476 273766
rect 325424 273702 325476 273708
rect 324780 271652 324832 271658
rect 324780 271594 324832 271600
rect 324596 270632 324648 270638
rect 324596 270574 324648 270580
rect 324136 265532 324188 265538
rect 324136 265474 324188 265480
rect 324148 264316 324176 265474
rect 324608 264316 324636 270574
rect 325436 264330 325464 273702
rect 325988 271930 326016 277780
rect 326804 273828 326856 273834
rect 326804 273770 326856 273776
rect 326344 273692 326396 273698
rect 326344 273634 326396 273640
rect 325976 271924 326028 271930
rect 325976 271866 326028 271872
rect 325608 271856 325660 271862
rect 325608 271798 325660 271804
rect 325620 267986 325648 271798
rect 325976 268456 326028 268462
rect 325976 268398 326028 268404
rect 325608 267980 325660 267986
rect 325608 267922 325660 267928
rect 325516 265600 325568 265606
rect 325516 265542 325568 265548
rect 325082 264302 325464 264330
rect 325528 264316 325556 265542
rect 325988 264316 326016 268398
rect 326356 264316 326384 273634
rect 326712 271924 326764 271930
rect 326712 271866 326764 271872
rect 326436 270768 326488 270774
rect 326436 270710 326488 270716
rect 326448 268190 326476 270710
rect 326436 268184 326488 268190
rect 326436 268126 326488 268132
rect 326724 268054 326752 271866
rect 326712 268048 326764 268054
rect 326712 267990 326764 267996
rect 326816 264316 326844 273770
rect 327092 271726 327120 277780
rect 327724 273964 327776 273970
rect 327724 273906 327776 273912
rect 327080 271720 327132 271726
rect 327080 271662 327132 271668
rect 327264 270836 327316 270842
rect 327264 270778 327316 270784
rect 327276 264316 327304 270778
rect 327736 264316 327764 273906
rect 328288 271590 328316 277780
rect 329012 273896 329064 273902
rect 329012 273838 329064 273844
rect 328276 271584 328328 271590
rect 328276 271526 328328 271532
rect 328644 269680 328696 269686
rect 328644 269622 328696 269628
rect 328000 267912 328052 267918
rect 328000 267854 328052 267860
rect 328012 264330 328040 267854
rect 328012 264302 328210 264330
rect 328656 264316 328684 269622
rect 329024 264316 329052 273838
rect 329484 273222 329512 277780
rect 330392 273556 330444 273562
rect 330392 273498 330444 273504
rect 329472 273216 329524 273222
rect 329472 273158 329524 273164
rect 329748 271244 329800 271250
rect 329748 271186 329800 271192
rect 329760 269006 329788 271186
rect 329932 270904 329984 270910
rect 329932 270846 329984 270852
rect 329748 269000 329800 269006
rect 329748 268942 329800 268948
rect 329472 265736 329524 265742
rect 329472 265678 329524 265684
rect 329484 264316 329512 265678
rect 329944 264316 329972 270846
rect 330404 264316 330432 273498
rect 330680 271794 330708 277780
rect 331680 274032 331732 274038
rect 331680 273974 331732 273980
rect 330668 271788 330720 271794
rect 330668 271730 330720 271736
rect 331312 270972 331364 270978
rect 331312 270914 331364 270920
rect 331128 270700 331180 270706
rect 331128 270642 331180 270648
rect 330852 269000 330904 269006
rect 330852 268942 330904 268948
rect 330864 264316 330892 268942
rect 331140 268938 331168 270642
rect 331128 268932 331180 268938
rect 331128 268874 331180 268880
rect 331324 264316 331352 270914
rect 331692 264316 331720 273974
rect 331876 273154 331904 277780
rect 332140 274168 332192 274174
rect 332140 274110 332192 274116
rect 331864 273148 331916 273154
rect 331864 273090 331916 273096
rect 332152 264316 332180 274110
rect 333072 269074 333100 277780
rect 333152 274304 333204 274310
rect 333152 274246 333204 274252
rect 333060 269068 333112 269074
rect 333060 269010 333112 269016
rect 332784 268456 332836 268462
rect 332784 268398 332836 268404
rect 332508 268388 332560 268394
rect 332508 268330 332560 268336
rect 332600 268388 332652 268394
rect 332600 268330 332652 268336
rect 332520 267782 332548 268330
rect 332508 267776 332560 267782
rect 332508 267718 332560 267724
rect 332612 264316 332640 268330
rect 332692 268252 332744 268258
rect 332692 268194 332744 268200
rect 332704 267918 332732 268194
rect 332796 268122 332824 268398
rect 332784 268116 332836 268122
rect 332784 268058 332836 268064
rect 332692 267912 332744 267918
rect 332692 267854 332744 267860
rect 333164 264330 333192 274246
rect 334176 273018 334204 277780
rect 334348 274236 334400 274242
rect 334348 274178 334400 274184
rect 334164 273012 334216 273018
rect 334164 272954 334216 272960
rect 333980 271040 334032 271046
rect 333980 270982 334032 270988
rect 333520 268456 333572 268462
rect 333520 268398 333572 268404
rect 333086 264302 333192 264330
rect 333532 264316 333560 268398
rect 333992 264316 334020 270982
rect 334360 264316 334388 274178
rect 335372 273086 335400 277780
rect 336096 274372 336148 274378
rect 336096 274314 336148 274320
rect 335360 273080 335412 273086
rect 335360 273022 335412 273028
rect 334808 271108 334860 271114
rect 334808 271050 334860 271056
rect 334820 264316 334848 271050
rect 335268 268524 335320 268530
rect 335268 268466 335320 268472
rect 335280 264316 335308 268466
rect 336108 264330 336136 274314
rect 336568 270434 336596 277780
rect 337108 274440 337160 274446
rect 337108 274382 337160 274388
rect 336740 271720 336792 271726
rect 336740 271662 336792 271668
rect 336648 271176 336700 271182
rect 336648 271118 336700 271124
rect 336556 270428 336608 270434
rect 336556 270370 336608 270376
rect 336188 268592 336240 268598
rect 336188 268534 336240 268540
rect 335754 264302 336136 264330
rect 336200 264316 336228 268534
rect 336660 264316 336688 271118
rect 336752 270366 336780 271662
rect 336740 270360 336792 270366
rect 336740 270302 336792 270308
rect 337120 264316 337148 274382
rect 337764 272338 337792 277780
rect 338960 272746 338988 277780
rect 339500 273216 339552 273222
rect 339500 273158 339552 273164
rect 338948 272740 339000 272746
rect 338948 272682 339000 272688
rect 337752 272332 337804 272338
rect 337752 272274 337804 272280
rect 339316 272332 339368 272338
rect 339316 272274 339368 272280
rect 337476 271312 337528 271318
rect 337476 271254 337528 271260
rect 337488 264316 337516 271254
rect 338856 268728 338908 268734
rect 338856 268670 338908 268676
rect 337936 268660 337988 268666
rect 337936 268602 337988 268608
rect 337948 264316 337976 268602
rect 338396 265872 338448 265878
rect 338396 265814 338448 265820
rect 338408 264316 338436 265814
rect 338868 264316 338896 268670
rect 339328 264316 339356 272274
rect 339512 270298 339540 273158
rect 340156 271250 340184 277780
rect 341064 274508 341116 274514
rect 341064 274450 341116 274456
rect 340236 271380 340288 271386
rect 340236 271322 340288 271328
rect 340144 271244 340196 271250
rect 340144 271186 340196 271192
rect 339500 270292 339552 270298
rect 339500 270234 339552 270240
rect 339776 265940 339828 265946
rect 339776 265882 339828 265888
rect 339788 264316 339816 265882
rect 340248 264330 340276 271322
rect 340788 270836 340840 270842
rect 340788 270778 340840 270784
rect 340800 270638 340828 270778
rect 340788 270632 340840 270638
rect 340788 270574 340840 270580
rect 340604 268796 340656 268802
rect 340604 268738 340656 268744
rect 340170 264302 340276 264330
rect 340616 264316 340644 268738
rect 341076 264316 341104 274450
rect 341352 272542 341380 277780
rect 341340 272536 341392 272542
rect 341340 272478 341392 272484
rect 342076 272536 342128 272542
rect 342076 272478 342128 272484
rect 341524 268864 341576 268870
rect 341524 268806 341576 268812
rect 341536 264316 341564 268806
rect 342088 264330 342116 272478
rect 342456 270230 342484 277780
rect 342536 274576 342588 274582
rect 342536 274518 342588 274524
rect 342444 270224 342496 270230
rect 342444 270166 342496 270172
rect 342548 264330 342576 274518
rect 343652 271726 343680 277780
rect 343732 275936 343784 275942
rect 343732 275878 343784 275884
rect 343640 271720 343692 271726
rect 343640 271662 343692 271668
rect 342812 271516 342864 271522
rect 342812 271458 342864 271464
rect 342010 264302 342116 264330
rect 342470 264302 342576 264330
rect 342824 264316 342852 271458
rect 343272 267912 343324 267918
rect 343272 267854 343324 267860
rect 343284 264316 343312 267854
rect 343744 264316 343772 275878
rect 344848 273222 344876 277780
rect 345112 276004 345164 276010
rect 345112 275946 345164 275952
rect 344836 273216 344888 273222
rect 344836 273158 344888 273164
rect 344008 273012 344060 273018
rect 344008 272954 344060 272960
rect 344020 270502 344048 272954
rect 344744 272740 344796 272746
rect 344744 272682 344796 272688
rect 344008 270496 344060 270502
rect 344008 270438 344060 270444
rect 344192 268932 344244 268938
rect 344192 268874 344244 268880
rect 344204 264316 344232 268874
rect 344756 264330 344784 272682
rect 344678 264302 344784 264330
rect 345124 264316 345152 275946
rect 346044 272950 346072 277780
rect 346032 272944 346084 272950
rect 346032 272886 346084 272892
rect 346860 270496 346912 270502
rect 346860 270438 346912 270444
rect 345480 270020 345532 270026
rect 345480 269962 345532 269968
rect 345492 264316 345520 269962
rect 345940 269000 345992 269006
rect 345940 268942 345992 268948
rect 345952 264316 345980 268942
rect 346400 266008 346452 266014
rect 346400 265950 346452 265956
rect 346412 264316 346440 265950
rect 346872 264316 346900 270438
rect 347240 270162 347268 277780
rect 348436 272882 348464 277780
rect 349068 275868 349120 275874
rect 349068 275810 349120 275816
rect 348424 272876 348476 272882
rect 348424 272818 348476 272824
rect 348240 271652 348292 271658
rect 348240 271594 348292 271600
rect 347596 271584 347648 271590
rect 347596 271526 347648 271532
rect 347228 270156 347280 270162
rect 347228 270098 347280 270104
rect 347608 264330 347636 271526
rect 347780 266076 347832 266082
rect 347780 266018 347832 266024
rect 347346 264302 347636 264330
rect 347792 264316 347820 266018
rect 348252 264316 348280 271594
rect 348608 270428 348660 270434
rect 348608 270370 348660 270376
rect 348620 264316 348648 270370
rect 349080 264316 349108 275810
rect 349528 270360 349580 270366
rect 349528 270302 349580 270308
rect 349540 264316 349568 270302
rect 349632 270094 349660 277780
rect 350172 275800 350224 275806
rect 350172 275742 350224 275748
rect 349988 271788 350040 271794
rect 349988 271730 350040 271736
rect 349620 270088 349672 270094
rect 349620 270030 349672 270036
rect 350000 264316 350028 271730
rect 350184 264330 350212 275742
rect 350736 267170 350764 277780
rect 351828 274100 351880 274106
rect 351828 274042 351880 274048
rect 351840 273562 351868 274042
rect 351828 273556 351880 273562
rect 351828 273498 351880 273504
rect 351932 272610 351960 277780
rect 353128 272814 353156 277780
rect 353116 272808 353168 272814
rect 353116 272750 353168 272756
rect 351920 272604 351972 272610
rect 351920 272546 351972 272552
rect 353116 272604 353168 272610
rect 353116 272546 353168 272552
rect 350908 271720 350960 271726
rect 350908 271662 350960 271668
rect 350724 267164 350776 267170
rect 350724 267106 350776 267112
rect 350184 264302 350474 264330
rect 350920 264316 350948 271662
rect 351736 270632 351788 270638
rect 351736 270574 351788 270580
rect 351276 270292 351328 270298
rect 351276 270234 351328 270240
rect 351288 264316 351316 270234
rect 351748 267986 351776 270574
rect 352196 270224 352248 270230
rect 352196 270166 352248 270172
rect 351920 269680 351972 269686
rect 351920 269622 351972 269628
rect 351828 269068 351880 269074
rect 351828 269010 351880 269016
rect 351840 268326 351868 269010
rect 351828 268320 351880 268326
rect 351828 268262 351880 268268
rect 351932 268190 351960 269622
rect 352012 269000 352064 269006
rect 352012 268942 352064 268948
rect 351920 268184 351972 268190
rect 351920 268126 351972 268132
rect 351736 267980 351788 267986
rect 351736 267922 351788 267928
rect 352024 267918 352052 268942
rect 352012 267912 352064 267918
rect 352012 267854 352064 267860
rect 351736 266144 351788 266150
rect 351736 266086 351788 266092
rect 351748 264316 351776 266086
rect 352208 264316 352236 270166
rect 353128 264974 353156 272546
rect 353576 270156 353628 270162
rect 353576 270098 353628 270104
rect 353208 266212 353260 266218
rect 353208 266154 353260 266160
rect 353036 264946 353156 264974
rect 353036 264330 353064 264946
rect 353220 264330 353248 266154
rect 352682 264302 353064 264330
rect 353142 264302 353248 264330
rect 353588 264316 353616 270098
rect 353942 268288 353998 268297
rect 353942 268223 353998 268232
rect 353956 264316 353984 268223
rect 354324 267102 354352 277780
rect 354404 275732 354456 275738
rect 354404 275674 354456 275680
rect 354312 267096 354364 267102
rect 354312 267038 354364 267044
rect 354416 264316 354444 275674
rect 354864 273216 354916 273222
rect 354864 273158 354916 273164
rect 354772 271448 354824 271454
rect 354772 271390 354824 271396
rect 354784 270026 354812 271390
rect 354772 270020 354824 270026
rect 354772 269962 354824 269968
rect 354876 264316 354904 273158
rect 355324 273148 355376 273154
rect 355324 273090 355376 273096
rect 355336 264316 355364 273090
rect 355520 272678 355548 277780
rect 355784 275664 355836 275670
rect 355784 275606 355836 275612
rect 355508 272672 355560 272678
rect 355508 272614 355560 272620
rect 355796 264316 355824 275606
rect 356716 272474 356744 277780
rect 356704 272468 356756 272474
rect 356704 272410 356756 272416
rect 357440 270564 357492 270570
rect 357440 270506 357492 270512
rect 356244 270088 356296 270094
rect 356244 270030 356296 270036
rect 356256 264316 356284 270030
rect 356610 268424 356666 268433
rect 356610 268359 356666 268368
rect 356624 264316 356652 268359
rect 357452 268054 357480 270506
rect 357440 268048 357492 268054
rect 357440 267990 357492 267996
rect 357532 268048 357584 268054
rect 357532 267990 357584 267996
rect 357072 266280 357124 266286
rect 357072 266222 357124 266228
rect 357084 264316 357112 266222
rect 357544 264316 357572 267990
rect 357912 267034 357940 277780
rect 358452 275596 358504 275602
rect 358452 275538 358504 275544
rect 357992 272944 358044 272950
rect 357992 272886 358044 272892
rect 357900 267028 357952 267034
rect 357900 266970 357952 266976
rect 358004 264316 358032 272886
rect 358464 264316 358492 275538
rect 358820 273080 358872 273086
rect 358820 273022 358872 273028
rect 358728 268048 358780 268054
rect 358832 268036 358860 273022
rect 359016 272270 359044 277780
rect 360212 272406 360240 277780
rect 361120 275528 361172 275534
rect 361120 275470 361172 275476
rect 360660 272876 360712 272882
rect 360660 272818 360712 272824
rect 360568 272808 360620 272814
rect 360568 272750 360620 272756
rect 360200 272400 360252 272406
rect 360200 272342 360252 272348
rect 359004 272264 359056 272270
rect 359004 272206 359056 272212
rect 358910 268696 358966 268705
rect 358910 268631 358966 268640
rect 358780 268008 358860 268036
rect 358728 267990 358780 267996
rect 358924 264316 358952 268631
rect 359370 268560 359426 268569
rect 359370 268495 359426 268504
rect 359384 264316 359412 268495
rect 359740 267708 359792 267714
rect 359740 267650 359792 267656
rect 359752 264316 359780 267650
rect 360580 264330 360608 272750
rect 360226 264302 360608 264330
rect 360672 264316 360700 272818
rect 361132 264316 361160 275470
rect 361408 266966 361436 277780
rect 362604 273018 362632 277780
rect 362960 273216 363012 273222
rect 362960 273158 363012 273164
rect 362592 273012 362644 273018
rect 362592 272954 362644 272960
rect 362972 272610 363000 273158
rect 363144 272672 363196 272678
rect 363144 272614 363196 272620
rect 362960 272604 363012 272610
rect 362960 272546 363012 272552
rect 361580 269680 361632 269686
rect 361580 269622 361632 269628
rect 361396 266960 361448 266966
rect 361396 266902 361448 266908
rect 361592 264316 361620 269622
rect 362038 268832 362094 268841
rect 362038 268767 362094 268776
rect 362052 264316 362080 268767
rect 362408 267640 362460 267646
rect 362408 267582 362460 267588
rect 362420 264316 362448 267582
rect 363156 264330 363184 272614
rect 363326 271416 363382 271425
rect 363326 271351 363382 271360
rect 362894 264302 363184 264330
rect 363340 264316 363368 271351
rect 363800 267850 363828 277780
rect 364064 275460 364116 275466
rect 364064 275402 364116 275408
rect 363788 267844 363840 267850
rect 363788 267786 363840 267792
rect 364076 264330 364104 275402
rect 364708 270020 364760 270026
rect 364708 269962 364760 269968
rect 364246 268968 364302 268977
rect 364246 268903 364302 268912
rect 363814 264302 364104 264330
rect 364260 264316 364288 268903
rect 364720 264316 364748 269962
rect 364996 266898 365024 277780
rect 365534 271688 365590 271697
rect 365534 271623 365590 271632
rect 365076 267572 365128 267578
rect 365076 267514 365128 267520
rect 364984 266892 365036 266898
rect 364984 266834 365036 266840
rect 365088 264316 365116 267514
rect 365548 264316 365576 271623
rect 365994 271552 366050 271561
rect 365994 271487 366050 271496
rect 366008 264316 366036 271487
rect 366100 269958 366128 277780
rect 366456 275392 366508 275398
rect 366456 275334 366508 275340
rect 366088 269952 366140 269958
rect 366088 269894 366140 269900
rect 366468 264316 366496 275334
rect 367296 272202 367324 277780
rect 368204 272604 368256 272610
rect 368204 272546 368256 272552
rect 367284 272196 367336 272202
rect 367284 272138 367336 272144
rect 366914 270464 366970 270473
rect 366914 270399 366970 270408
rect 366928 264316 366956 270399
rect 367376 269952 367428 269958
rect 367376 269894 367428 269900
rect 367388 264316 367416 269894
rect 367744 267504 367796 267510
rect 367744 267446 367796 267452
rect 367756 264316 367784 267446
rect 368216 264316 368244 272546
rect 368492 266830 368520 277780
rect 369124 275324 369176 275330
rect 369124 275266 369176 275272
rect 368662 273184 368718 273193
rect 368662 273119 368718 273128
rect 368480 266824 368532 266830
rect 368480 266766 368532 266772
rect 368676 264316 368704 273119
rect 369136 264316 369164 275266
rect 369582 270328 369638 270337
rect 369582 270263 369638 270272
rect 369596 264316 369624 270263
rect 369688 269890 369716 277780
rect 369676 269884 369728 269890
rect 369676 269826 369728 269832
rect 370044 269884 370096 269890
rect 370044 269826 370096 269832
rect 370056 264316 370084 269826
rect 370884 269822 370912 277780
rect 371792 275256 371844 275262
rect 371792 275198 371844 275204
rect 371238 273048 371294 273057
rect 371238 272983 371294 272992
rect 370872 269816 370924 269822
rect 370872 269758 370924 269764
rect 370504 267436 370556 267442
rect 370504 267378 370556 267384
rect 370516 264316 370544 267378
rect 371252 264330 371280 272983
rect 371330 272912 371386 272921
rect 371330 272847 371386 272856
rect 370898 264302 371280 264330
rect 371344 264316 371372 272847
rect 371804 264316 371832 275198
rect 372080 266762 372108 277780
rect 373172 272468 373224 272474
rect 373172 272410 373224 272416
rect 372250 270192 372306 270201
rect 372250 270127 372306 270136
rect 372068 266756 372120 266762
rect 372068 266698 372120 266704
rect 372264 264316 372292 270127
rect 372712 268048 372764 268054
rect 372712 267990 372764 267996
rect 372724 264316 372752 267990
rect 373184 264316 373212 272410
rect 373276 269822 373304 277780
rect 373998 272776 374054 272785
rect 373998 272711 374054 272720
rect 373264 269816 373316 269822
rect 373264 269758 373316 269764
rect 373540 267368 373592 267374
rect 373540 267310 373592 267316
rect 373552 264316 373580 267310
rect 374012 264316 374040 272711
rect 374380 272134 374408 277780
rect 374920 275188 374972 275194
rect 374920 275130 374972 275136
rect 374368 272128 374420 272134
rect 374368 272070 374420 272076
rect 374460 267300 374512 267306
rect 374460 267242 374512 267248
rect 374472 264316 374500 267242
rect 374932 264316 374960 275130
rect 375380 269748 375432 269754
rect 375380 269690 375432 269696
rect 375392 264316 375420 269690
rect 375576 266694 375604 277780
rect 376668 272400 376720 272406
rect 376668 272342 376720 272348
rect 376208 267232 376260 267238
rect 376208 267174 376260 267180
rect 375840 267164 375892 267170
rect 375840 267106 375892 267112
rect 375564 266688 375616 266694
rect 375564 266630 375616 266636
rect 375852 264316 375880 267106
rect 376220 264316 376248 267174
rect 376680 264316 376708 272342
rect 376772 267782 376800 277780
rect 377588 275120 377640 275126
rect 377588 275062 377640 275068
rect 376760 267776 376812 267782
rect 376760 267718 376812 267724
rect 377128 267096 377180 267102
rect 377128 267038 377180 267044
rect 377140 264316 377168 267038
rect 377600 264316 377628 275062
rect 377968 270706 377996 277780
rect 377956 270700 378008 270706
rect 377956 270642 378008 270648
rect 378046 270056 378102 270065
rect 378046 269991 378102 270000
rect 378060 264316 378088 269991
rect 378508 267028 378560 267034
rect 378508 266970 378560 266976
rect 378520 264316 378548 266970
rect 378876 266960 378928 266966
rect 378876 266902 378928 266908
rect 378888 264316 378916 266902
rect 379164 266626 379192 277780
rect 380256 275052 380308 275058
rect 380256 274994 380308 275000
rect 379334 272640 379390 272649
rect 379334 272575 379390 272584
rect 379152 266620 379204 266626
rect 379152 266562 379204 266568
rect 379348 264316 379376 272575
rect 379796 266892 379848 266898
rect 379796 266834 379848 266840
rect 379808 264316 379836 266834
rect 380268 264316 380296 274994
rect 380360 269618 380388 277780
rect 381556 272066 381584 277780
rect 382004 272264 382056 272270
rect 382004 272206 382056 272212
rect 381544 272060 381596 272066
rect 381544 272002 381596 272008
rect 380348 269612 380400 269618
rect 380348 269554 380400 269560
rect 380716 269612 380768 269618
rect 380716 269554 380768 269560
rect 380728 264316 380756 269554
rect 381636 266824 381688 266830
rect 381636 266766 381688 266772
rect 381176 266756 381228 266762
rect 381176 266698 381228 266704
rect 381188 264316 381216 266698
rect 381648 264316 381676 266766
rect 382016 264316 382044 272206
rect 382464 270020 382516 270026
rect 382464 269962 382516 269968
rect 382476 269906 382504 269962
rect 382292 269878 382504 269906
rect 382292 269686 382320 269878
rect 382464 269748 382516 269754
rect 382464 269690 382516 269696
rect 382280 269680 382332 269686
rect 382280 269622 382332 269628
rect 382476 268054 382504 269690
rect 382464 268048 382516 268054
rect 382464 267990 382516 267996
rect 382464 266688 382516 266694
rect 382464 266630 382516 266636
rect 382188 266348 382240 266354
rect 382188 266290 382240 266296
rect 382200 265810 382228 266290
rect 382096 265804 382148 265810
rect 382096 265746 382148 265752
rect 382188 265804 382240 265810
rect 382188 265746 382240 265752
rect 382108 265690 382136 265746
rect 382108 265674 382320 265690
rect 382108 265668 382332 265674
rect 382108 265662 382280 265668
rect 382280 265610 382332 265616
rect 382476 264316 382504 266630
rect 382660 266558 382688 277780
rect 382924 274984 382976 274990
rect 382924 274926 382976 274932
rect 382648 266552 382700 266558
rect 382648 266494 382700 266500
rect 382936 264316 382964 274926
rect 383382 269920 383438 269929
rect 383382 269855 383438 269864
rect 383396 264316 383424 269855
rect 383856 269550 383884 277780
rect 384672 272196 384724 272202
rect 384672 272138 384724 272144
rect 383844 269544 383896 269550
rect 383844 269486 383896 269492
rect 384304 266620 384356 266626
rect 384304 266562 384356 266568
rect 383844 266552 383896 266558
rect 383844 266494 383896 266500
rect 383856 264316 383884 266494
rect 384316 264316 384344 266562
rect 384684 264316 384712 272138
rect 385052 270570 385080 277780
rect 385592 274916 385644 274922
rect 385592 274858 385644 274864
rect 385040 270564 385092 270570
rect 385040 270506 385092 270512
rect 385130 266112 385186 266121
rect 385130 266047 385186 266056
rect 385144 264316 385172 266047
rect 385604 264316 385632 274858
rect 386052 269544 386104 269550
rect 386052 269486 386104 269492
rect 386064 264316 386092 269486
rect 386248 266490 386276 277780
rect 387340 272128 387392 272134
rect 387340 272070 387392 272076
rect 386970 267608 387026 267617
rect 386970 267543 387026 267552
rect 386236 266484 386288 266490
rect 386236 266426 386288 266432
rect 386510 266248 386566 266257
rect 386510 266183 386566 266192
rect 386524 264316 386552 266183
rect 386984 264316 387012 267543
rect 387352 264316 387380 272070
rect 387444 269482 387472 277780
rect 388258 275904 388314 275913
rect 388258 275839 388314 275848
rect 387432 269476 387484 269482
rect 387432 269418 387484 269424
rect 387798 267744 387854 267753
rect 387798 267679 387854 267688
rect 387812 264316 387840 267679
rect 388272 264316 388300 275839
rect 388640 271998 388668 277780
rect 388628 271992 388680 271998
rect 388628 271934 388680 271940
rect 388720 269476 388772 269482
rect 388720 269418 388772 269424
rect 388732 264316 388760 269418
rect 389638 267472 389694 267481
rect 389638 267407 389694 267416
rect 389180 266484 389232 266490
rect 389180 266426 389232 266432
rect 389192 264316 389220 266426
rect 389652 264316 389680 267407
rect 389744 265266 389772 277780
rect 390940 269414 390968 277780
rect 391294 275768 391350 275777
rect 391294 275703 391350 275712
rect 390928 269408 390980 269414
rect 390928 269350 390980 269356
rect 390008 268048 390060 268054
rect 390008 267990 390060 267996
rect 389732 265260 389784 265266
rect 389732 265202 389784 265208
rect 390020 264316 390048 267990
rect 390466 267336 390522 267345
rect 390466 267271 390522 267280
rect 390480 264316 390508 267271
rect 391308 264330 391336 275703
rect 391386 269784 391442 269793
rect 391386 269719 391442 269728
rect 390954 264302 391336 264330
rect 391400 264316 391428 269719
rect 392136 269346 392164 277780
rect 392766 272504 392822 272513
rect 392766 272439 392822 272448
rect 392124 269340 392176 269346
rect 392124 269282 392176 269288
rect 391846 267200 391902 267209
rect 391846 267135 391902 267144
rect 391860 264316 391888 267135
rect 392308 266416 392360 266422
rect 392308 266358 392360 266364
rect 392320 264316 392348 266358
rect 392780 264316 392808 272439
rect 393134 267064 393190 267073
rect 393134 266999 393190 267008
rect 393148 264316 393176 266999
rect 393332 266354 393360 277780
rect 393594 275632 393650 275641
rect 393594 275567 393650 275576
rect 393320 266348 393372 266354
rect 393320 266290 393372 266296
rect 393608 264316 393636 275567
rect 394528 270638 394556 277780
rect 394608 272060 394660 272066
rect 394608 272002 394660 272008
rect 394516 270632 394568 270638
rect 394516 270574 394568 270580
rect 394056 269408 394108 269414
rect 394056 269350 394108 269356
rect 394068 264316 394096 269350
rect 394620 268054 394648 272002
rect 395436 271992 395488 271998
rect 395436 271934 395488 271940
rect 394608 268048 394660 268054
rect 394608 267990 394660 267996
rect 394514 266928 394570 266937
rect 394514 266863 394570 266872
rect 394528 264316 394556 266863
rect 394976 266348 395028 266354
rect 394976 266290 395028 266296
rect 394988 264316 395016 266290
rect 395448 264316 395476 271934
rect 395724 270774 395752 277780
rect 396262 275496 396318 275505
rect 396262 275431 396318 275440
rect 395712 270768 395764 270774
rect 395712 270710 395764 270716
rect 395802 266792 395858 266801
rect 395802 266727 395858 266736
rect 395816 264316 395844 266727
rect 396276 264316 396304 275431
rect 396724 269340 396776 269346
rect 396724 269282 396776 269288
rect 396736 264316 396764 269282
rect 396920 265810 396948 277780
rect 397182 266656 397238 266665
rect 397182 266591 397238 266600
rect 396908 265804 396960 265810
rect 396908 265746 396960 265752
rect 397196 264316 397224 266591
rect 397644 265804 397696 265810
rect 397644 265746 397696 265752
rect 397656 264316 397684 265746
rect 398024 265674 398052 277780
rect 398930 275360 398986 275369
rect 398930 275295 398986 275304
rect 398102 272368 398158 272377
rect 398102 272303 398158 272312
rect 398012 265668 398064 265674
rect 398012 265610 398064 265616
rect 398116 264316 398144 272303
rect 398470 266520 398526 266529
rect 398470 266455 398526 266464
rect 398484 264316 398512 266455
rect 398944 264316 398972 275295
rect 399220 269278 399248 277780
rect 399208 269272 399260 269278
rect 399208 269214 399260 269220
rect 399392 269272 399444 269278
rect 399392 269214 399444 269220
rect 399404 264316 399432 269214
rect 399850 266384 399906 266393
rect 399850 266319 399906 266328
rect 399864 264316 399892 266319
rect 400312 265668 400364 265674
rect 400312 265610 400364 265616
rect 400324 264316 400352 265610
rect 400416 265334 400444 277780
rect 401612 274854 401640 277780
rect 401690 275224 401746 275233
rect 401690 275159 401746 275168
rect 401600 274848 401652 274854
rect 401600 274790 401652 274796
rect 401140 273488 401192 273494
rect 401140 273430 401192 273436
rect 400772 268048 400824 268054
rect 400772 267990 400824 267996
rect 400404 265328 400456 265334
rect 400404 265270 400456 265276
rect 400784 264316 400812 267990
rect 401152 264316 401180 273430
rect 401704 264330 401732 275159
rect 402702 274952 402758 274961
rect 402702 274887 402758 274896
rect 402058 269648 402114 269657
rect 402058 269583 402114 269592
rect 401626 264302 401732 264330
rect 402072 264316 402100 269583
rect 402716 264330 402744 274887
rect 402808 271930 402836 277780
rect 403900 274848 403952 274854
rect 403900 274790 403952 274796
rect 403438 272232 403494 272241
rect 403438 272167 403494 272176
rect 402796 271924 402848 271930
rect 402796 271866 402848 271872
rect 402888 271924 402940 271930
rect 402888 271866 402940 271872
rect 402900 268054 402928 271866
rect 402888 268048 402940 268054
rect 402888 267990 402940 267996
rect 402980 265328 403032 265334
rect 402980 265270 403032 265276
rect 402546 264302 402744 264330
rect 402992 264316 403020 265270
rect 403452 264316 403480 272167
rect 403912 264316 403940 274790
rect 404004 265198 404032 277780
rect 404266 275088 404322 275097
rect 404266 275023 404322 275032
rect 403992 265192 404044 265198
rect 403992 265134 404044 265140
rect 404280 264316 404308 275023
rect 405200 274786 405228 277780
rect 405370 274816 405426 274825
rect 405188 274780 405240 274786
rect 405370 274751 405426 274760
rect 405188 274722 405240 274728
rect 404726 269512 404782 269521
rect 404726 269447 404782 269456
rect 404740 264316 404768 269447
rect 405384 264330 405412 274751
rect 406304 269210 406332 277780
rect 406568 274780 406620 274786
rect 406568 274722 406620 274728
rect 406292 269204 406344 269210
rect 406292 269146 406344 269152
rect 406108 268048 406160 268054
rect 406108 267990 406160 267996
rect 405462 265976 405518 265985
rect 405462 265911 405518 265920
rect 405214 264302 405412 264330
rect 405476 264330 405504 265911
rect 405476 264302 405674 264330
rect 406120 264316 406148 267990
rect 406580 264316 406608 274722
rect 407500 274718 407528 277780
rect 407488 274712 407540 274718
rect 406934 274680 406990 274689
rect 407488 274654 407540 274660
rect 406934 274615 406990 274624
rect 406948 264316 406976 274615
rect 408222 274544 408278 274553
rect 408222 274479 408278 274488
rect 407394 269376 407450 269385
rect 407394 269311 407450 269320
rect 407408 264316 407436 269311
rect 408236 264330 408264 274479
rect 408314 265840 408370 265849
rect 408314 265775 408370 265784
rect 407882 264302 408264 264330
rect 408328 264316 408356 265775
rect 408696 265402 408724 277780
rect 409236 274712 409288 274718
rect 409236 274654 409288 274660
rect 408774 272096 408830 272105
rect 408774 272031 408830 272040
rect 408684 265396 408736 265402
rect 408684 265338 408736 265344
rect 408788 264316 408816 272031
rect 409248 264316 409276 274654
rect 409892 271862 409920 277780
rect 411088 274650 411116 277780
rect 411076 274644 411128 274650
rect 411076 274586 411128 274592
rect 410890 271960 410946 271969
rect 410890 271895 410946 271904
rect 409880 271856 409932 271862
rect 409880 271798 409932 271804
rect 409602 269240 409658 269249
rect 409602 269175 409658 269184
rect 409616 264316 409644 269175
rect 410062 269104 410118 269113
rect 410062 269039 410118 269048
rect 410076 264316 410104 269039
rect 410904 264330 410932 271895
rect 411996 271856 412048 271862
rect 411074 271824 411130 271833
rect 411996 271798 412048 271804
rect 411074 271759 411130 271768
rect 411088 264330 411116 271759
rect 411812 270564 411864 270570
rect 411812 270506 411864 270512
rect 411444 269204 411496 269210
rect 411444 269146 411496 269152
rect 410550 264302 410932 264330
rect 411010 264302 411116 264330
rect 411456 264316 411484 269146
rect 411824 269142 411852 270506
rect 411812 269136 411864 269142
rect 411812 269078 411864 269084
rect 411904 269136 411956 269142
rect 411904 269078 411956 269084
rect 411916 264316 411944 269078
rect 412008 268054 412036 271798
rect 411996 268048 412048 268054
rect 411996 267990 412048 267996
rect 412284 265470 412312 277780
rect 413112 277766 413402 277794
rect 413112 270570 413140 277766
rect 414584 273562 414612 277780
rect 414572 273556 414624 273562
rect 414572 273498 414624 273504
rect 415308 271176 415360 271182
rect 415308 271118 415360 271124
rect 415320 271046 415348 271118
rect 415308 271040 415360 271046
rect 415308 270982 415360 270988
rect 413100 270564 413152 270570
rect 413100 270506 413152 270512
rect 415780 265538 415808 277780
rect 416976 270638 417004 277780
rect 418172 273766 418200 277780
rect 418160 273760 418212 273766
rect 418160 273702 418212 273708
rect 416964 270632 417016 270638
rect 416964 270574 417016 270580
rect 419368 265606 419396 277780
rect 420564 268122 420592 277780
rect 420920 274848 420972 274854
rect 420920 274790 420972 274796
rect 420932 273494 420960 274790
rect 421668 273630 421696 277780
rect 422864 273834 422892 277780
rect 422852 273828 422904 273834
rect 422852 273770 422904 273776
rect 421656 273624 421708 273630
rect 421656 273566 421708 273572
rect 420920 273488 420972 273494
rect 420920 273430 420972 273436
rect 420920 271176 420972 271182
rect 420748 271124 420920 271130
rect 420748 271118 420972 271124
rect 420748 271114 420960 271118
rect 420736 271108 420960 271114
rect 420788 271102 420960 271108
rect 420736 271050 420788 271056
rect 424060 270706 424088 277780
rect 425256 273970 425284 277780
rect 425244 273964 425296 273970
rect 425244 273906 425296 273912
rect 424048 270700 424100 270706
rect 424048 270642 424100 270648
rect 426452 268258 426480 277780
rect 426440 268252 426492 268258
rect 426440 268194 426492 268200
rect 427648 268190 427676 277780
rect 428844 273902 428872 277780
rect 428832 273896 428884 273902
rect 428832 273838 428884 273844
rect 427636 268184 427688 268190
rect 427636 268126 427688 268132
rect 420552 268116 420604 268122
rect 420552 268058 420604 268064
rect 429948 265742 429976 277780
rect 431144 270842 431172 277780
rect 432340 274106 432368 277780
rect 432328 274100 432380 274106
rect 432328 274042 432380 274048
rect 431132 270836 431184 270842
rect 431132 270778 431184 270784
rect 433536 268326 433564 277780
rect 434732 270910 434760 277780
rect 435928 274038 435956 277780
rect 437032 274174 437060 277780
rect 437020 274168 437072 274174
rect 437020 274110 437072 274116
rect 435916 274032 435968 274038
rect 435916 273974 435968 273980
rect 434720 270904 434772 270910
rect 434720 270846 434772 270852
rect 438228 268394 438256 277780
rect 439424 274310 439452 277780
rect 439412 274304 439464 274310
rect 439412 274246 439464 274252
rect 440620 268462 440648 277780
rect 441816 271182 441844 277780
rect 443012 274242 443040 277780
rect 443000 274236 443052 274242
rect 443000 274178 443052 274184
rect 441804 271176 441856 271182
rect 441804 271118 441856 271124
rect 444208 271114 444236 277780
rect 444196 271108 444248 271114
rect 444196 271050 444248 271056
rect 445312 268530 445340 277780
rect 446508 274378 446536 277780
rect 446496 274372 446548 274378
rect 446496 274314 446548 274320
rect 447704 268598 447732 277780
rect 448900 271250 448928 277780
rect 450096 274446 450124 277780
rect 450084 274440 450136 274446
rect 450084 274382 450136 274388
rect 451292 271318 451320 277780
rect 451280 271312 451332 271318
rect 451280 271254 451332 271260
rect 448888 271244 448940 271250
rect 448888 271186 448940 271192
rect 452488 268666 452516 277780
rect 452476 268660 452528 268666
rect 452476 268602 452528 268608
rect 447692 268592 447744 268598
rect 447692 268534 447744 268540
rect 445300 268524 445352 268530
rect 445300 268466 445352 268472
rect 440608 268456 440660 268462
rect 440608 268398 440660 268404
rect 438216 268388 438268 268394
rect 438216 268330 438268 268336
rect 433524 268320 433576 268326
rect 433524 268262 433576 268268
rect 453592 265878 453620 277780
rect 454788 268734 454816 277780
rect 455984 272338 456012 277780
rect 455972 272332 456024 272338
rect 455972 272274 456024 272280
rect 454776 268728 454828 268734
rect 454776 268670 454828 268676
rect 457180 265946 457208 277780
rect 458376 271386 458404 277780
rect 459468 272332 459520 272338
rect 459468 272274 459520 272280
rect 458364 271380 458416 271386
rect 458364 271322 458416 271328
rect 457168 265940 457220 265946
rect 457168 265882 457220 265888
rect 453580 265872 453632 265878
rect 459480 265849 459508 272274
rect 459572 268802 459600 277780
rect 460676 274514 460704 277780
rect 460664 274508 460716 274514
rect 460664 274450 460716 274456
rect 461872 268870 461900 277780
rect 463068 272542 463096 277780
rect 464264 274582 464292 277780
rect 464252 274576 464304 274582
rect 464252 274518 464304 274524
rect 463056 272536 463108 272542
rect 463056 272478 463108 272484
rect 465460 271522 465488 277780
rect 465908 272536 465960 272542
rect 465908 272478 465960 272484
rect 465448 271516 465500 271522
rect 465448 271458 465500 271464
rect 461860 268864 461912 268870
rect 461860 268806 461912 268812
rect 459560 268796 459612 268802
rect 459560 268738 459612 268744
rect 465920 265985 465948 272478
rect 466656 269006 466684 277780
rect 467852 275942 467880 277780
rect 467840 275936 467892 275942
rect 467840 275878 467892 275884
rect 466644 269000 466696 269006
rect 466644 268942 466696 268948
rect 468956 268938 468984 277780
rect 470152 272746 470180 277780
rect 471348 276010 471376 277780
rect 471336 276004 471388 276010
rect 471336 275946 471388 275952
rect 470140 272740 470192 272746
rect 470140 272682 470192 272688
rect 471980 272740 472032 272746
rect 471980 272682 472032 272688
rect 468944 268932 468996 268938
rect 468944 268874 468996 268880
rect 465906 265976 465962 265985
rect 465906 265911 465962 265920
rect 453580 265814 453632 265820
rect 459466 265840 459522 265849
rect 459466 265775 459522 265784
rect 429936 265736 429988 265742
rect 429936 265678 429988 265684
rect 419356 265600 419408 265606
rect 419356 265542 419408 265548
rect 415768 265532 415820 265538
rect 415768 265474 415820 265480
rect 412272 265464 412324 265470
rect 412272 265406 412324 265412
rect 471992 265334 472020 272682
rect 472544 271454 472572 277780
rect 472532 271448 472584 271454
rect 472532 271390 472584 271396
rect 473740 269074 473768 277780
rect 473728 269068 473780 269074
rect 473728 269010 473780 269016
rect 474936 266014 474964 277780
rect 476132 270502 476160 277780
rect 477236 271590 477264 277780
rect 477224 271584 477276 271590
rect 477224 271526 477276 271532
rect 476120 270496 476172 270502
rect 476120 270438 476172 270444
rect 478432 266082 478460 277780
rect 479628 271658 479656 277780
rect 479616 271652 479668 271658
rect 479616 271594 479668 271600
rect 480824 270434 480852 277780
rect 482020 275874 482048 277780
rect 482008 275868 482060 275874
rect 482008 275810 482060 275816
rect 480812 270428 480864 270434
rect 480812 270370 480864 270376
rect 483216 270366 483244 277780
rect 484320 271794 484348 277780
rect 485516 275806 485544 277780
rect 485504 275800 485556 275806
rect 485504 275742 485556 275748
rect 484308 271788 484360 271794
rect 484308 271730 484360 271736
rect 486712 271726 486740 277780
rect 486700 271720 486752 271726
rect 486700 271662 486752 271668
rect 483204 270360 483256 270366
rect 483204 270302 483256 270308
rect 487908 270298 487936 277780
rect 487896 270292 487948 270298
rect 487896 270234 487948 270240
rect 489104 266150 489132 277780
rect 490300 270230 490328 277780
rect 491496 273222 491524 277780
rect 491484 273216 491536 273222
rect 491484 273158 491536 273164
rect 490288 270224 490340 270230
rect 490288 270166 490340 270172
rect 492600 266218 492628 277780
rect 493796 270162 493824 277780
rect 493784 270156 493836 270162
rect 493784 270098 493836 270104
rect 494992 268297 495020 277780
rect 496188 275738 496216 277780
rect 496176 275732 496228 275738
rect 496176 275674 496228 275680
rect 497384 273154 497412 277780
rect 497372 273148 497424 273154
rect 497372 273090 497424 273096
rect 498580 273086 498608 277780
rect 499776 275670 499804 277780
rect 499764 275664 499816 275670
rect 499764 275606 499816 275612
rect 498568 273080 498620 273086
rect 498568 273022 498620 273028
rect 498844 273080 498896 273086
rect 498844 273022 498896 273028
rect 494978 268288 495034 268297
rect 494978 268223 495034 268232
rect 492588 266212 492640 266218
rect 492588 266154 492640 266160
rect 489092 266144 489144 266150
rect 489092 266086 489144 266092
rect 478420 266076 478472 266082
rect 478420 266018 478472 266024
rect 474924 266008 474976 266014
rect 474924 265950 474976 265956
rect 498856 265674 498884 273022
rect 500880 270094 500908 277780
rect 500868 270088 500920 270094
rect 500868 270030 500920 270036
rect 502076 268433 502104 277780
rect 502062 268424 502118 268433
rect 502062 268359 502118 268368
rect 503272 266286 503300 277780
rect 504468 273018 504496 277780
rect 504456 273012 504508 273018
rect 504456 272954 504508 272960
rect 505664 272950 505692 277780
rect 506860 275602 506888 277780
rect 506848 275596 506900 275602
rect 506848 275538 506900 275544
rect 505652 272944 505704 272950
rect 505652 272886 505704 272892
rect 507964 268705 507992 277780
rect 507950 268696 508006 268705
rect 507950 268631 508006 268640
rect 509160 268569 509188 277780
rect 509146 268560 509202 268569
rect 509146 268495 509202 268504
rect 510356 267714 510384 277780
rect 511552 272814 511580 277780
rect 512748 272882 512776 277780
rect 513944 275534 513972 277780
rect 513932 275528 513984 275534
rect 513932 275470 513984 275476
rect 512736 272876 512788 272882
rect 512736 272818 512788 272824
rect 511540 272808 511592 272814
rect 511540 272750 511592 272756
rect 511632 272808 511684 272814
rect 511632 272750 511684 272756
rect 510344 267708 510396 267714
rect 510344 267650 510396 267656
rect 503260 266280 503312 266286
rect 503260 266222 503312 266228
rect 511644 265810 511672 272750
rect 515140 270026 515168 277780
rect 515128 270020 515180 270026
rect 515128 269962 515180 269968
rect 516244 268841 516272 277780
rect 516230 268832 516286 268841
rect 516230 268767 516286 268776
rect 517440 267646 517468 277780
rect 518636 272678 518664 277780
rect 518624 272672 518676 272678
rect 518624 272614 518676 272620
rect 519832 271425 519860 277780
rect 521028 275466 521056 277780
rect 521016 275460 521068 275466
rect 521016 275402 521068 275408
rect 519818 271416 519874 271425
rect 519818 271351 519874 271360
rect 522224 268977 522252 277780
rect 523420 269958 523448 277780
rect 523408 269952 523460 269958
rect 523408 269894 523460 269900
rect 522210 268968 522266 268977
rect 522210 268903 522266 268912
rect 517428 267640 517480 267646
rect 517428 267582 517480 267588
rect 524524 267578 524552 277780
rect 525720 271697 525748 277780
rect 525706 271688 525762 271697
rect 525706 271623 525762 271632
rect 526916 271561 526944 277780
rect 528112 275398 528140 277780
rect 528100 275392 528152 275398
rect 528100 275334 528152 275340
rect 526902 271552 526958 271561
rect 526902 271487 526958 271496
rect 529308 270473 529336 277780
rect 529294 270464 529350 270473
rect 529294 270399 529350 270408
rect 530504 269890 530532 277780
rect 530492 269884 530544 269890
rect 530492 269826 530544 269832
rect 524512 267572 524564 267578
rect 524512 267514 524564 267520
rect 531608 267510 531636 277780
rect 532804 272610 532832 277780
rect 534000 273193 534028 277780
rect 535196 275330 535224 277780
rect 535184 275324 535236 275330
rect 535184 275266 535236 275272
rect 533986 273184 534042 273193
rect 533986 273119 534042 273128
rect 532792 272604 532844 272610
rect 532792 272546 532844 272552
rect 536392 270337 536420 277780
rect 536378 270328 536434 270337
rect 536378 270263 536434 270272
rect 537588 269822 537616 277780
rect 537576 269816 537628 269822
rect 537576 269758 537628 269764
rect 531596 267504 531648 267510
rect 531596 267446 531648 267452
rect 538784 267442 538812 277780
rect 539888 273057 539916 277780
rect 539874 273048 539930 273057
rect 539874 272983 539930 272992
rect 541084 272921 541112 277780
rect 542280 275262 542308 277780
rect 542268 275256 542320 275262
rect 542268 275198 542320 275204
rect 541070 272912 541126 272921
rect 541070 272847 541126 272856
rect 543476 270201 543504 277780
rect 543462 270192 543518 270201
rect 543462 270127 543518 270136
rect 544672 269754 544700 277780
rect 545868 272474 545896 277780
rect 545856 272468 545908 272474
rect 545856 272410 545908 272416
rect 544660 269748 544712 269754
rect 544660 269690 544712 269696
rect 538772 267436 538824 267442
rect 538772 267378 538824 267384
rect 547064 267374 547092 277780
rect 548168 272785 548196 277780
rect 548154 272776 548210 272785
rect 548154 272711 548210 272720
rect 547052 267368 547104 267374
rect 547052 267310 547104 267316
rect 549364 267306 549392 277780
rect 550560 275194 550588 277780
rect 550548 275188 550600 275194
rect 550548 275130 550600 275136
rect 551756 269686 551784 277780
rect 551744 269680 551796 269686
rect 551744 269622 551796 269628
rect 549352 267300 549404 267306
rect 549352 267242 549404 267248
rect 552952 267170 552980 277780
rect 554148 267238 554176 277780
rect 555252 272406 555280 277780
rect 555240 272400 555292 272406
rect 555240 272342 555292 272348
rect 554136 267232 554188 267238
rect 554136 267174 554188 267180
rect 552940 267164 552992 267170
rect 552940 267106 552992 267112
rect 556448 267102 556476 277780
rect 557644 275126 557672 277780
rect 557632 275120 557684 275126
rect 557632 275062 557684 275068
rect 558840 270065 558868 277780
rect 558826 270056 558882 270065
rect 558826 269991 558882 270000
rect 556436 267096 556488 267102
rect 556436 267038 556488 267044
rect 560036 267034 560064 277780
rect 560024 267028 560076 267034
rect 560024 266970 560076 266976
rect 561232 266966 561260 277780
rect 562428 272649 562456 277780
rect 562414 272640 562470 272649
rect 562414 272575 562470 272584
rect 561220 266960 561272 266966
rect 561220 266902 561272 266908
rect 563532 266898 563560 277780
rect 564728 275058 564756 277780
rect 564716 275052 564768 275058
rect 564716 274994 564768 275000
rect 565924 269618 565952 277780
rect 565912 269612 565964 269618
rect 565912 269554 565964 269560
rect 563520 266892 563572 266898
rect 563520 266834 563572 266840
rect 567120 266762 567148 277780
rect 568316 266830 568344 277780
rect 569512 272270 569540 277780
rect 569500 272264 569552 272270
rect 569500 272206 569552 272212
rect 568304 266824 568356 266830
rect 568304 266766 568356 266772
rect 567108 266756 567160 266762
rect 567108 266698 567160 266704
rect 570708 266694 570736 277780
rect 571812 274990 571840 277780
rect 571800 274984 571852 274990
rect 571800 274926 571852 274932
rect 573008 269929 573036 277780
rect 572994 269920 573050 269929
rect 572994 269855 573050 269864
rect 570696 266688 570748 266694
rect 570696 266630 570748 266636
rect 574204 266558 574232 277780
rect 575400 266626 575428 277780
rect 576596 272202 576624 277780
rect 576584 272196 576636 272202
rect 576584 272138 576636 272144
rect 575388 266620 575440 266626
rect 575388 266562 575440 266568
rect 574192 266552 574244 266558
rect 574192 266494 574244 266500
rect 577792 266121 577820 277780
rect 578896 274922 578924 277780
rect 578884 274916 578936 274922
rect 578884 274858 578936 274864
rect 580092 269550 580120 277780
rect 580080 269544 580132 269550
rect 580080 269486 580132 269492
rect 581288 266257 581316 277780
rect 582484 267617 582512 277780
rect 583680 272134 583708 277780
rect 583668 272128 583720 272134
rect 583668 272070 583720 272076
rect 584876 267753 584904 277780
rect 586072 275913 586100 277780
rect 586058 275904 586114 275913
rect 586058 275839 586114 275848
rect 587176 269482 587204 277780
rect 587164 269476 587216 269482
rect 587164 269418 587216 269424
rect 584862 267744 584918 267753
rect 584862 267679 584918 267688
rect 582470 267608 582526 267617
rect 582470 267543 582526 267552
rect 588372 266490 588400 277780
rect 589568 267481 589596 277780
rect 590764 272066 590792 277780
rect 590752 272060 590804 272066
rect 590752 272002 590804 272008
rect 589554 267472 589610 267481
rect 589554 267407 589610 267416
rect 591960 267345 591988 277780
rect 593156 275777 593184 277780
rect 593142 275768 593198 275777
rect 593142 275703 593198 275712
rect 594352 269793 594380 277780
rect 594338 269784 594394 269793
rect 594338 269719 594394 269728
rect 591946 267336 592002 267345
rect 591946 267271 592002 267280
rect 595456 267209 595484 277780
rect 595442 267200 595498 267209
rect 595442 267135 595498 267144
rect 588360 266484 588412 266490
rect 588360 266426 588412 266432
rect 596652 266422 596680 277780
rect 597848 272513 597876 277780
rect 597834 272504 597890 272513
rect 597834 272439 597890 272448
rect 599044 267073 599072 277780
rect 600240 275641 600268 277780
rect 600226 275632 600282 275641
rect 600226 275567 600282 275576
rect 601436 269414 601464 277780
rect 601424 269408 601476 269414
rect 601424 269350 601476 269356
rect 599030 267064 599086 267073
rect 599030 266999 599086 267008
rect 602540 266937 602568 277780
rect 602526 266928 602582 266937
rect 602526 266863 602582 266872
rect 596640 266416 596692 266422
rect 596640 266358 596692 266364
rect 603736 266354 603764 277780
rect 604932 271998 604960 277780
rect 604920 271992 604972 271998
rect 604920 271934 604972 271940
rect 606128 266801 606156 277780
rect 607324 275505 607352 277780
rect 607310 275496 607366 275505
rect 607310 275431 607366 275440
rect 608520 269346 608548 277780
rect 608508 269340 608560 269346
rect 608508 269282 608560 269288
rect 606114 266792 606170 266801
rect 606114 266727 606170 266736
rect 609716 266665 609744 277780
rect 610820 272814 610848 277780
rect 610808 272808 610860 272814
rect 610808 272750 610860 272756
rect 612016 272377 612044 277780
rect 612002 272368 612058 272377
rect 612002 272303 612058 272312
rect 609702 266656 609758 266665
rect 609702 266591 609758 266600
rect 613212 266529 613240 277780
rect 614408 275369 614436 277780
rect 614394 275360 614450 275369
rect 614394 275295 614450 275304
rect 615604 269278 615632 277780
rect 615592 269272 615644 269278
rect 615592 269214 615644 269220
rect 613198 266520 613254 266529
rect 613198 266455 613254 266464
rect 616800 266393 616828 277780
rect 617996 273086 618024 277780
rect 617984 273080 618036 273086
rect 617984 273022 618036 273028
rect 619100 271930 619128 277780
rect 620296 274854 620324 277780
rect 621492 275233 621520 277780
rect 621478 275224 621534 275233
rect 621478 275159 621534 275168
rect 620284 274848 620336 274854
rect 620284 274790 620336 274796
rect 619088 271924 619140 271930
rect 619088 271866 619140 271872
rect 622688 269657 622716 277780
rect 623884 274961 623912 277780
rect 623870 274952 623926 274961
rect 623870 274887 623926 274896
rect 625080 272746 625108 277780
rect 625068 272740 625120 272746
rect 625068 272682 625120 272688
rect 626184 272241 626212 277780
rect 627380 274786 627408 277780
rect 628576 275097 628604 277780
rect 628562 275088 628618 275097
rect 628562 275023 628618 275032
rect 627368 274780 627420 274786
rect 627368 274722 627420 274728
rect 626170 272232 626226 272241
rect 626170 272167 626226 272176
rect 622674 269648 622730 269657
rect 622674 269583 622730 269592
rect 629772 269521 629800 277780
rect 630968 274825 630996 277780
rect 630954 274816 631010 274825
rect 630954 274751 631010 274760
rect 632164 272542 632192 277780
rect 632152 272536 632204 272542
rect 632152 272478 632204 272484
rect 633360 271862 633388 277780
rect 634464 274718 634492 277780
rect 634452 274712 634504 274718
rect 635660 274689 635688 277780
rect 634452 274654 634504 274660
rect 635646 274680 635702 274689
rect 635646 274615 635702 274624
rect 633348 271856 633400 271862
rect 633348 271798 633400 271804
rect 629758 269512 629814 269521
rect 629758 269447 629814 269456
rect 636856 269385 636884 277780
rect 638052 274553 638080 277780
rect 638038 274544 638094 274553
rect 638038 274479 638094 274488
rect 639248 272338 639276 277780
rect 639236 272332 639288 272338
rect 639236 272274 639288 272280
rect 640444 272105 640472 277780
rect 641640 274650 641668 277780
rect 641628 274644 641680 274650
rect 641628 274586 641680 274592
rect 640430 272096 640486 272105
rect 640430 272031 640486 272040
rect 636842 269376 636898 269385
rect 636842 269311 636898 269320
rect 642744 269249 642772 277780
rect 642730 269240 642786 269249
rect 642730 269175 642786 269184
rect 643940 269113 643968 277780
rect 645136 271969 645164 277780
rect 645122 271960 645178 271969
rect 645122 271895 645178 271904
rect 646332 271833 646360 277780
rect 646318 271824 646374 271833
rect 646318 271759 646374 271768
rect 647528 269210 647556 277780
rect 647516 269204 647568 269210
rect 647516 269146 647568 269152
rect 648724 269142 648752 277780
rect 648712 269136 648764 269142
rect 643926 269104 643982 269113
rect 648712 269078 648764 269084
rect 643926 269039 643982 269048
rect 616786 266384 616842 266393
rect 603724 266348 603776 266354
rect 616786 266319 616842 266328
rect 603724 266290 603776 266296
rect 581274 266248 581330 266257
rect 581274 266183 581330 266192
rect 577778 266112 577834 266121
rect 577778 266047 577834 266056
rect 511632 265804 511684 265810
rect 511632 265746 511684 265752
rect 498844 265668 498896 265674
rect 498844 265610 498896 265616
rect 471980 265328 472032 265334
rect 471980 265270 472032 265276
rect 418066 262712 418122 262721
rect 418066 262647 418122 262656
rect 418080 262274 418108 262647
rect 418068 262268 418120 262274
rect 418068 262210 418120 262216
rect 571708 262268 571760 262274
rect 571708 262210 571760 262216
rect 417790 260264 417846 260273
rect 417790 260199 417846 260208
rect 184938 259992 184994 260001
rect 184938 259927 184994 259936
rect 184952 259486 184980 259927
rect 417804 259486 417832 260199
rect 184940 259480 184992 259486
rect 184940 259422 184992 259428
rect 417792 259480 417844 259486
rect 417792 259422 417844 259428
rect 418342 257952 418398 257961
rect 418342 257887 418398 257896
rect 418356 256766 418384 257887
rect 418344 256760 418396 256766
rect 418344 256702 418396 256708
rect 571524 256760 571576 256766
rect 571524 256702 571576 256708
rect 416778 255504 416834 255513
rect 416778 255439 416834 255448
rect 416792 253978 416820 255439
rect 416780 253972 416832 253978
rect 416780 253914 416832 253920
rect 416778 253192 416834 253201
rect 416778 253127 416834 253136
rect 184938 251968 184994 251977
rect 184938 251903 184994 251912
rect 184952 251258 184980 251903
rect 416792 251258 416820 253127
rect 184940 251252 184992 251258
rect 184940 251194 184992 251200
rect 416780 251252 416832 251258
rect 416780 251194 416832 251200
rect 416778 250744 416834 250753
rect 416778 250679 416834 250688
rect 416792 248470 416820 250679
rect 416780 248464 416832 248470
rect 416780 248406 416832 248412
rect 569868 248464 569920 248470
rect 569868 248406 569920 248412
rect 418066 248296 418122 248305
rect 418066 248231 418122 248240
rect 184938 244080 184994 244089
rect 184938 244015 184994 244024
rect 184952 242962 184980 244015
rect 184940 242956 184992 242962
rect 184940 242898 184992 242904
rect 161388 237380 161440 237386
rect 161388 237322 161440 237328
rect 142160 237244 142212 237250
rect 142160 237186 142212 237192
rect 106186 237008 106242 237017
rect 106186 236943 106242 236952
rect 136548 236972 136600 236978
rect 89626 236872 89682 236881
rect 89626 236807 89682 236816
rect 81346 236464 81402 236473
rect 81346 236399 81402 236408
rect 73066 236328 73122 236337
rect 73066 236263 73122 236272
rect 67548 236088 67600 236094
rect 67548 236030 67600 236036
rect 62026 235920 62082 235929
rect 62026 235855 62082 235864
rect 61936 227860 61988 227866
rect 61936 227802 61988 227808
rect 60280 225004 60332 225010
rect 60280 224946 60332 224952
rect 60292 217410 60320 224946
rect 61106 222184 61162 222193
rect 61106 222119 61162 222128
rect 61120 217410 61148 222119
rect 61948 217410 61976 227802
rect 62040 221406 62068 235855
rect 66996 225072 67048 225078
rect 63406 225040 63462 225049
rect 66996 225014 67048 225020
rect 63406 224975 63462 224984
rect 62764 222760 62816 222766
rect 62764 222702 62816 222708
rect 62028 221400 62080 221406
rect 62028 221342 62080 221348
rect 62776 217410 62804 222702
rect 63420 217410 63448 224975
rect 65340 222964 65392 222970
rect 65340 222906 65392 222912
rect 64512 220992 64564 220998
rect 64512 220934 64564 220940
rect 64524 217410 64552 220934
rect 65352 217410 65380 222906
rect 66166 222320 66222 222329
rect 66166 222255 66222 222264
rect 66180 217410 66208 222255
rect 67008 217410 67036 225014
rect 67560 221338 67588 236030
rect 70398 225176 70454 225185
rect 70398 225111 70454 225120
rect 67822 222456 67878 222465
rect 67822 222391 67878 222400
rect 67548 221332 67600 221338
rect 67548 221274 67600 221280
rect 67836 217410 67864 222391
rect 68652 221060 68704 221066
rect 68652 221002 68704 221008
rect 68664 217410 68692 221002
rect 69480 220924 69532 220930
rect 69480 220866 69532 220872
rect 69492 217410 69520 220866
rect 70412 217410 70440 225111
rect 72056 223100 72108 223106
rect 72056 223042 72108 223048
rect 71228 222692 71280 222698
rect 71228 222634 71280 222640
rect 71240 217410 71268 222634
rect 72068 217410 72096 223042
rect 72882 222728 72938 222737
rect 72882 222663 72938 222672
rect 72896 217410 72924 222663
rect 73080 222426 73108 236263
rect 75826 236192 75882 236201
rect 75826 236127 75882 236136
rect 73160 236020 73212 236026
rect 73160 235962 73212 235968
rect 73068 222420 73120 222426
rect 73068 222362 73120 222368
rect 73172 220930 73200 235962
rect 73712 225140 73764 225146
rect 73712 225082 73764 225088
rect 73160 220924 73212 220930
rect 73160 220866 73212 220872
rect 73724 217410 73752 225082
rect 74446 222592 74502 222601
rect 74446 222527 74502 222536
rect 74460 217410 74488 222527
rect 75368 222420 75420 222426
rect 75368 222362 75420 222368
rect 75380 217410 75408 222362
rect 75840 220998 75868 236127
rect 78586 236056 78642 236065
rect 78586 235991 78642 236000
rect 77114 225312 77170 225321
rect 77114 225247 77170 225256
rect 76288 221400 76340 221406
rect 76288 221342 76340 221348
rect 75828 220992 75880 220998
rect 75828 220934 75880 220940
rect 76300 217410 76328 221342
rect 77128 217410 77156 225247
rect 78600 221406 78628 235991
rect 80426 225448 80482 225457
rect 80426 225383 80482 225392
rect 78772 223236 78824 223242
rect 78772 223178 78824 223184
rect 78588 221400 78640 221406
rect 78588 221342 78640 221348
rect 77944 221332 77996 221338
rect 77944 221274 77996 221280
rect 77956 217410 77984 221274
rect 78784 217410 78812 223178
rect 79598 222864 79654 222873
rect 79598 222799 79654 222808
rect 79612 217410 79640 222799
rect 80440 217410 80468 225383
rect 81360 222698 81388 236399
rect 86868 236156 86920 236162
rect 86868 236098 86920 236104
rect 83830 225584 83886 225593
rect 83830 225519 83886 225528
rect 82728 222896 82780 222902
rect 82728 222838 82780 222844
rect 81348 222692 81400 222698
rect 81348 222634 81400 222640
rect 82176 222624 82228 222630
rect 82176 222566 82228 222572
rect 81256 222488 81308 222494
rect 81256 222430 81308 222436
rect 81268 217410 81296 222430
rect 82188 217410 82216 222566
rect 82740 217410 82768 222838
rect 83844 217410 83872 225519
rect 86316 223372 86368 223378
rect 86316 223314 86368 223320
rect 85488 222556 85540 222562
rect 85488 222498 85540 222504
rect 84660 221264 84712 221270
rect 84660 221206 84712 221212
rect 84672 217410 84700 221206
rect 85500 217410 85528 222498
rect 86328 217410 86356 223314
rect 86880 221338 86908 236098
rect 87144 227996 87196 228002
rect 87144 227938 87196 227944
rect 86868 221332 86920 221338
rect 86868 221274 86920 221280
rect 87156 217410 87184 227938
rect 88890 225856 88946 225865
rect 88890 225791 88946 225800
rect 88064 223032 88116 223038
rect 88064 222974 88116 222980
rect 88076 217410 88104 222974
rect 88904 217410 88932 225791
rect 89640 222766 89668 236807
rect 97906 236736 97962 236745
rect 97906 236671 97962 236680
rect 95146 236600 95202 236609
rect 95146 236535 95202 236544
rect 93768 228064 93820 228070
rect 93768 228006 93820 228012
rect 90548 227928 90600 227934
rect 90548 227870 90600 227876
rect 89628 222760 89680 222766
rect 89628 222702 89680 222708
rect 89720 222692 89772 222698
rect 89720 222634 89772 222640
rect 89732 217410 89760 222634
rect 90560 217410 90588 227870
rect 92202 225720 92258 225729
rect 92202 225655 92258 225664
rect 91376 220924 91428 220930
rect 91376 220866 91428 220872
rect 91388 217410 91416 220866
rect 92216 217410 92244 225655
rect 93032 221944 93084 221950
rect 93032 221886 93084 221892
rect 93044 217410 93072 221886
rect 93780 217410 93808 228006
rect 94780 223168 94832 223174
rect 94780 223110 94832 223116
rect 94792 217410 94820 223110
rect 95160 221270 95188 236535
rect 97264 228132 97316 228138
rect 97264 228074 97316 228080
rect 95608 225208 95660 225214
rect 95608 225150 95660 225156
rect 95148 221264 95200 221270
rect 95148 221206 95200 221212
rect 95620 217410 95648 225150
rect 96434 223000 96490 223009
rect 96434 222935 96490 222944
rect 96448 217410 96476 222935
rect 97276 217410 97304 228074
rect 97920 222902 97948 236671
rect 103428 236292 103480 236298
rect 103428 236234 103480 236240
rect 102046 226128 102102 226137
rect 102046 226063 102102 226072
rect 98918 225992 98974 226001
rect 98918 225927 98974 225936
rect 97908 222896 97960 222902
rect 97908 222838 97960 222844
rect 98092 222828 98144 222834
rect 98092 222770 98144 222776
rect 98104 217410 98132 222770
rect 98932 217410 98960 225927
rect 100668 225344 100720 225350
rect 100668 225286 100720 225292
rect 99840 221740 99892 221746
rect 99840 221682 99892 221688
rect 99852 217410 99880 221682
rect 100680 217410 100708 225286
rect 101496 223304 101548 223310
rect 101496 223246 101548 223252
rect 101508 217410 101536 223246
rect 102060 217410 102088 226063
rect 103440 222970 103468 236234
rect 105728 225480 105780 225486
rect 105728 225422 105780 225428
rect 103980 225276 104032 225282
rect 103980 225218 104032 225224
rect 103428 222964 103480 222970
rect 103428 222906 103480 222912
rect 103152 222896 103204 222902
rect 103152 222838 103204 222844
rect 103164 217410 103192 222838
rect 103992 217410 104020 225218
rect 104806 223136 104862 223145
rect 104806 223071 104862 223080
rect 104820 217410 104848 223071
rect 105740 217410 105768 225422
rect 106200 223038 106228 236943
rect 136548 236914 136600 236920
rect 128268 236904 128320 236910
rect 128268 236846 128320 236852
rect 117228 236700 117280 236706
rect 117228 236642 117280 236648
rect 111708 236224 111760 236230
rect 111708 236166 111760 236172
rect 110696 225752 110748 225758
rect 110696 225694 110748 225700
rect 109040 225548 109092 225554
rect 109040 225490 109092 225496
rect 107384 225412 107436 225418
rect 107384 225354 107436 225360
rect 106556 223440 106608 223446
rect 106556 223382 106608 223388
rect 106188 223032 106240 223038
rect 106188 222974 106240 222980
rect 106568 217410 106596 223382
rect 107396 217410 107424 225354
rect 108212 223508 108264 223514
rect 108212 223450 108264 223456
rect 108224 217410 108252 223450
rect 109052 217410 109080 225490
rect 109868 222964 109920 222970
rect 109868 222906 109920 222912
rect 109880 217410 109908 222906
rect 110708 217410 110736 225694
rect 111614 223272 111670 223281
rect 111614 223207 111670 223216
rect 111628 217410 111656 223207
rect 111720 223174 111748 236166
rect 114100 225956 114152 225962
rect 114100 225898 114152 225904
rect 112444 225616 112496 225622
rect 112444 225558 112496 225564
rect 111708 223168 111760 223174
rect 111708 223110 111760 223116
rect 112456 217410 112484 225558
rect 113088 223576 113140 223582
rect 113088 223518 113140 223524
rect 113100 217410 113128 223518
rect 114112 217410 114140 225898
rect 115756 225684 115808 225690
rect 115756 225626 115808 225632
rect 114928 222148 114980 222154
rect 114928 222090 114980 222096
rect 114940 217410 114968 222090
rect 115768 217410 115796 225626
rect 116584 223168 116636 223174
rect 116584 223110 116636 223116
rect 116596 217410 116624 223110
rect 117240 223106 117268 236642
rect 119988 236496 120040 236502
rect 119988 236438 120040 236444
rect 119160 228200 119212 228206
rect 119160 228142 119212 228148
rect 117504 225888 117556 225894
rect 117504 225830 117556 225836
rect 117228 223100 117280 223106
rect 117228 223042 117280 223048
rect 117516 217410 117544 225830
rect 118332 223032 118384 223038
rect 118332 222974 118384 222980
rect 118344 217410 118372 222974
rect 119172 217410 119200 228142
rect 120000 223242 120028 236438
rect 125508 236428 125560 236434
rect 125508 236370 125560 236376
rect 122748 236360 122800 236366
rect 122748 236302 122800 236308
rect 122472 228268 122524 228274
rect 122472 228210 122524 228216
rect 120816 225820 120868 225826
rect 120816 225762 120868 225768
rect 119988 223236 120040 223242
rect 119988 223178 120040 223184
rect 119988 223100 120040 223106
rect 119988 223042 120040 223048
rect 120000 217410 120028 223042
rect 120828 217410 120856 225762
rect 121366 223408 121422 223417
rect 121366 223343 121422 223352
rect 121380 217410 121408 223343
rect 122484 217410 122512 228210
rect 122760 223310 122788 236302
rect 124128 226024 124180 226030
rect 124128 225966 124180 225972
rect 122748 223304 122800 223310
rect 122748 223246 122800 223252
rect 123392 221876 123444 221882
rect 123392 221818 123444 221824
rect 123404 217410 123432 221818
rect 124140 217410 124168 225966
rect 125520 223446 125548 236370
rect 125876 228336 125928 228342
rect 125876 228278 125928 228284
rect 125508 223440 125560 223446
rect 125508 223382 125560 223388
rect 125048 221808 125100 221814
rect 125048 221750 125100 221756
rect 125060 217410 125088 221750
rect 125888 217410 125916 228278
rect 127532 226092 127584 226098
rect 127532 226034 127584 226040
rect 126704 223236 126756 223242
rect 126704 223178 126756 223184
rect 126716 217410 126744 223178
rect 127544 217410 127572 226034
rect 128280 223378 128308 236846
rect 135996 228540 136048 228546
rect 135996 228482 136048 228488
rect 132408 228472 132460 228478
rect 132408 228414 132460 228420
rect 129280 228404 129332 228410
rect 129280 228346 129332 228352
rect 128268 223372 128320 223378
rect 128268 223314 128320 223320
rect 128360 223304 128412 223310
rect 128360 223246 128412 223252
rect 128372 217410 128400 223246
rect 129292 217410 129320 228346
rect 130936 226160 130988 226166
rect 130936 226102 130988 226108
rect 130108 221672 130160 221678
rect 130108 221614 130160 221620
rect 130120 217410 130148 221614
rect 130948 217410 130976 226102
rect 131764 221332 131816 221338
rect 131764 221274 131816 221280
rect 131776 217410 131804 221274
rect 132420 217410 132448 228414
rect 134248 226228 134300 226234
rect 134248 226170 134300 226176
rect 133420 220856 133472 220862
rect 133420 220798 133472 220804
rect 133432 217410 133460 220798
rect 134260 217410 134288 226170
rect 135168 223440 135220 223446
rect 135168 223382 135220 223388
rect 135180 217410 135208 223382
rect 136008 217410 136036 228482
rect 136560 223514 136588 236914
rect 139308 236768 139360 236774
rect 139308 236710 139360 236716
rect 139216 228608 139268 228614
rect 139216 228550 139268 228556
rect 137652 226296 137704 226302
rect 137652 226238 137704 226244
rect 136548 223508 136600 223514
rect 136548 223450 136600 223456
rect 136824 221536 136876 221542
rect 136824 221478 136876 221484
rect 136836 217410 136864 221478
rect 137664 217410 137692 226238
rect 138480 221400 138532 221406
rect 138480 221342 138532 221348
rect 138492 217410 138520 221342
rect 139228 217410 139256 228550
rect 139320 223582 139348 236710
rect 142068 236564 142120 236570
rect 142068 236506 142120 236512
rect 141056 224868 141108 224874
rect 141056 224810 141108 224816
rect 139308 223576 139360 223582
rect 139308 223518 139360 223524
rect 140136 223508 140188 223514
rect 140136 223450 140188 223456
rect 140148 217410 140176 223450
rect 141068 217410 141096 224810
rect 141884 223576 141936 223582
rect 141884 223518 141936 223524
rect 141896 217410 141924 223518
rect 142080 221338 142108 236506
rect 142172 222154 142200 237186
rect 159824 237176 159876 237182
rect 153106 237144 153162 237153
rect 159824 237118 159876 237124
rect 153106 237079 153162 237088
rect 153200 237108 153252 237114
rect 147588 237040 147640 237046
rect 147588 236982 147640 236988
rect 146024 228744 146076 228750
rect 146024 228686 146076 228692
rect 142712 228676 142764 228682
rect 142712 228618 142764 228624
rect 142160 222148 142212 222154
rect 142160 222090 142212 222096
rect 142068 221332 142120 221338
rect 142068 221274 142120 221280
rect 142724 217410 142752 228618
rect 144368 224800 144420 224806
rect 144368 224742 144420 224748
rect 143448 221604 143500 221610
rect 143448 221546 143500 221552
rect 143460 217410 143488 221546
rect 144380 217410 144408 224742
rect 145196 221332 145248 221338
rect 145196 221274 145248 221280
rect 145208 217410 145236 221274
rect 146036 217410 146064 228686
rect 146944 222080 146996 222086
rect 146944 222022 146996 222028
rect 146956 217410 146984 222022
rect 147600 221406 147628 236982
rect 150348 236632 150400 236638
rect 150348 236574 150400 236580
rect 149428 228812 149480 228818
rect 149428 228754 149480 228760
rect 147772 224732 147824 224738
rect 147772 224674 147824 224680
rect 147588 221400 147640 221406
rect 147588 221342 147640 221348
rect 147784 217410 147812 224674
rect 148600 222148 148652 222154
rect 148600 222090 148652 222096
rect 148612 217410 148640 222090
rect 149440 217410 149468 228754
rect 150360 221406 150388 236574
rect 152832 228880 152884 228886
rect 152832 228822 152884 228828
rect 151084 224596 151136 224602
rect 151084 224538 151136 224544
rect 150348 221400 150400 221406
rect 150348 221342 150400 221348
rect 150256 221332 150308 221338
rect 150256 221274 150308 221280
rect 150268 217410 150296 221274
rect 151096 217410 151124 224538
rect 151728 221400 151780 221406
rect 151728 221342 151780 221348
rect 151740 217410 151768 221342
rect 152844 217410 152872 228822
rect 153120 221950 153148 237079
rect 153200 237050 153252 237056
rect 153108 221944 153160 221950
rect 153108 221886 153160 221892
rect 153212 221338 153240 237050
rect 155868 236836 155920 236842
rect 155868 236778 155920 236784
rect 154488 224664 154540 224670
rect 154488 224606 154540 224612
rect 153660 222012 153712 222018
rect 153660 221954 153712 221960
rect 153200 221332 153252 221338
rect 153200 221274 153252 221280
rect 153672 217410 153700 221954
rect 154500 217410 154528 224606
rect 155316 221944 155368 221950
rect 155316 221886 155368 221892
rect 155328 217410 155356 221886
rect 155880 221406 155908 236778
rect 158628 235612 158680 235618
rect 158628 235554 158680 235560
rect 155960 235544 156012 235550
rect 155960 235486 156012 235492
rect 155972 221882 156000 235486
rect 156052 235408 156104 235414
rect 156052 235350 156104 235356
rect 155960 221876 156012 221882
rect 155960 221818 156012 221824
rect 156064 221814 156092 235350
rect 156144 228948 156196 228954
rect 156144 228890 156196 228896
rect 156052 221808 156104 221814
rect 156052 221750 156104 221756
rect 155868 221400 155920 221406
rect 155868 221342 155920 221348
rect 156156 217410 156184 228890
rect 157800 224460 157852 224466
rect 157800 224402 157852 224408
rect 156972 221332 157024 221338
rect 156972 221274 157024 221280
rect 156984 217410 157012 221274
rect 157812 217410 157840 224402
rect 158640 221678 158668 235554
rect 159548 229016 159600 229022
rect 159548 228958 159600 228964
rect 158628 221672 158680 221678
rect 158628 221614 158680 221620
rect 158720 221400 158772 221406
rect 158720 221342 158772 221348
rect 158732 217410 158760 221342
rect 159560 217410 159588 228958
rect 159836 221406 159864 237118
rect 161204 224528 161256 224534
rect 161204 224470 161256 224476
rect 160376 221876 160428 221882
rect 160376 221818 160428 221824
rect 159824 221400 159876 221406
rect 159824 221342 159876 221348
rect 160388 217410 160416 221818
rect 161216 217410 161244 224470
rect 161400 221338 161428 237322
rect 165436 237312 165488 237318
rect 165436 237254 165488 237260
rect 165344 235884 165396 235890
rect 165344 235826 165396 235832
rect 161572 235476 161624 235482
rect 161572 235418 161624 235424
rect 161480 235000 161532 235006
rect 161480 234942 161532 234948
rect 161492 221746 161520 234942
rect 161480 221740 161532 221746
rect 161480 221682 161532 221688
rect 161584 221542 161612 235418
rect 162768 230580 162820 230586
rect 162768 230522 162820 230528
rect 162032 221808 162084 221814
rect 162032 221750 162084 221756
rect 161572 221536 161624 221542
rect 161572 221478 161624 221484
rect 161388 221332 161440 221338
rect 161388 221274 161440 221280
rect 162044 217410 162072 221750
rect 162780 217410 162808 230522
rect 164608 224392 164660 224398
rect 164608 224334 164660 224340
rect 163688 221400 163740 221406
rect 163688 221342 163740 221348
rect 163700 217410 163728 221342
rect 164620 217410 164648 224334
rect 165356 221406 165384 235826
rect 165344 221400 165396 221406
rect 165344 221342 165396 221348
rect 165448 217410 165476 237254
rect 168104 235952 168156 235958
rect 168104 235894 168156 235900
rect 166264 230716 166316 230722
rect 166264 230658 166316 230664
rect 166276 217410 166304 230658
rect 167920 224324 167972 224330
rect 167920 224266 167972 224272
rect 167092 221332 167144 221338
rect 167092 221274 167144 221280
rect 167104 217410 167132 221274
rect 167932 217410 167960 224266
rect 168116 221338 168144 235894
rect 173716 235816 173768 235822
rect 173716 235758 173768 235764
rect 169668 235136 169720 235142
rect 169668 235078 169720 235084
rect 169576 230648 169628 230654
rect 169576 230590 169628 230596
rect 168748 221672 168800 221678
rect 168748 221614 168800 221620
rect 168104 221332 168156 221338
rect 168104 221274 168156 221280
rect 168760 217410 168788 221614
rect 169588 217410 169616 230590
rect 169680 221610 169708 235078
rect 172980 230852 173032 230858
rect 172980 230794 173032 230800
rect 171048 224256 171100 224262
rect 171048 224198 171100 224204
rect 170496 221740 170548 221746
rect 170496 221682 170548 221688
rect 169668 221604 169720 221610
rect 169668 221546 169720 221552
rect 170508 217410 170536 221682
rect 171060 217410 171088 224198
rect 172152 221400 172204 221406
rect 172152 221342 172204 221348
rect 172164 217410 172192 221342
rect 172992 217410 173020 230794
rect 173728 217410 173756 235758
rect 173808 235748 173860 235754
rect 173808 235690 173860 235696
rect 173820 221406 173848 235690
rect 183468 235340 183520 235346
rect 183468 235282 183520 235288
rect 179328 235068 179380 235074
rect 179328 235010 179380 235016
rect 176384 230784 176436 230790
rect 176384 230726 176436 230732
rect 174636 224188 174688 224194
rect 174636 224130 174688 224136
rect 173808 221400 173860 221406
rect 173808 221342 173860 221348
rect 174648 217410 174676 224130
rect 175464 221604 175516 221610
rect 175464 221546 175516 221552
rect 175476 217410 175504 221546
rect 176396 217410 176424 230726
rect 178040 224120 178092 224126
rect 178040 224062 178092 224068
rect 177212 221536 177264 221542
rect 177212 221478 177264 221484
rect 177224 217410 177252 221478
rect 178052 217410 178080 224062
rect 179340 221338 179368 235010
rect 179696 230988 179748 230994
rect 179696 230930 179748 230936
rect 178868 221332 178920 221338
rect 178868 221274 178920 221280
rect 179328 221332 179380 221338
rect 179328 221274 179380 221280
rect 178880 217410 178908 221274
rect 179708 217410 179736 230930
rect 183100 230920 183152 230926
rect 183100 230862 183152 230868
rect 181352 224052 181404 224058
rect 181352 223994 181404 224000
rect 180524 221060 180576 221066
rect 180524 221002 180576 221008
rect 180536 217410 180564 221002
rect 181364 217410 181392 223994
rect 182088 221468 182140 221474
rect 182088 221410 182140 221416
rect 182100 217410 182128 221410
rect 183112 217410 183140 230862
rect 183480 221066 183508 235282
rect 190368 235272 190420 235278
rect 190368 235214 190420 235220
rect 187608 235204 187660 235210
rect 187608 235146 187660 235152
rect 186412 231056 186464 231062
rect 186412 230998 186464 231004
rect 184756 223984 184808 223990
rect 184756 223926 184808 223932
rect 183928 221400 183980 221406
rect 183928 221342 183980 221348
rect 183468 221060 183520 221066
rect 183468 221002 183520 221008
rect 183940 217410 183968 221342
rect 184768 217410 184796 223926
rect 185584 221332 185636 221338
rect 185584 221274 185636 221280
rect 185596 217410 185624 221274
rect 186424 217410 186452 230998
rect 187620 221338 187648 235146
rect 188160 223916 188212 223922
rect 188160 223858 188212 223864
rect 187608 221332 187660 221338
rect 187608 221274 187660 221280
rect 187240 221264 187292 221270
rect 187240 221206 187292 221212
rect 187252 217410 187280 221206
rect 188172 217410 188200 223858
rect 189540 222760 189592 222766
rect 189540 222702 189592 222708
rect 189552 222562 189580 222702
rect 189540 222556 189592 222562
rect 189540 222498 189592 222504
rect 189724 222488 189776 222494
rect 189724 222430 189776 222436
rect 188988 221060 189040 221066
rect 188988 221002 189040 221008
rect 189000 217410 189028 221002
rect 189736 220930 189764 222430
rect 189724 220924 189776 220930
rect 189724 220866 189776 220872
rect 189816 220924 189868 220930
rect 189816 220866 189868 220872
rect 189828 217410 189856 220866
rect 190380 217410 190408 235214
rect 190644 233028 190696 233034
rect 190644 232970 190696 232976
rect 190656 224942 190684 232970
rect 192312 227730 192340 239700
rect 192404 239686 192602 239714
rect 192404 233034 192432 239686
rect 192956 236094 192984 239700
rect 192944 236088 192996 236094
rect 192944 236030 192996 236036
rect 193036 236088 193088 236094
rect 193036 236030 193088 236036
rect 193048 235090 193076 236030
rect 192956 235062 193076 235090
rect 192392 233028 192444 233034
rect 192392 232970 192444 232976
rect 192300 227724 192352 227730
rect 192300 227666 192352 227672
rect 190644 224936 190696 224942
rect 190644 224878 190696 224884
rect 191472 224936 191524 224942
rect 191472 224878 191524 224884
rect 191484 217410 191512 224878
rect 192956 221338 192984 235062
rect 193036 234932 193088 234938
rect 193036 234874 193088 234880
rect 192300 221332 192352 221338
rect 192300 221274 192352 221280
rect 192944 221332 192996 221338
rect 192944 221274 192996 221280
rect 192312 217410 192340 221274
rect 193048 217410 193076 234874
rect 193324 222222 193352 239700
rect 193416 239686 193706 239714
rect 193416 224913 193444 239686
rect 193680 233096 193732 233102
rect 193680 233038 193732 233044
rect 193496 233028 193548 233034
rect 193496 232970 193548 232976
rect 193508 225010 193536 232970
rect 193496 225004 193548 225010
rect 193496 224946 193548 224952
rect 193402 224904 193458 224913
rect 193402 224839 193458 224848
rect 193312 222216 193364 222222
rect 193312 222158 193364 222164
rect 193692 221202 193720 233038
rect 194060 227798 194088 239700
rect 194428 236337 194456 239700
rect 194414 236328 194470 236337
rect 194414 236263 194470 236272
rect 194796 235929 194824 239700
rect 194888 239686 195178 239714
rect 194782 235920 194838 235929
rect 194782 235855 194838 235864
rect 194888 233034 194916 239686
rect 194876 233028 194928 233034
rect 194876 232970 194928 232976
rect 195440 227866 195468 239700
rect 195532 239686 195822 239714
rect 196190 239686 196388 239714
rect 196558 239686 196664 239714
rect 195532 233102 195560 239686
rect 196360 233186 196388 239686
rect 196360 233158 196572 233186
rect 195520 233096 195572 233102
rect 195520 233038 195572 233044
rect 196164 233096 196216 233102
rect 196164 233038 196216 233044
rect 195428 227860 195480 227866
rect 195428 227802 195480 227808
rect 194048 227792 194100 227798
rect 194048 227734 194100 227740
rect 194876 225004 194928 225010
rect 194876 224946 194928 224952
rect 194048 222284 194100 222290
rect 194048 222226 194100 222232
rect 193680 221196 193732 221202
rect 193680 221138 193732 221144
rect 194060 217410 194088 222226
rect 194888 217410 194916 224946
rect 196176 222329 196204 233038
rect 196348 233028 196400 233034
rect 196348 232970 196400 232976
rect 196256 232892 196308 232898
rect 196256 232834 196308 232840
rect 196268 225049 196296 232834
rect 196254 225040 196310 225049
rect 196254 224975 196310 224984
rect 196162 222320 196218 222329
rect 196162 222255 196218 222264
rect 195704 222216 195756 222222
rect 195704 222158 195756 222164
rect 195716 217410 195744 222158
rect 196360 221134 196388 232970
rect 196440 232960 196492 232966
rect 196440 232902 196492 232908
rect 196452 225078 196480 232902
rect 196440 225072 196492 225078
rect 196440 225014 196492 225020
rect 196544 222193 196572 233158
rect 196636 232898 196664 239686
rect 196912 236298 196940 239700
rect 197004 239686 197294 239714
rect 197004 236881 197032 239686
rect 197268 236904 197320 236910
rect 196990 236872 197046 236881
rect 197268 236846 197320 236852
rect 196990 236807 197046 236816
rect 196900 236292 196952 236298
rect 196900 236234 196952 236240
rect 197280 236230 197308 236846
rect 197176 236224 197228 236230
rect 197176 236166 197228 236172
rect 197268 236224 197320 236230
rect 197648 236201 197676 239700
rect 197740 239686 198030 239714
rect 198108 239686 198306 239714
rect 198384 239686 198674 239714
rect 198752 239686 199042 239714
rect 199120 239686 199410 239714
rect 197268 236166 197320 236172
rect 197634 236192 197690 236201
rect 197188 234734 197216 236166
rect 197634 236127 197690 236136
rect 197268 235680 197320 235686
rect 197268 235622 197320 235628
rect 197280 235074 197308 235622
rect 197268 235068 197320 235074
rect 197268 235010 197320 235016
rect 197176 234728 197228 234734
rect 197176 234670 197228 234676
rect 197740 232966 197768 239686
rect 198108 233034 198136 239686
rect 198384 233102 198412 239686
rect 198648 234932 198700 234938
rect 198648 234874 198700 234880
rect 198372 233096 198424 233102
rect 198372 233038 198424 233044
rect 198096 233028 198148 233034
rect 198096 232970 198148 232976
rect 197728 232960 197780 232966
rect 197728 232902 197780 232908
rect 196624 232892 196676 232898
rect 196624 232834 196676 232840
rect 198188 225072 198240 225078
rect 198188 225014 198240 225020
rect 196530 222184 196586 222193
rect 196530 222119 196586 222128
rect 196532 221332 196584 221338
rect 196532 221274 196584 221280
rect 196348 221128 196400 221134
rect 196348 221070 196400 221076
rect 196544 217410 196572 221274
rect 197360 220992 197412 220998
rect 197360 220934 197412 220940
rect 197372 217410 197400 220934
rect 198200 217410 198228 225014
rect 198660 220998 198688 234874
rect 198752 222465 198780 239686
rect 199120 225185 199148 239686
rect 199764 236706 199792 239700
rect 199752 236700 199804 236706
rect 199752 236642 199804 236648
rect 200132 236026 200160 239700
rect 200500 236473 200528 239700
rect 200592 239686 200882 239714
rect 200960 239686 201158 239714
rect 201526 239686 201724 239714
rect 200486 236464 200542 236473
rect 200486 236399 200542 236408
rect 200120 236020 200172 236026
rect 200120 235962 200172 235968
rect 199106 225176 199162 225185
rect 200592 225146 200620 239686
rect 200856 236700 200908 236706
rect 200856 236642 200908 236648
rect 199106 225111 199162 225120
rect 200580 225140 200632 225146
rect 200580 225082 200632 225088
rect 198844 223378 199056 223394
rect 198844 223372 199068 223378
rect 198844 223366 199016 223372
rect 198844 223242 198872 223366
rect 199016 223314 199068 223320
rect 198832 223236 198884 223242
rect 198832 223178 198884 223184
rect 198924 223236 198976 223242
rect 198924 223178 198976 223184
rect 198936 222970 198964 223178
rect 198924 222964 198976 222970
rect 198924 222906 198976 222912
rect 199016 222964 199068 222970
rect 199016 222906 199068 222912
rect 198738 222456 198794 222465
rect 198738 222391 198794 222400
rect 198648 220992 198700 220998
rect 198648 220934 198700 220940
rect 199028 217410 199056 222906
rect 200868 221338 200896 236642
rect 200960 222426 200988 239686
rect 201408 236020 201460 236026
rect 201408 235962 201460 235968
rect 201316 225140 201368 225146
rect 201316 225082 201368 225088
rect 200948 222420 201000 222426
rect 200948 222362 201000 222368
rect 200856 221332 200908 221338
rect 200856 221274 200908 221280
rect 200764 221196 200816 221202
rect 200764 221138 200816 221144
rect 199936 221128 199988 221134
rect 199936 221070 199988 221076
rect 199948 217410 199976 221070
rect 200776 217410 200804 221138
rect 201328 217410 201356 225082
rect 201420 222970 201448 235962
rect 201408 222964 201460 222970
rect 201408 222906 201460 222912
rect 201696 222737 201724 239686
rect 201682 222728 201738 222737
rect 201682 222663 201738 222672
rect 201880 222601 201908 239700
rect 202064 239686 202262 239714
rect 202064 225321 202092 239686
rect 202616 236502 202644 239700
rect 202604 236496 202656 236502
rect 202604 236438 202656 236444
rect 202984 236065 203012 239700
rect 203248 236496 203300 236502
rect 203248 236438 203300 236444
rect 202970 236056 203026 236065
rect 202970 235991 203026 236000
rect 202050 225312 202106 225321
rect 202050 225247 202106 225256
rect 201866 222592 201922 222601
rect 201866 222527 201922 222536
rect 202420 222352 202472 222358
rect 202420 222294 202472 222300
rect 202432 217410 202460 222294
rect 203260 217410 203288 236438
rect 203352 236162 203380 239700
rect 203444 239686 203734 239714
rect 203812 239686 204010 239714
rect 203340 236156 203392 236162
rect 203340 236098 203392 236104
rect 203444 225457 203472 239686
rect 203430 225448 203486 225457
rect 203430 225383 203486 225392
rect 203812 222630 203840 239686
rect 204168 236156 204220 236162
rect 204168 236098 204220 236104
rect 203800 222624 203852 222630
rect 203800 222566 203852 222572
rect 204180 217410 204208 236098
rect 204364 222873 204392 239700
rect 204456 239686 204746 239714
rect 204824 239686 205114 239714
rect 205192 239686 205482 239714
rect 204350 222864 204406 222873
rect 204350 222799 204406 222808
rect 204456 222562 204484 239686
rect 204824 225593 204852 239686
rect 204904 227792 204956 227798
rect 204904 227734 204956 227740
rect 204810 225584 204866 225593
rect 204810 225519 204866 225528
rect 204444 222556 204496 222562
rect 204444 222498 204496 222504
rect 204916 217410 204944 227734
rect 205192 222766 205220 239686
rect 205836 236745 205864 239700
rect 205822 236736 205878 236745
rect 205822 236671 205878 236680
rect 206204 236609 206232 239700
rect 206376 236904 206428 236910
rect 206376 236846 206428 236852
rect 206190 236600 206246 236609
rect 206388 236570 206416 236846
rect 206190 236535 206246 236544
rect 206376 236564 206428 236570
rect 206376 236506 206428 236512
rect 205732 236292 205784 236298
rect 205732 236234 205784 236240
rect 205744 234938 205772 236234
rect 205732 234932 205784 234938
rect 205732 234874 205784 234880
rect 206572 228002 206600 239700
rect 206664 239686 206862 239714
rect 206560 227996 206612 228002
rect 206560 227938 206612 227944
rect 206664 225865 206692 239686
rect 207216 236230 207244 239700
rect 207584 237017 207612 239700
rect 207570 237008 207626 237017
rect 207570 236943 207626 236952
rect 207204 236224 207256 236230
rect 207204 236166 207256 236172
rect 207952 227934 207980 239700
rect 208044 239686 208334 239714
rect 208412 239686 208702 239714
rect 208780 239686 209070 239714
rect 207940 227928 207992 227934
rect 207940 227870 207992 227876
rect 206650 225856 206706 225865
rect 206650 225791 206706 225800
rect 208044 225729 208072 239686
rect 208412 237374 208440 239686
rect 208412 237346 208532 237374
rect 208124 235612 208176 235618
rect 208124 235554 208176 235560
rect 208136 235006 208164 235554
rect 208216 235476 208268 235482
rect 208216 235418 208268 235424
rect 208124 235000 208176 235006
rect 208124 234942 208176 234948
rect 208228 234734 208256 235418
rect 208400 235408 208452 235414
rect 208400 235350 208452 235356
rect 208412 235142 208440 235350
rect 208400 235136 208452 235142
rect 208400 235078 208452 235084
rect 208216 234728 208268 234734
rect 208216 234670 208268 234676
rect 208504 229786 208532 237346
rect 208412 229758 208532 229786
rect 208030 225720 208086 225729
rect 208030 225655 208086 225664
rect 207940 223236 207992 223242
rect 207940 223178 207992 223184
rect 207952 222970 207980 223178
rect 207940 222964 207992 222970
rect 207940 222906 207992 222912
rect 205180 222760 205232 222766
rect 205180 222702 205232 222708
rect 207388 222760 207440 222766
rect 207388 222702 207440 222708
rect 205824 222420 205876 222426
rect 205824 222362 205876 222368
rect 205836 217410 205864 222362
rect 206652 220992 206704 220998
rect 206652 220934 206704 220940
rect 206664 217410 206692 220934
rect 207400 217410 207428 222702
rect 208412 222698 208440 229758
rect 208492 227724 208544 227730
rect 208492 227666 208544 227672
rect 208400 222692 208452 222698
rect 208400 222634 208452 222640
rect 208032 221332 208084 221338
rect 208032 221274 208084 221280
rect 208044 221066 208072 221274
rect 208124 221128 208176 221134
rect 208176 221076 208440 221082
rect 208124 221070 208440 221076
rect 208136 221066 208440 221070
rect 208032 221060 208084 221066
rect 208136 221060 208452 221066
rect 208136 221054 208400 221060
rect 208032 221002 208084 221008
rect 208400 221002 208452 221008
rect 208124 220992 208176 220998
rect 208176 220940 208348 220946
rect 208124 220934 208348 220940
rect 208136 220930 208348 220934
rect 208136 220924 208360 220930
rect 208136 220918 208308 220924
rect 208308 220866 208360 220872
rect 208504 218054 208532 227666
rect 208780 222494 208808 239686
rect 209424 228070 209452 239700
rect 209516 239686 209714 239714
rect 209412 228064 209464 228070
rect 209412 228006 209464 228012
rect 209516 225214 209544 239686
rect 210068 237153 210096 239700
rect 210054 237144 210110 237153
rect 210054 237079 210110 237088
rect 209688 236496 209740 236502
rect 209688 236438 209740 236444
rect 209504 225208 209556 225214
rect 209504 225150 209556 225156
rect 209136 222624 209188 222630
rect 209136 222566 209188 222572
rect 208768 222488 208820 222494
rect 208768 222430 208820 222436
rect 208320 218026 208532 218054
rect 208320 217410 208348 218026
rect 209148 217410 209176 222566
rect 209700 217410 209728 236438
rect 210436 234802 210464 239700
rect 210424 234796 210476 234802
rect 210424 234738 210476 234744
rect 210804 228138 210832 239700
rect 210896 239686 211186 239714
rect 211264 239686 211554 239714
rect 211632 239686 211922 239714
rect 212000 239686 212290 239714
rect 212566 239686 212856 239714
rect 210792 228132 210844 228138
rect 210792 228074 210844 228080
rect 210896 226001 210924 239686
rect 210976 236224 211028 236230
rect 210976 236166 211028 236172
rect 210882 225992 210938 226001
rect 210882 225927 210938 225936
rect 210988 218054 211016 236166
rect 211264 223009 211292 239686
rect 211250 223000 211306 223009
rect 211250 222935 211306 222944
rect 211632 222834 211660 239686
rect 211712 227860 211764 227866
rect 211712 227802 211764 227808
rect 211620 222828 211672 222834
rect 211620 222770 211672 222776
rect 210804 218026 211016 218054
rect 210804 217410 210832 218026
rect 211724 217410 211752 227802
rect 212000 225350 212028 239686
rect 212540 234796 212592 234802
rect 212540 234738 212592 234744
rect 211988 225344 212040 225350
rect 211988 225286 212040 225292
rect 212552 222970 212580 234738
rect 212828 226137 212856 239686
rect 212920 234938 212948 239700
rect 213288 236366 213316 239700
rect 213380 239686 213670 239714
rect 213748 239686 214038 239714
rect 214116 239686 214406 239714
rect 214484 239686 214774 239714
rect 214852 239686 215142 239714
rect 215418 239686 215708 239714
rect 213276 236360 213328 236366
rect 213276 236302 213328 236308
rect 212908 234932 212960 234938
rect 212908 234874 212960 234880
rect 212814 226128 212870 226137
rect 212814 226063 212870 226072
rect 213380 225282 213408 239686
rect 213748 225486 213776 239686
rect 213736 225480 213788 225486
rect 213736 225422 213788 225428
rect 213368 225276 213420 225282
rect 213368 225218 213420 225224
rect 212540 222964 212592 222970
rect 212540 222906 212592 222912
rect 214116 222902 214144 239686
rect 214484 223145 214512 239686
rect 214852 225418 214880 239686
rect 215300 234660 215352 234666
rect 215300 234602 215352 234608
rect 215024 227928 215076 227934
rect 215024 227870 215076 227876
rect 214840 225412 214892 225418
rect 214840 225354 214892 225360
rect 214470 223136 214526 223145
rect 214470 223071 214526 223080
rect 214104 222896 214156 222902
rect 214104 222838 214156 222844
rect 214196 222896 214248 222902
rect 214196 222838 214248 222844
rect 212356 222556 212408 222562
rect 212356 222498 212408 222504
rect 212368 217410 212396 222498
rect 213368 222488 213420 222494
rect 213368 222430 213420 222436
rect 213380 217410 213408 222430
rect 214208 217410 214236 222838
rect 215036 217410 215064 227870
rect 215312 223242 215340 234602
rect 215680 225554 215708 239686
rect 215772 236434 215800 239700
rect 216140 236978 216168 239700
rect 216232 239686 216522 239714
rect 216600 239686 216890 239714
rect 216128 236972 216180 236978
rect 216128 236914 216180 236920
rect 215760 236428 215812 236434
rect 215760 236370 215812 236376
rect 216232 225758 216260 239686
rect 216220 225752 216272 225758
rect 216220 225694 216272 225700
rect 216600 225622 216628 239686
rect 216680 236360 216732 236366
rect 216680 236302 216732 236308
rect 216588 225616 216640 225622
rect 216588 225558 216640 225564
rect 215668 225548 215720 225554
rect 215668 225490 215720 225496
rect 215300 223236 215352 223242
rect 215300 223178 215352 223184
rect 215852 222828 215904 222834
rect 215852 222770 215904 222776
rect 215864 217410 215892 222770
rect 216692 217410 216720 236302
rect 217244 234802 217272 239700
rect 217336 239686 217626 239714
rect 217704 239686 217994 239714
rect 217232 234796 217284 234802
rect 217232 234738 217284 234744
rect 217336 223281 217364 239686
rect 217704 237374 217732 239686
rect 217612 237346 217732 237374
rect 217612 225962 217640 237346
rect 217690 235920 217746 235929
rect 217690 235855 217746 235864
rect 217600 225956 217652 225962
rect 217600 225898 217652 225904
rect 217322 223272 217378 223281
rect 217322 223207 217378 223216
rect 217704 217410 217732 235855
rect 218256 225690 218284 239700
rect 218624 236774 218652 239700
rect 218992 237250 219020 239700
rect 219084 239686 219374 239714
rect 218980 237244 219032 237250
rect 218980 237186 219032 237192
rect 218612 236768 218664 236774
rect 218612 236710 218664 236716
rect 218428 233028 218480 233034
rect 218428 232970 218480 232976
rect 218336 227996 218388 228002
rect 218336 227938 218388 227944
rect 218244 225684 218296 225690
rect 218244 225626 218296 225632
rect 218348 217410 218376 227938
rect 218440 223106 218468 232970
rect 219084 225894 219112 239686
rect 219728 228206 219756 239700
rect 220096 234666 220124 239700
rect 220188 239686 220478 239714
rect 220846 239686 221044 239714
rect 221122 239686 221228 239714
rect 220084 234660 220136 234666
rect 220084 234602 220136 234608
rect 220188 233034 220216 239686
rect 220728 236768 220780 236774
rect 220728 236710 220780 236716
rect 220636 236428 220688 236434
rect 220636 236370 220688 236376
rect 220176 233028 220228 233034
rect 220176 232970 220228 232976
rect 219716 228200 219768 228206
rect 219716 228142 219768 228148
rect 219072 225888 219124 225894
rect 219072 225830 219124 225836
rect 220084 223168 220136 223174
rect 220084 223110 220136 223116
rect 218428 223100 218480 223106
rect 218428 223042 218480 223048
rect 219256 220924 219308 220930
rect 219256 220866 219308 220872
rect 219268 217410 219296 220866
rect 220096 217410 220124 223110
rect 220648 220930 220676 236370
rect 220636 220924 220688 220930
rect 220636 220866 220688 220872
rect 220740 217410 220768 236710
rect 221016 225826 221044 239686
rect 221096 233028 221148 233034
rect 221096 232970 221148 232976
rect 221108 226030 221136 232970
rect 221200 228274 221228 239686
rect 221292 239686 221490 239714
rect 221568 239686 221858 239714
rect 221936 239686 222226 239714
rect 221188 228268 221240 228274
rect 221188 228210 221240 228216
rect 221096 226024 221148 226030
rect 221096 225966 221148 225972
rect 221004 225820 221056 225826
rect 221004 225762 221056 225768
rect 221292 223242 221320 239686
rect 221568 223417 221596 239686
rect 221936 233034 221964 239686
rect 221924 233028 221976 233034
rect 221924 232970 221976 232976
rect 222580 228342 222608 239700
rect 222948 235618 222976 239700
rect 222936 235612 222988 235618
rect 222936 235554 222988 235560
rect 223316 235550 223344 239700
rect 223698 239686 223896 239714
rect 223488 236972 223540 236978
rect 223488 236914 223540 236920
rect 223304 235544 223356 235550
rect 223304 235486 223356 235492
rect 222568 228336 222620 228342
rect 222568 228278 222620 228284
rect 221740 228064 221792 228070
rect 221740 228006 221792 228012
rect 221554 223408 221610 223417
rect 221554 223343 221610 223352
rect 221280 223236 221332 223242
rect 221280 223178 221332 223184
rect 220820 222488 220872 222494
rect 220820 222430 220872 222436
rect 220832 220930 220860 222430
rect 220820 220924 220872 220930
rect 220820 220866 220872 220872
rect 221752 217410 221780 228006
rect 222568 222692 222620 222698
rect 222568 222634 222620 222640
rect 222580 217410 222608 222634
rect 223500 217410 223528 236914
rect 223764 233028 223816 233034
rect 223764 232970 223816 232976
rect 223776 226166 223804 232970
rect 223764 226160 223816 226166
rect 223764 226102 223816 226108
rect 223868 226098 223896 239686
rect 223960 228410 223988 239700
rect 224144 239686 224342 239714
rect 224144 238610 224172 239686
rect 224132 238604 224184 238610
rect 224132 238546 224184 238552
rect 224132 238400 224184 238406
rect 224132 238342 224184 238348
rect 224040 235612 224092 235618
rect 224040 235554 224092 235560
rect 223948 228404 224000 228410
rect 223948 228346 224000 228352
rect 223856 226092 223908 226098
rect 223856 226034 223908 226040
rect 224052 223310 224080 235554
rect 224144 223378 224172 238342
rect 224696 235618 224724 239700
rect 224788 239686 225078 239714
rect 224684 235612 224736 235618
rect 224684 235554 224736 235560
rect 224788 233034 224816 239686
rect 224776 233028 224828 233034
rect 224776 232970 224828 232976
rect 225432 228478 225460 239700
rect 225800 235006 225828 239700
rect 226168 236910 226196 239700
rect 226156 236904 226208 236910
rect 226156 236846 226208 236852
rect 226248 236904 226300 236910
rect 226248 236846 226300 236852
rect 226260 236586 226288 236846
rect 226168 236558 226288 236586
rect 226168 236502 226196 236558
rect 226156 236496 226208 236502
rect 226156 236438 226208 236444
rect 226246 236056 226302 236065
rect 226246 235991 226302 236000
rect 225788 235000 225840 235006
rect 225788 234942 225840 234948
rect 225420 228472 225472 228478
rect 225420 228414 225472 228420
rect 226260 226334 226288 235991
rect 226076 226306 226288 226334
rect 225144 225208 225196 225214
rect 225144 225150 225196 225156
rect 224132 223372 224184 223378
rect 224132 223314 224184 223320
rect 224040 223304 224092 223310
rect 224040 223246 224092 223252
rect 224316 223032 224368 223038
rect 224316 222974 224368 222980
rect 224328 217410 224356 222974
rect 225156 217410 225184 225150
rect 226076 217410 226104 226306
rect 226536 226234 226564 239700
rect 226720 239686 226826 239714
rect 226904 239686 227194 239714
rect 227272 239686 227562 239714
rect 227640 239686 227930 239714
rect 226616 233096 226668 233102
rect 226616 233038 226668 233044
rect 226628 226302 226656 233038
rect 226720 228546 226748 239686
rect 226800 233028 226852 233034
rect 226800 232970 226852 232976
rect 226708 228540 226760 228546
rect 226708 228482 226760 228488
rect 226616 226296 226668 226302
rect 226616 226238 226668 226244
rect 226524 226228 226576 226234
rect 226524 226170 226576 226176
rect 226812 223446 226840 232970
rect 226800 223440 226852 223446
rect 226800 223382 226852 223388
rect 226616 223100 226668 223106
rect 226616 223042 226668 223048
rect 226628 221270 226656 223042
rect 226616 221264 226668 221270
rect 226616 221206 226668 221212
rect 226708 221264 226760 221270
rect 226708 221206 226760 221212
rect 226720 221134 226748 221206
rect 226708 221128 226760 221134
rect 226708 221070 226760 221076
rect 226800 221128 226852 221134
rect 226800 221070 226852 221076
rect 226812 217410 226840 221070
rect 226904 220862 226932 239686
rect 227272 233034 227300 239686
rect 227640 233102 227668 239686
rect 227628 233096 227680 233102
rect 227628 233038 227680 233044
rect 227260 233028 227312 233034
rect 227260 232970 227312 232976
rect 228284 228614 228312 239700
rect 228652 234734 228680 239700
rect 229020 237046 229048 239700
rect 229008 237040 229060 237046
rect 229008 236982 229060 236988
rect 229006 236192 229062 236201
rect 229006 236127 229062 236136
rect 228640 234728 228692 234734
rect 228640 234670 228692 234676
rect 228272 228608 228324 228614
rect 228272 228550 228324 228556
rect 228456 225344 228508 225350
rect 228456 225286 228508 225292
rect 227536 223440 227588 223446
rect 227536 223382 227588 223388
rect 227548 221406 227576 223382
rect 227536 221400 227588 221406
rect 227536 221342 227588 221348
rect 227628 221400 227680 221406
rect 227628 221342 227680 221348
rect 226892 220856 226944 220862
rect 226892 220798 226944 220804
rect 227640 217410 227668 221342
rect 228468 217410 228496 225286
rect 229020 221406 229048 236127
rect 229284 233096 229336 233102
rect 229284 233038 229336 233044
rect 229192 233028 229244 233034
rect 229192 232970 229244 232976
rect 229204 223582 229232 232970
rect 229296 224806 229324 233038
rect 229388 224874 229416 239700
rect 229664 228682 229692 239700
rect 229756 239686 230046 239714
rect 230124 239686 230414 239714
rect 230492 239686 230782 239714
rect 229652 228676 229704 228682
rect 229652 228618 229704 228624
rect 229376 224868 229428 224874
rect 229376 224810 229428 224816
rect 229284 224800 229336 224806
rect 229284 224742 229336 224748
rect 229192 223576 229244 223582
rect 229192 223518 229244 223524
rect 229756 223514 229784 239686
rect 230124 233034 230152 239686
rect 230492 233102 230520 239686
rect 230480 233096 230532 233102
rect 230480 233038 230532 233044
rect 230112 233028 230164 233034
rect 230112 232970 230164 232976
rect 231136 228750 231164 239700
rect 231504 235414 231532 239700
rect 231872 236638 231900 239700
rect 232148 239686 232254 239714
rect 231860 236632 231912 236638
rect 231860 236574 231912 236580
rect 231492 235408 231544 235414
rect 231492 235350 231544 235356
rect 232044 233096 232096 233102
rect 232044 233038 232096 233044
rect 231124 228744 231176 228750
rect 231124 228686 231176 228692
rect 231768 225276 231820 225282
rect 231768 225218 231820 225224
rect 229744 223508 229796 223514
rect 229744 223450 229796 223456
rect 230940 223508 230992 223514
rect 230940 223450 230992 223456
rect 229284 223372 229336 223378
rect 229284 223314 229336 223320
rect 229296 221542 229324 223314
rect 230952 223106 230980 223450
rect 230940 223100 230992 223106
rect 230940 223042 230992 223048
rect 231032 223100 231084 223106
rect 231032 223042 231084 223048
rect 229376 222964 229428 222970
rect 229376 222906 229428 222912
rect 229284 221536 229336 221542
rect 229284 221478 229336 221484
rect 229008 221400 229060 221406
rect 229008 221342 229060 221348
rect 229388 217410 229416 222906
rect 229560 221536 229612 221542
rect 229560 221478 229612 221484
rect 229572 220930 229600 221478
rect 230204 221060 230256 221066
rect 230204 221002 230256 221008
rect 229560 220924 229612 220930
rect 229560 220866 229612 220872
rect 230216 217410 230244 221002
rect 231044 217410 231072 223042
rect 231780 217410 231808 225218
rect 232056 224602 232084 233038
rect 232148 224738 232176 239686
rect 232320 233028 232372 233034
rect 232320 232970 232372 232976
rect 232136 224732 232188 224738
rect 232136 224674 232188 224680
rect 232044 224596 232096 224602
rect 232044 224538 232096 224544
rect 232332 222154 232360 232970
rect 232516 228818 232544 239700
rect 232608 239686 232898 239714
rect 232976 239686 233266 239714
rect 233344 239686 233634 239714
rect 232504 228812 232556 228818
rect 232504 228754 232556 228760
rect 232320 222148 232372 222154
rect 232320 222090 232372 222096
rect 232608 222086 232636 239686
rect 232976 233034 233004 239686
rect 233148 234932 233200 234938
rect 233148 234874 233200 234880
rect 232964 233028 233016 233034
rect 232964 232970 233016 232976
rect 232596 222080 232648 222086
rect 232596 222022 232648 222028
rect 232228 221808 232280 221814
rect 232504 221808 232556 221814
rect 232280 221768 232504 221796
rect 232228 221750 232280 221756
rect 232504 221750 232556 221756
rect 232228 221672 232280 221678
rect 232412 221672 232464 221678
rect 232280 221620 232412 221626
rect 232228 221614 232464 221620
rect 232136 221604 232188 221610
rect 232240 221598 232452 221614
rect 232136 221546 232188 221552
rect 232148 221406 232176 221546
rect 232136 221400 232188 221406
rect 232136 221342 232188 221348
rect 233160 220998 233188 234874
rect 233240 234864 233292 234870
rect 233240 234806 233292 234812
rect 233252 221270 233280 234806
rect 233344 233102 233372 239686
rect 233424 235408 233476 235414
rect 233424 235350 233476 235356
rect 233332 233096 233384 233102
rect 233332 233038 233384 233044
rect 233240 221264 233292 221270
rect 233240 221206 233292 221212
rect 233148 220992 233200 220998
rect 233148 220934 233200 220940
rect 233436 220930 233464 235350
rect 233988 228886 234016 239700
rect 234356 237114 234384 239700
rect 234344 237108 234396 237114
rect 234344 237050 234396 237056
rect 234724 236842 234752 239700
rect 234908 239686 235106 239714
rect 234712 236836 234764 236842
rect 234712 236778 234764 236784
rect 234526 236328 234582 236337
rect 234526 236263 234582 236272
rect 233976 228880 234028 228886
rect 233976 228822 234028 228828
rect 233516 222080 233568 222086
rect 233516 222022 233568 222028
rect 233528 221338 233556 222022
rect 234344 221876 234396 221882
rect 234344 221818 234396 221824
rect 233516 221332 233568 221338
rect 233516 221274 233568 221280
rect 233424 220924 233476 220930
rect 233424 220866 233476 220872
rect 233516 220924 233568 220930
rect 233516 220866 233568 220872
rect 232688 220856 232740 220862
rect 232688 220798 232740 220804
rect 232700 217410 232728 220798
rect 233528 217410 233556 220866
rect 234356 217410 234384 221818
rect 234540 220862 234568 236263
rect 234804 233096 234856 233102
rect 234804 233038 234856 233044
rect 234816 224466 234844 233038
rect 234908 224670 234936 239686
rect 235172 233028 235224 233034
rect 235172 232970 235224 232976
rect 234896 224664 234948 224670
rect 234896 224606 234948 224612
rect 234804 224460 234856 224466
rect 234804 224402 234856 224408
rect 235184 221950 235212 232970
rect 235368 228954 235396 239700
rect 235460 239686 235750 239714
rect 235828 239686 236118 239714
rect 236196 239686 236486 239714
rect 235356 228948 235408 228954
rect 235356 228890 235408 228896
rect 235460 222018 235488 239686
rect 235828 233034 235856 239686
rect 236092 235476 236144 235482
rect 236092 235418 236144 235424
rect 236000 235136 236052 235142
rect 236000 235078 236052 235084
rect 235816 233028 235868 233034
rect 235816 232970 235868 232976
rect 236012 230738 236040 235078
rect 235920 230710 236040 230738
rect 235920 223174 235948 230710
rect 236104 226334 236132 235418
rect 236196 233102 236224 239686
rect 236276 235204 236328 235210
rect 236276 235146 236328 235152
rect 236288 234938 236316 235146
rect 236276 234932 236328 234938
rect 236276 234874 236328 234880
rect 236184 233096 236236 233102
rect 236184 233038 236236 233044
rect 236840 229022 236868 239700
rect 237208 237386 237236 239700
rect 237196 237380 237248 237386
rect 237196 237322 237248 237328
rect 237576 237182 237604 239700
rect 237668 239686 237958 239714
rect 237564 237176 237616 237182
rect 237564 237118 237616 237124
rect 237288 236632 237340 236638
rect 237288 236574 237340 236580
rect 236828 229016 236880 229022
rect 236828 228958 236880 228964
rect 236012 226306 236132 226334
rect 235908 223168 235960 223174
rect 235908 223110 235960 223116
rect 235816 222828 235868 222834
rect 235816 222770 235868 222776
rect 235828 222630 235856 222770
rect 235816 222624 235868 222630
rect 235816 222566 235868 222572
rect 235448 222012 235500 222018
rect 235448 221954 235500 221960
rect 235172 221944 235224 221950
rect 235172 221886 235224 221892
rect 236012 221542 236040 226306
rect 236092 222964 236144 222970
rect 236092 222906 236144 222912
rect 236000 221536 236052 221542
rect 236000 221478 236052 221484
rect 235264 221400 235316 221406
rect 235264 221342 235316 221348
rect 234528 220856 234580 220862
rect 234528 220798 234580 220804
rect 235276 217410 235304 221342
rect 236104 217410 236132 222906
rect 236920 221536 236972 221542
rect 236920 221478 236972 221484
rect 236932 217410 236960 221478
rect 237300 221406 237328 236574
rect 237668 233050 237696 239686
rect 237576 233022 237696 233050
rect 237748 233028 237800 233034
rect 237576 224534 237604 233022
rect 237748 232970 237800 232976
rect 237656 232960 237708 232966
rect 237656 232902 237708 232908
rect 237564 224528 237616 224534
rect 237564 224470 237616 224476
rect 237668 224398 237696 232902
rect 237656 224392 237708 224398
rect 237656 224334 237708 224340
rect 237760 223394 237788 232970
rect 238220 230586 238248 239700
rect 238312 239686 238602 239714
rect 238680 239686 238970 239714
rect 239048 239686 239338 239714
rect 238208 230580 238260 230586
rect 238208 230522 238260 230528
rect 237668 223366 237788 223394
rect 237668 221814 237696 223366
rect 237748 223236 237800 223242
rect 237748 223178 237800 223184
rect 237656 221808 237708 221814
rect 237656 221750 237708 221756
rect 237288 221400 237340 221406
rect 237288 221342 237340 221348
rect 237760 217410 237788 223178
rect 238312 221746 238340 239686
rect 238680 233034 238708 239686
rect 238944 237380 238996 237386
rect 238944 237322 238996 237328
rect 238852 237176 238904 237182
rect 238852 237118 238904 237124
rect 238758 236600 238814 236609
rect 238758 236535 238814 236544
rect 238668 233028 238720 233034
rect 238668 232970 238720 232976
rect 238772 231418 238800 236535
rect 238680 231390 238800 231418
rect 238300 221740 238352 221746
rect 238300 221682 238352 221688
rect 238576 221264 238628 221270
rect 238576 221206 238628 221212
rect 238588 217410 238616 221206
rect 238680 220930 238708 231390
rect 238864 231282 238892 237118
rect 238772 231254 238892 231282
rect 238772 221134 238800 231254
rect 238760 221128 238812 221134
rect 238760 221070 238812 221076
rect 238956 221066 238984 237322
rect 239048 232966 239076 239686
rect 239036 232960 239088 232966
rect 239036 232902 239088 232908
rect 239692 230722 239720 239700
rect 239784 239686 240074 239714
rect 239784 235890 239812 239686
rect 240428 237318 240456 239700
rect 240612 239686 240810 239714
rect 240416 237312 240468 237318
rect 240416 237254 240468 237260
rect 239956 236564 240008 236570
rect 239956 236506 240008 236512
rect 239772 235884 239824 235890
rect 239772 235826 239824 235832
rect 239680 230716 239732 230722
rect 239680 230658 239732 230664
rect 239404 221332 239456 221338
rect 239404 221274 239456 221280
rect 238944 221060 238996 221066
rect 238944 221002 238996 221008
rect 238668 220924 238720 220930
rect 238668 220866 238720 220872
rect 239416 217410 239444 221274
rect 239968 221270 239996 236506
rect 240046 236464 240102 236473
rect 240046 236399 240102 236408
rect 240060 221338 240088 236399
rect 240324 233096 240376 233102
rect 240324 233038 240376 233044
rect 240336 224262 240364 233038
rect 240508 233028 240560 233034
rect 240508 232970 240560 232976
rect 240324 224256 240376 224262
rect 240324 224198 240376 224204
rect 240520 221678 240548 232970
rect 240612 224330 240640 239686
rect 241072 230654 241100 239700
rect 241164 239686 241454 239714
rect 241532 239686 241822 239714
rect 241900 239686 242190 239714
rect 241164 235958 241192 239686
rect 241428 236836 241480 236842
rect 241428 236778 241480 236784
rect 241152 235952 241204 235958
rect 241152 235894 241204 235900
rect 241060 230648 241112 230654
rect 241060 230590 241112 230596
rect 240600 224324 240652 224330
rect 240600 224266 240652 224272
rect 241152 223304 241204 223310
rect 241152 223246 241204 223252
rect 240508 221672 240560 221678
rect 240508 221614 240560 221620
rect 240048 221332 240100 221338
rect 240048 221274 240100 221280
rect 239956 221264 240008 221270
rect 239956 221206 240008 221212
rect 240048 221128 240100 221134
rect 240048 221070 240100 221076
rect 240060 217410 240088 221070
rect 241164 217410 241192 223246
rect 241440 221134 241468 236778
rect 241532 233034 241560 239686
rect 241612 237312 241664 237318
rect 241612 237254 241664 237260
rect 241520 233028 241572 233034
rect 241520 232970 241572 232976
rect 241624 231962 241652 237254
rect 241796 234660 241848 234666
rect 241796 234602 241848 234608
rect 241532 231934 241652 231962
rect 241532 221542 241560 231934
rect 241808 231690 241836 234602
rect 241900 233102 241928 239686
rect 241888 233096 241940 233102
rect 241888 233038 241940 233044
rect 241624 231662 241836 231690
rect 241624 221610 241652 231662
rect 242544 230858 242572 239700
rect 242808 237108 242860 237114
rect 242808 237050 242860 237056
rect 242532 230852 242584 230858
rect 242532 230794 242584 230800
rect 242716 223168 242768 223174
rect 242716 223110 242768 223116
rect 241612 221604 241664 221610
rect 241612 221546 241664 221552
rect 241520 221536 241572 221542
rect 241520 221478 241572 221484
rect 241980 221332 242032 221338
rect 241980 221274 242032 221280
rect 241428 221128 241480 221134
rect 241428 221070 241480 221076
rect 241992 217410 242020 221274
rect 242728 217410 242756 223110
rect 242820 221338 242848 237050
rect 242912 234666 242940 239700
rect 243280 235754 243308 239700
rect 243464 239686 243662 239714
rect 243268 235748 243320 235754
rect 243268 235690 243320 235696
rect 242900 234660 242952 234666
rect 242900 234602 242952 234608
rect 243084 233096 243136 233102
rect 243084 233038 243136 233044
rect 243096 224126 243124 233038
rect 243268 233028 243320 233034
rect 243268 232970 243320 232976
rect 243084 224120 243136 224126
rect 243084 224062 243136 224068
rect 243280 221406 243308 232970
rect 243464 224194 243492 239686
rect 243924 230790 243952 239700
rect 244292 235822 244320 239700
rect 244384 239686 244674 239714
rect 244752 239686 245042 239714
rect 244280 235816 244332 235822
rect 244280 235758 244332 235764
rect 244280 235544 244332 235550
rect 244280 235486 244332 235492
rect 244188 235408 244240 235414
rect 244188 235350 244240 235356
rect 243912 230784 243964 230790
rect 243912 230726 243964 230732
rect 243452 224188 243504 224194
rect 243452 224130 243504 224136
rect 244200 223378 244228 235350
rect 244292 223514 244320 235486
rect 244384 233034 244412 239686
rect 244464 234728 244516 234734
rect 244464 234670 244516 234676
rect 244372 233028 244424 233034
rect 244372 232970 244424 232976
rect 244476 223514 244504 234670
rect 244752 233102 244780 239686
rect 244740 233096 244792 233102
rect 244740 233038 244792 233044
rect 245396 230994 245424 239700
rect 245476 237040 245528 237046
rect 245476 236982 245528 236988
rect 245384 230988 245436 230994
rect 245384 230930 245436 230936
rect 245488 226334 245516 236982
rect 245568 235952 245620 235958
rect 245568 235894 245620 235900
rect 245396 226306 245516 226334
rect 244280 223508 244332 223514
rect 244280 223450 244332 223456
rect 244464 223508 244516 223514
rect 244464 223450 244516 223456
rect 244188 223372 244240 223378
rect 244188 223314 244240 223320
rect 244464 223372 244516 223378
rect 244464 223314 244516 223320
rect 243268 221400 243320 221406
rect 243268 221342 243320 221348
rect 242808 221332 242860 221338
rect 242808 221274 242860 221280
rect 243636 220856 243688 220862
rect 243636 220798 243688 220804
rect 243648 217410 243676 220798
rect 244476 217410 244504 223314
rect 245396 217410 245424 226306
rect 245580 220862 245608 235894
rect 245764 235414 245792 239700
rect 246132 235686 246160 239700
rect 246224 239686 246514 239714
rect 246120 235680 246172 235686
rect 246120 235622 246172 235628
rect 245752 235408 245804 235414
rect 245752 235350 245804 235356
rect 245844 233096 245896 233102
rect 245844 233038 245896 233044
rect 245856 223990 245884 233038
rect 246028 233028 246080 233034
rect 246028 232970 246080 232976
rect 245844 223984 245896 223990
rect 245844 223926 245896 223932
rect 246040 221474 246068 232970
rect 246224 224058 246252 239686
rect 246776 230926 246804 239700
rect 247144 235618 247172 239700
rect 247236 239686 247526 239714
rect 247604 239686 247894 239714
rect 247132 235612 247184 235618
rect 247132 235554 247184 235560
rect 246948 235136 247000 235142
rect 246948 235078 247000 235084
rect 247132 235136 247184 235142
rect 247132 235078 247184 235084
rect 246960 234802 246988 235078
rect 247040 234864 247092 234870
rect 247040 234806 247092 234812
rect 246948 234796 247000 234802
rect 246948 234738 247000 234744
rect 246948 234660 247000 234666
rect 246948 234602 247000 234608
rect 246764 230920 246816 230926
rect 246764 230862 246816 230868
rect 246212 224052 246264 224058
rect 246212 223994 246264 224000
rect 246960 222290 246988 234602
rect 246948 222284 247000 222290
rect 246948 222226 247000 222232
rect 246120 221536 246172 221542
rect 247052 221490 247080 234806
rect 247144 222766 247172 235078
rect 247236 233034 247264 239686
rect 247316 235748 247368 235754
rect 247316 235690 247368 235696
rect 247224 233028 247276 233034
rect 247224 232970 247276 232976
rect 247328 222834 247356 235690
rect 247604 233102 247632 239686
rect 247592 233096 247644 233102
rect 247592 233038 247644 233044
rect 248248 231062 248276 239700
rect 248328 235952 248380 235958
rect 248328 235894 248380 235900
rect 248236 231056 248288 231062
rect 248236 230998 248288 231004
rect 247316 222828 247368 222834
rect 247316 222770 247368 222776
rect 247132 222760 247184 222766
rect 247132 222702 247184 222708
rect 246120 221478 246172 221484
rect 246028 221468 246080 221474
rect 246028 221410 246080 221416
rect 245568 220856 245620 220862
rect 245568 220798 245620 220804
rect 246132 217410 246160 221478
rect 246960 221462 247080 221490
rect 246960 221202 246988 221462
rect 248340 221406 248368 235894
rect 248616 234734 248644 239700
rect 248984 235074 249012 239700
rect 249076 239686 249366 239714
rect 248972 235068 249024 235074
rect 248972 235010 249024 235016
rect 248604 234728 248656 234734
rect 248604 234670 248656 234676
rect 248604 233028 248656 233034
rect 248604 232970 248656 232976
rect 248616 224942 248644 232970
rect 248788 228132 248840 228138
rect 248788 228074 248840 228080
rect 248604 224936 248656 224942
rect 248604 224878 248656 224884
rect 248800 222086 248828 228074
rect 249076 223922 249104 239686
rect 249628 234938 249656 239700
rect 249890 237008 249946 237017
rect 249890 236943 249946 236952
rect 249706 236736 249762 236745
rect 249706 236671 249762 236680
rect 249616 234932 249668 234938
rect 249616 234874 249668 234880
rect 249064 223916 249116 223922
rect 249064 223858 249116 223864
rect 248788 222080 248840 222086
rect 248788 222022 248840 222028
rect 249720 221882 249748 236671
rect 249904 223106 249932 236943
rect 249996 235550 250024 239700
rect 250088 239686 250378 239714
rect 250456 239686 250746 239714
rect 250824 239686 251114 239714
rect 249984 235544 250036 235550
rect 249984 235486 250036 235492
rect 250088 228138 250116 239686
rect 250166 237280 250222 237289
rect 250166 237215 250222 237224
rect 250076 228132 250128 228138
rect 250076 228074 250128 228080
rect 249892 223100 249944 223106
rect 249892 223042 249944 223048
rect 250180 223038 250208 237215
rect 250456 233034 250484 239686
rect 250824 235006 250852 239686
rect 250996 235816 251048 235822
rect 250996 235758 251048 235764
rect 250812 235000 250864 235006
rect 250812 234942 250864 234948
rect 250444 233028 250496 233034
rect 250444 232970 250496 232976
rect 250168 223032 250220 223038
rect 250168 222974 250220 222980
rect 249708 221876 249760 221882
rect 249708 221818 249760 221824
rect 249524 221468 249576 221474
rect 249524 221410 249576 221416
rect 247040 221400 247092 221406
rect 247040 221342 247092 221348
rect 248328 221400 248380 221406
rect 248328 221342 248380 221348
rect 246948 221196 247000 221202
rect 246948 221138 247000 221144
rect 247052 217410 247080 221342
rect 247868 221264 247920 221270
rect 247868 221206 247920 221212
rect 247880 217410 247908 221206
rect 248696 220856 248748 220862
rect 248696 220798 248748 220804
rect 248708 217410 248736 220798
rect 249536 217410 249564 221410
rect 251008 221338 251036 235758
rect 251088 235680 251140 235686
rect 251088 235622 251140 235628
rect 250352 221332 250404 221338
rect 250352 221274 250404 221280
rect 250996 221332 251048 221338
rect 250996 221274 251048 221280
rect 250364 217410 250392 221274
rect 250996 221128 251048 221134
rect 250996 221070 251048 221076
rect 251008 217410 251036 221070
rect 251100 220862 251128 235622
rect 251468 235278 251496 239700
rect 251836 236094 251864 239700
rect 251928 239686 252218 239714
rect 251824 236088 251876 236094
rect 251824 236030 251876 236036
rect 251456 235272 251508 235278
rect 251456 235214 251508 235220
rect 251364 233096 251416 233102
rect 251364 233038 251416 233044
rect 251376 225078 251404 233038
rect 251456 233028 251508 233034
rect 251456 232970 251508 232976
rect 251364 225072 251416 225078
rect 251364 225014 251416 225020
rect 251468 222222 251496 232970
rect 251928 225010 251956 239686
rect 252480 236706 252508 239700
rect 252558 236872 252614 236881
rect 252558 236807 252614 236816
rect 252468 236700 252520 236706
rect 252468 236642 252520 236648
rect 252572 234954 252600 236807
rect 252480 234926 252600 234954
rect 251916 225004 251968 225010
rect 251916 224946 251968 224952
rect 252480 223242 252508 234926
rect 252560 234796 252612 234802
rect 252560 234738 252612 234744
rect 252572 223310 252600 234738
rect 252848 234666 252876 239700
rect 252940 239686 253230 239714
rect 253308 239686 253598 239714
rect 252836 234660 252888 234666
rect 252836 234602 252888 234608
rect 252940 233034 252968 239686
rect 253204 236700 253256 236706
rect 253204 236642 253256 236648
rect 253216 236434 253244 236642
rect 253204 236428 253256 236434
rect 253204 236370 253256 236376
rect 253308 233102 253336 239686
rect 253756 236088 253808 236094
rect 253756 236030 253808 236036
rect 253296 233096 253348 233102
rect 253296 233038 253348 233044
rect 252928 233028 252980 233034
rect 252928 232970 252980 232976
rect 252560 223304 252612 223310
rect 252560 223246 252612 223252
rect 252468 223236 252520 223242
rect 252468 223178 252520 223184
rect 251456 222216 251508 222222
rect 251456 222158 251508 222164
rect 252928 221332 252980 221338
rect 252928 221274 252980 221280
rect 252008 221196 252060 221202
rect 252008 221138 252060 221144
rect 251088 220856 251140 220862
rect 251088 220798 251140 220804
rect 252020 217410 252048 221138
rect 252940 217410 252968 221274
rect 253768 221202 253796 236030
rect 253952 235210 253980 239700
rect 254320 236298 254348 239700
rect 254308 236292 254360 236298
rect 254308 236234 254360 236240
rect 254688 236026 254716 239700
rect 254780 239686 255070 239714
rect 254676 236020 254728 236026
rect 254676 235962 254728 235968
rect 253940 235204 253992 235210
rect 253940 235146 253992 235152
rect 253848 234728 253900 234734
rect 253848 234670 253900 234676
rect 253756 221196 253808 221202
rect 253756 221138 253808 221144
rect 253860 217410 253888 234670
rect 254216 233028 254268 233034
rect 254216 232970 254268 232976
rect 254228 222358 254256 232970
rect 254780 225146 254808 239686
rect 254860 237244 254912 237250
rect 254860 237186 254912 237192
rect 254872 236978 254900 237186
rect 254860 236972 254912 236978
rect 254860 236914 254912 236920
rect 255332 236502 255360 239700
rect 255320 236496 255372 236502
rect 255320 236438 255372 236444
rect 255412 236020 255464 236026
rect 255412 235962 255464 235968
rect 255320 235408 255372 235414
rect 255320 235350 255372 235356
rect 255228 235340 255280 235346
rect 255228 235282 255280 235288
rect 254768 225140 254820 225146
rect 254768 225082 254820 225088
rect 254216 222352 254268 222358
rect 254216 222294 254268 222300
rect 254584 221400 254636 221406
rect 254584 221342 254636 221348
rect 254596 217410 254624 221342
rect 255240 221270 255268 235282
rect 255332 223378 255360 235350
rect 255320 223372 255372 223378
rect 255320 223314 255372 223320
rect 255228 221264 255280 221270
rect 255228 221206 255280 221212
rect 255424 221134 255452 235962
rect 255504 234932 255556 234938
rect 255504 234874 255556 234880
rect 255516 223174 255544 234874
rect 255700 234870 255728 239700
rect 255792 239686 256082 239714
rect 255688 234864 255740 234870
rect 255688 234806 255740 234812
rect 255792 233034 255820 239686
rect 255780 233028 255832 233034
rect 255780 232970 255832 232976
rect 256436 227798 256464 239700
rect 256516 236292 256568 236298
rect 256516 236234 256568 236240
rect 256424 227792 256476 227798
rect 256424 227734 256476 227740
rect 255504 223168 255556 223174
rect 255504 223110 255556 223116
rect 256528 221406 256556 236234
rect 256608 235476 256660 235482
rect 256608 235418 256660 235424
rect 256516 221400 256568 221406
rect 256516 221342 256568 221348
rect 256240 221264 256292 221270
rect 256240 221206 256292 221212
rect 255412 221128 255464 221134
rect 255412 221070 255464 221076
rect 255412 220924 255464 220930
rect 255412 220866 255464 220872
rect 255424 217410 255452 220866
rect 256252 217410 256280 221206
rect 256620 220930 256648 235418
rect 256804 235278 256832 239700
rect 257172 236162 257200 239700
rect 257356 239686 257554 239714
rect 257160 236156 257212 236162
rect 257160 236098 257212 236104
rect 256792 235272 256844 235278
rect 256792 235214 256844 235220
rect 257068 233028 257120 233034
rect 257068 232970 257120 232976
rect 257080 222562 257108 232970
rect 257068 222556 257120 222562
rect 257068 222498 257120 222504
rect 257356 222426 257384 239686
rect 257908 227730 257936 239700
rect 258080 236972 258132 236978
rect 258080 236914 258132 236920
rect 257988 235068 258040 235074
rect 257988 235010 258040 235016
rect 257896 227724 257948 227730
rect 257896 227666 257948 227672
rect 257344 222420 257396 222426
rect 257344 222362 257396 222368
rect 258000 221542 258028 235010
rect 257988 221536 258040 221542
rect 257988 221478 258040 221484
rect 257068 221400 257120 221406
rect 257068 221342 257120 221348
rect 256608 220924 256660 220930
rect 256608 220866 256660 220872
rect 257080 217410 257108 221342
rect 258092 221338 258120 236914
rect 258184 236910 258212 239700
rect 258172 236904 258224 236910
rect 258172 236846 258224 236852
rect 258172 235544 258224 235550
rect 258172 235486 258224 235492
rect 258184 221474 258212 235486
rect 258552 235142 258580 239700
rect 258644 239686 258934 239714
rect 259012 239686 259302 239714
rect 258540 235136 258592 235142
rect 258540 235078 258592 235084
rect 258644 233034 258672 239686
rect 258632 233028 258684 233034
rect 258632 232970 258684 232976
rect 259012 227866 259040 239686
rect 259276 236496 259328 236502
rect 259276 236438 259328 236444
rect 259184 235204 259236 235210
rect 259184 235146 259236 235152
rect 259000 227860 259052 227866
rect 259000 227802 259052 227808
rect 258172 221468 258224 221474
rect 258172 221410 258224 221416
rect 259196 221406 259224 235146
rect 259184 221400 259236 221406
rect 259184 221342 259236 221348
rect 258080 221332 258132 221338
rect 258080 221274 258132 221280
rect 258816 221332 258868 221338
rect 258816 221274 258868 221280
rect 257896 220856 257948 220862
rect 257896 220798 257948 220804
rect 257908 217410 257936 220798
rect 258828 217410 258856 221274
rect 259288 220862 259316 236438
rect 259368 236156 259420 236162
rect 259368 236098 259420 236104
rect 259380 221338 259408 236098
rect 259656 235618 259684 239700
rect 260024 236230 260052 239700
rect 260116 239686 260406 239714
rect 260484 239686 260774 239714
rect 260012 236224 260064 236230
rect 260012 236166 260064 236172
rect 259644 235612 259696 235618
rect 259644 235554 259696 235560
rect 259828 233028 259880 233034
rect 259828 232970 259880 232976
rect 259840 222630 259868 232970
rect 259828 222624 259880 222630
rect 259828 222566 259880 222572
rect 260116 222494 260144 239686
rect 260484 227934 260512 239686
rect 261036 236434 261064 239700
rect 261024 236428 261076 236434
rect 261024 236370 261076 236376
rect 260840 236360 260892 236366
rect 260840 236302 260892 236308
rect 260748 236224 260800 236230
rect 260748 236166 260800 236172
rect 260472 227928 260524 227934
rect 260472 227870 260524 227876
rect 260104 222488 260156 222494
rect 260104 222430 260156 222436
rect 259368 221332 259420 221338
rect 259368 221274 259420 221280
rect 260760 221202 260788 236166
rect 260852 221270 260880 236302
rect 261404 235754 261432 239700
rect 261496 239686 261786 239714
rect 261864 239686 262154 239714
rect 261392 235748 261444 235754
rect 261392 235690 261444 235696
rect 261496 233034 261524 239686
rect 261484 233028 261536 233034
rect 261484 232970 261536 232976
rect 261864 228002 261892 239686
rect 261944 235612 261996 235618
rect 261944 235554 261996 235560
rect 261852 227996 261904 228002
rect 261852 227938 261904 227944
rect 260840 221264 260892 221270
rect 260840 221206 260892 221212
rect 259368 221196 259420 221202
rect 259368 221138 259420 221144
rect 260748 221196 260800 221202
rect 260748 221138 260800 221144
rect 259276 220856 259328 220862
rect 259276 220798 259328 220804
rect 259380 217410 259408 221138
rect 261956 221066 261984 235554
rect 262036 235272 262088 235278
rect 262036 235214 262088 235220
rect 260472 221060 260524 221066
rect 260472 221002 260524 221008
rect 261944 221060 261996 221066
rect 261944 221002 261996 221008
rect 260484 217410 260512 221002
rect 262048 220930 262076 235214
rect 262128 235136 262180 235142
rect 262128 235078 262180 235084
rect 261300 220924 261352 220930
rect 261300 220866 261352 220872
rect 262036 220924 262088 220930
rect 262036 220866 262088 220872
rect 261312 217410 261340 220866
rect 262140 217410 262168 235078
rect 262508 234666 262536 239700
rect 262876 235929 262904 239700
rect 263244 236706 263272 239700
rect 263232 236700 263284 236706
rect 263232 236642 263284 236648
rect 262862 235920 262918 235929
rect 262862 235855 262918 235864
rect 263508 235000 263560 235006
rect 263508 234942 263560 234948
rect 262496 234660 262548 234666
rect 262496 234602 262548 234608
rect 262588 233028 262640 233034
rect 262588 232970 262640 232976
rect 262600 222698 262628 232970
rect 263520 222902 263548 234942
rect 263612 228070 263640 239700
rect 263888 237250 263916 239700
rect 263876 237244 263928 237250
rect 263876 237186 263928 237192
rect 264256 236774 264284 239700
rect 264348 239686 264638 239714
rect 265006 239686 265296 239714
rect 264244 236768 264296 236774
rect 264244 236710 264296 236716
rect 264348 233034 264376 239686
rect 264704 236972 264756 236978
rect 264704 236914 264756 236920
rect 264336 233028 264388 233034
rect 264336 232970 264388 232976
rect 263600 228064 263652 228070
rect 263600 228006 263652 228012
rect 263508 222896 263560 222902
rect 263508 222838 263560 222844
rect 262588 222692 262640 222698
rect 262588 222634 262640 222640
rect 264716 221202 264744 236914
rect 264888 236768 264940 236774
rect 264888 236710 264940 236716
rect 264796 236428 264848 236434
rect 264796 236370 264848 236376
rect 263784 221196 263836 221202
rect 263784 221138 263836 221144
rect 264704 221196 264756 221202
rect 264704 221138 264756 221144
rect 262956 220856 263008 220862
rect 262956 220798 263008 220804
rect 262968 217410 262996 220798
rect 263796 217410 263824 221138
rect 264808 217410 264836 236370
rect 264900 220862 264928 236710
rect 265268 225214 265296 239686
rect 265360 237182 265388 239700
rect 265728 237289 265756 239700
rect 265714 237280 265770 237289
rect 265714 237215 265770 237224
rect 265348 237176 265400 237182
rect 265348 237118 265400 237124
rect 266096 236065 266124 239700
rect 266188 239686 266478 239714
rect 266082 236056 266138 236065
rect 266082 235991 266138 236000
rect 266188 225350 266216 239686
rect 266740 237386 266768 239700
rect 266728 237380 266780 237386
rect 266728 237322 266780 237328
rect 267108 236201 267136 239700
rect 267094 236192 267150 236201
rect 267094 236127 267150 236136
rect 267188 235748 267240 235754
rect 267188 235690 267240 235696
rect 267200 235278 267228 235690
rect 267188 235272 267240 235278
rect 267188 235214 267240 235220
rect 267280 235272 267332 235278
rect 267280 235214 267332 235220
rect 267292 235142 267320 235214
rect 267280 235136 267332 235142
rect 267280 235078 267332 235084
rect 267372 235136 267424 235142
rect 267372 235078 267424 235084
rect 267384 234734 267412 235078
rect 267476 235006 267504 239700
rect 267464 235000 267516 235006
rect 267464 234942 267516 234948
rect 267464 234796 267516 234802
rect 267464 234738 267516 234744
rect 267372 234728 267424 234734
rect 267372 234670 267424 234676
rect 266176 225344 266228 225350
rect 266176 225286 266228 225292
rect 265256 225208 265308 225214
rect 265256 225150 265308 225156
rect 267476 220930 267504 234738
rect 267556 234728 267608 234734
rect 267556 234670 267608 234676
rect 266360 220924 266412 220930
rect 266360 220866 266412 220872
rect 267464 220924 267516 220930
rect 267464 220866 267516 220872
rect 264888 220856 264940 220862
rect 264888 220798 264940 220804
rect 265532 220856 265584 220862
rect 265532 220798 265584 220804
rect 265544 217410 265572 220798
rect 266372 217410 266400 220866
rect 267568 217546 267596 234670
rect 267648 234660 267700 234666
rect 267648 234602 267700 234608
rect 267660 220862 267688 234602
rect 267844 225282 267872 239700
rect 268212 236609 268240 239700
rect 268580 237017 268608 239700
rect 268566 237008 268622 237017
rect 268566 236943 268622 236952
rect 268198 236600 268254 236609
rect 268198 236535 268254 236544
rect 268948 236337 268976 239700
rect 269316 236706 269344 239700
rect 269592 237318 269620 239700
rect 269580 237312 269632 237318
rect 269580 237254 269632 237260
rect 269960 236745 269988 239700
rect 270052 239686 270342 239714
rect 269946 236736 270002 236745
rect 269304 236700 269356 236706
rect 269946 236671 270002 236680
rect 269304 236642 269356 236648
rect 268934 236328 268990 236337
rect 268934 236263 268990 236272
rect 270052 233034 270080 239686
rect 270408 236632 270460 236638
rect 270408 236574 270460 236580
rect 268200 233028 268252 233034
rect 268200 232970 268252 232976
rect 270040 233028 270092 233034
rect 270040 232970 270092 232976
rect 267832 225276 267884 225282
rect 267832 225218 267884 225224
rect 268212 222970 268240 232970
rect 268200 222964 268252 222970
rect 268200 222906 268252 222912
rect 268844 221332 268896 221338
rect 268844 221274 268896 221280
rect 267648 220856 267700 220862
rect 267648 220798 267700 220804
rect 268016 220856 268068 220862
rect 268016 220798 268068 220804
rect 267292 217518 267596 217546
rect 267292 217410 267320 217518
rect 268028 217410 268056 220798
rect 268856 217410 268884 221274
rect 270420 221202 270448 236574
rect 270696 236570 270724 239700
rect 271064 236842 271092 239700
rect 271432 236881 271460 239700
rect 271418 236872 271474 236881
rect 271052 236836 271104 236842
rect 271418 236807 271474 236816
rect 271052 236778 271104 236784
rect 270684 236564 270736 236570
rect 270684 236506 270736 236512
rect 271800 236473 271828 239700
rect 272168 237114 272196 239700
rect 272156 237108 272208 237114
rect 272156 237050 272208 237056
rect 271786 236464 271842 236473
rect 271786 236399 271842 236408
rect 272444 235890 272472 239700
rect 272432 235884 272484 235890
rect 272432 235826 272484 235832
rect 272812 234870 272840 239700
rect 273180 234938 273208 239700
rect 273548 237046 273576 239700
rect 273536 237040 273588 237046
rect 273536 236982 273588 236988
rect 273916 235958 273944 239700
rect 273904 235952 273956 235958
rect 273904 235894 273956 235900
rect 274284 235414 274312 239700
rect 274272 235408 274324 235414
rect 274272 235350 274324 235356
rect 274652 235074 274680 239700
rect 275020 235686 275048 239700
rect 275296 235822 275324 239700
rect 275284 235816 275336 235822
rect 275284 235758 275336 235764
rect 275008 235680 275060 235686
rect 275008 235622 275060 235628
rect 275664 235346 275692 239700
rect 276032 235550 276060 239700
rect 276400 236094 276428 239700
rect 276388 236088 276440 236094
rect 276388 236030 276440 236036
rect 276020 235544 276072 235550
rect 276020 235486 276072 235492
rect 275652 235340 275704 235346
rect 275652 235282 275704 235288
rect 276768 235142 276796 239700
rect 277136 236026 277164 239700
rect 277504 236910 277532 239700
rect 277492 236904 277544 236910
rect 277492 236846 277544 236852
rect 277124 236020 277176 236026
rect 277124 235962 277176 235968
rect 277872 235482 277900 239700
rect 277860 235476 277912 235482
rect 277860 235418 277912 235424
rect 278148 235210 278176 239700
rect 278516 236298 278544 239700
rect 278884 236366 278912 239700
rect 278872 236360 278924 236366
rect 278872 236302 278924 236308
rect 278504 236292 278556 236298
rect 278504 236234 278556 236240
rect 279252 236162 279280 239700
rect 279240 236156 279292 236162
rect 279240 236098 279292 236104
rect 279620 235618 279648 239700
rect 279988 236502 280016 239700
rect 279976 236496 280028 236502
rect 279976 236438 280028 236444
rect 280356 236230 280384 239700
rect 280344 236224 280396 236230
rect 280344 236166 280396 236172
rect 279608 235612 279660 235618
rect 279608 235554 279660 235560
rect 280724 235278 280752 239700
rect 281000 236978 281028 239700
rect 280988 236972 281040 236978
rect 280988 236914 281040 236920
rect 281368 235754 281396 239700
rect 281736 236774 281764 239700
rect 281724 236768 281776 236774
rect 281724 236710 281776 236716
rect 281356 235748 281408 235754
rect 281356 235690 281408 235696
rect 280712 235272 280764 235278
rect 280712 235214 280764 235220
rect 278136 235204 278188 235210
rect 278136 235146 278188 235152
rect 276756 235136 276808 235142
rect 276756 235078 276808 235084
rect 274640 235068 274692 235074
rect 274640 235010 274692 235016
rect 273168 234932 273220 234938
rect 273168 234874 273220 234880
rect 272800 234864 272852 234870
rect 272800 234806 272852 234812
rect 282104 234666 282132 239700
rect 282472 234734 282500 239700
rect 282840 236434 282868 239700
rect 282828 236428 282880 236434
rect 282828 236370 282880 236376
rect 283208 234802 283236 239700
rect 283300 239686 283590 239714
rect 283668 239686 283866 239714
rect 283944 239686 284234 239714
rect 283196 234796 283248 234802
rect 283196 234738 283248 234744
rect 282460 234728 282512 234734
rect 282460 234670 282512 234676
rect 282092 234660 282144 234666
rect 282092 234602 282144 234608
rect 283300 233102 283328 239686
rect 281724 233096 281776 233102
rect 281724 233038 281776 233044
rect 283288 233096 283340 233102
rect 283288 233038 283340 233044
rect 272248 223576 272300 223582
rect 272248 223518 272300 223524
rect 271420 221468 271472 221474
rect 271420 221410 271472 221416
rect 269672 221196 269724 221202
rect 269672 221138 269724 221144
rect 270408 221196 270460 221202
rect 270408 221138 270460 221144
rect 269684 217410 269712 221138
rect 270408 221060 270460 221066
rect 270408 221002 270460 221008
rect 270420 217410 270448 221002
rect 271432 217410 271460 221410
rect 272260 217410 272288 223518
rect 273076 223508 273128 223514
rect 273076 223450 273128 223456
rect 273088 217410 273116 223450
rect 278688 223440 278740 223446
rect 278688 223382 278740 223388
rect 278136 223372 278188 223378
rect 278136 223314 278188 223320
rect 274732 222012 274784 222018
rect 274732 221954 274784 221960
rect 273904 220924 273956 220930
rect 273904 220866 273956 220872
rect 273916 217410 273944 220866
rect 274744 217410 274772 221954
rect 275560 221876 275612 221882
rect 275560 221818 275612 221824
rect 275572 217410 275600 221818
rect 276480 221604 276532 221610
rect 276480 221546 276532 221552
rect 276492 217410 276520 221546
rect 277308 221128 277360 221134
rect 277308 221070 277360 221076
rect 277320 217410 277348 221070
rect 278148 217410 278176 223314
rect 278700 217410 278728 223382
rect 281448 222760 281500 222766
rect 281448 222702 281500 222708
rect 280620 222148 280672 222154
rect 280620 222090 280672 222096
rect 279792 221672 279844 221678
rect 279792 221614 279844 221620
rect 279804 217410 279832 221614
rect 280632 217410 280660 222090
rect 281460 217410 281488 222702
rect 281736 221338 281764 233038
rect 283668 233034 283696 239686
rect 282000 233028 282052 233034
rect 282000 232970 282052 232976
rect 283656 233028 283708 233034
rect 283656 232970 283708 232976
rect 281816 232960 281868 232966
rect 281816 232902 281868 232908
rect 281724 221332 281776 221338
rect 281724 221274 281776 221280
rect 281828 220862 281856 232902
rect 282012 221066 282040 232970
rect 283944 232966 283972 239686
rect 284588 236638 284616 239700
rect 284680 239686 284970 239714
rect 285048 239686 285338 239714
rect 285416 239686 285706 239714
rect 285784 239686 286074 239714
rect 286152 239686 286442 239714
rect 286520 239686 286718 239714
rect 284576 236632 284628 236638
rect 284576 236574 284628 236580
rect 284392 233164 284444 233170
rect 284392 233106 284444 233112
rect 283932 232960 283984 232966
rect 283932 232902 283984 232908
rect 283196 222420 283248 222426
rect 283196 222362 283248 222368
rect 282000 221060 282052 221066
rect 282000 221002 282052 221008
rect 282368 221060 282420 221066
rect 282368 221002 282420 221008
rect 281816 220856 281868 220862
rect 281816 220798 281868 220804
rect 282380 217410 282408 221002
rect 283208 217410 283236 222362
rect 283932 221196 283984 221202
rect 283932 221138 283984 221144
rect 283944 217410 283972 221138
rect 284404 220930 284432 233106
rect 284680 233050 284708 239686
rect 285048 233170 285076 239686
rect 285036 233164 285088 233170
rect 285036 233106 285088 233112
rect 285416 233050 285444 239686
rect 284484 233028 284536 233034
rect 284484 232970 284536 232976
rect 284588 233022 284708 233050
rect 284772 233022 285444 233050
rect 284496 221134 284524 232970
rect 284588 223582 284616 233022
rect 284772 232948 284800 233022
rect 284680 232920 284800 232948
rect 284576 223576 284628 223582
rect 284576 223518 284628 223524
rect 284680 221474 284708 232920
rect 285784 232778 285812 239686
rect 284772 232750 285812 232778
rect 284772 223514 284800 232750
rect 286152 232694 286180 239686
rect 286520 233034 286548 239686
rect 287072 233170 287100 239700
rect 287164 239686 287454 239714
rect 287532 239686 287822 239714
rect 287900 239686 288190 239714
rect 288268 239686 288558 239714
rect 288636 239686 288926 239714
rect 289004 239686 289294 239714
rect 289372 239686 289570 239714
rect 287060 233164 287112 233170
rect 287060 233106 287112 233112
rect 287164 233050 287192 239686
rect 287244 233232 287296 233238
rect 287244 233174 287296 233180
rect 286508 233028 286560 233034
rect 286508 232970 286560 232976
rect 287072 233022 287192 233050
rect 284852 232688 284904 232694
rect 284852 232630 284904 232636
rect 286140 232688 286192 232694
rect 286140 232630 286192 232636
rect 284760 223508 284812 223514
rect 284760 223450 284812 223456
rect 284864 221882 284892 232630
rect 284852 221876 284904 221882
rect 284852 221818 284904 221824
rect 287072 221610 287100 233022
rect 287152 232892 287204 232898
rect 287152 232834 287204 232840
rect 287164 223378 287192 232834
rect 287152 223372 287204 223378
rect 287152 223314 287204 223320
rect 287256 222154 287284 233174
rect 287532 233050 287560 239686
rect 287900 233238 287928 239686
rect 287888 233232 287940 233238
rect 287888 233174 287940 233180
rect 287612 233164 287664 233170
rect 287612 233106 287664 233112
rect 287348 233022 287560 233050
rect 287348 223446 287376 233022
rect 287428 232960 287480 232966
rect 287428 232902 287480 232908
rect 287336 223440 287388 223446
rect 287336 223382 287388 223388
rect 287244 222148 287296 222154
rect 287244 222090 287296 222096
rect 287440 221678 287468 232902
rect 287624 222018 287652 233106
rect 287888 233028 287940 233034
rect 287888 232970 287940 232976
rect 287796 231532 287848 231538
rect 287796 231474 287848 231480
rect 287612 222012 287664 222018
rect 287612 221954 287664 221960
rect 287428 221672 287480 221678
rect 287428 221614 287480 221620
rect 287060 221604 287112 221610
rect 287060 221546 287112 221552
rect 284668 221468 284720 221474
rect 284668 221410 284720 221416
rect 286508 221332 286560 221338
rect 286508 221274 286560 221280
rect 285680 221264 285732 221270
rect 285680 221206 285732 221212
rect 284484 221128 284536 221134
rect 284484 221070 284536 221076
rect 284852 221060 284904 221066
rect 284852 221002 284904 221008
rect 284392 220924 284444 220930
rect 284392 220866 284444 220872
rect 284864 217410 284892 221002
rect 285692 217410 285720 221206
rect 286520 217410 286548 221274
rect 287336 221128 287388 221134
rect 287336 221070 287388 221076
rect 287348 217410 287376 221070
rect 287808 220998 287836 231474
rect 287900 221202 287928 232970
rect 288268 232898 288296 239686
rect 288636 232966 288664 239686
rect 288624 232960 288676 232966
rect 288624 232902 288676 232908
rect 288256 232892 288308 232898
rect 288256 232834 288308 232840
rect 289004 231538 289032 239686
rect 289372 233034 289400 239686
rect 289820 234660 289872 234666
rect 289820 234602 289872 234608
rect 289360 233028 289412 233034
rect 289360 232970 289412 232976
rect 288992 231532 289044 231538
rect 288992 231474 289044 231480
rect 289728 221400 289780 221406
rect 289728 221342 289780 221348
rect 287888 221196 287940 221202
rect 287888 221138 287940 221144
rect 288256 221196 288308 221202
rect 288256 221138 288308 221144
rect 287796 220992 287848 220998
rect 287796 220934 287848 220940
rect 288268 217410 288296 221138
rect 289084 220992 289136 220998
rect 289084 220934 289136 220940
rect 289096 217410 289124 220934
rect 289740 217410 289768 221342
rect 289832 217546 289860 234602
rect 289924 222766 289952 239700
rect 290108 239686 290306 239714
rect 290476 239686 290674 239714
rect 290752 239686 291042 239714
rect 291120 239686 291410 239714
rect 291488 239686 291778 239714
rect 291856 239686 292146 239714
rect 290004 227180 290056 227186
rect 290004 227122 290056 227128
rect 289912 222760 289964 222766
rect 289912 222702 289964 222708
rect 290016 221134 290044 227122
rect 290108 222426 290136 239686
rect 290280 233096 290332 233102
rect 290280 233038 290332 233044
rect 290188 232960 290240 232966
rect 290188 232902 290240 232908
rect 290096 222420 290148 222426
rect 290096 222362 290148 222368
rect 290004 221128 290056 221134
rect 290004 221070 290056 221076
rect 290200 220998 290228 232902
rect 290292 221066 290320 233038
rect 290372 233028 290424 233034
rect 290372 232970 290424 232976
rect 290384 221338 290412 232970
rect 290372 221332 290424 221338
rect 290372 221274 290424 221280
rect 290476 221270 290504 239686
rect 290752 227186 290780 239686
rect 291120 233102 291148 239686
rect 291108 233096 291160 233102
rect 291108 233038 291160 233044
rect 291488 233034 291516 239686
rect 291476 233028 291528 233034
rect 291476 232970 291528 232976
rect 291856 232966 291884 239686
rect 292408 234666 292436 239700
rect 292790 239686 292896 239714
rect 292580 234728 292632 234734
rect 292580 234670 292632 234676
rect 292396 234660 292448 234666
rect 292396 234602 292448 234608
rect 291844 232960 291896 232966
rect 291844 232902 291896 232908
rect 290740 227180 290792 227186
rect 290740 227122 290792 227128
rect 292396 221332 292448 221338
rect 292396 221274 292448 221280
rect 290464 221264 290516 221270
rect 290464 221206 290516 221212
rect 290280 221060 290332 221066
rect 290280 221002 290332 221008
rect 290188 220992 290240 220998
rect 290188 220934 290240 220940
rect 291568 220992 291620 220998
rect 291568 220934 291620 220940
rect 289832 217518 290044 217546
rect 59984 217382 60320 217410
rect 60812 217382 61148 217410
rect 61640 217382 61976 217410
rect 62468 217382 62804 217410
rect 63296 217382 63448 217410
rect 64216 217382 64552 217410
rect 65044 217382 65380 217410
rect 65872 217382 66208 217410
rect 66700 217382 67036 217410
rect 67528 217382 67864 217410
rect 68356 217382 68692 217410
rect 69184 217382 69520 217410
rect 70104 217382 70440 217410
rect 70932 217382 71268 217410
rect 71760 217382 72096 217410
rect 72588 217382 72924 217410
rect 73416 217382 73752 217410
rect 74244 217382 74488 217410
rect 75072 217382 75408 217410
rect 75992 217382 76328 217410
rect 76820 217382 77156 217410
rect 77648 217382 77984 217410
rect 78476 217382 78812 217410
rect 79304 217382 79640 217410
rect 80132 217382 80468 217410
rect 80960 217382 81296 217410
rect 81880 217382 82216 217410
rect 82708 217382 82768 217410
rect 83536 217382 83872 217410
rect 84364 217382 84700 217410
rect 85192 217382 85528 217410
rect 86020 217382 86356 217410
rect 86848 217382 87184 217410
rect 87768 217382 88104 217410
rect 88596 217382 88932 217410
rect 89424 217382 89760 217410
rect 90252 217382 90588 217410
rect 91080 217382 91416 217410
rect 91908 217382 92244 217410
rect 92736 217382 93072 217410
rect 93656 217382 93808 217410
rect 94484 217382 94820 217410
rect 95312 217382 95648 217410
rect 96140 217382 96476 217410
rect 96968 217382 97304 217410
rect 97796 217382 98132 217410
rect 98624 217382 98960 217410
rect 99544 217382 99880 217410
rect 100372 217382 100708 217410
rect 101200 217382 101536 217410
rect 102028 217382 102088 217410
rect 102856 217382 103192 217410
rect 103684 217382 104020 217410
rect 104512 217382 104848 217410
rect 105432 217382 105768 217410
rect 106260 217382 106596 217410
rect 107088 217382 107424 217410
rect 107916 217382 108252 217410
rect 108744 217382 109080 217410
rect 109572 217382 109908 217410
rect 110400 217382 110736 217410
rect 111320 217382 111656 217410
rect 112148 217382 112484 217410
rect 112976 217382 113128 217410
rect 113804 217382 114140 217410
rect 114632 217382 114968 217410
rect 115460 217382 115796 217410
rect 116288 217382 116624 217410
rect 117208 217382 117544 217410
rect 118036 217382 118372 217410
rect 118864 217382 119200 217410
rect 119692 217382 120028 217410
rect 120520 217382 120856 217410
rect 121348 217382 121408 217410
rect 122176 217382 122512 217410
rect 123096 217382 123432 217410
rect 123924 217382 124168 217410
rect 124752 217382 125088 217410
rect 125580 217382 125916 217410
rect 126408 217382 126744 217410
rect 127236 217382 127572 217410
rect 128064 217382 128400 217410
rect 128984 217382 129320 217410
rect 129812 217382 130148 217410
rect 130640 217382 130976 217410
rect 131468 217382 131804 217410
rect 132296 217382 132448 217410
rect 133124 217382 133460 217410
rect 133952 217382 134288 217410
rect 134872 217382 135208 217410
rect 135700 217382 136036 217410
rect 136528 217382 136864 217410
rect 137356 217382 137692 217410
rect 138184 217382 138520 217410
rect 139012 217382 139256 217410
rect 139840 217382 140176 217410
rect 140760 217382 141096 217410
rect 141588 217382 141924 217410
rect 142416 217382 142752 217410
rect 143244 217382 143488 217410
rect 144072 217382 144408 217410
rect 144900 217382 145236 217410
rect 145728 217382 146064 217410
rect 146648 217382 146984 217410
rect 147476 217382 147812 217410
rect 148304 217382 148640 217410
rect 149132 217382 149468 217410
rect 149960 217382 150296 217410
rect 150788 217382 151124 217410
rect 151616 217382 151768 217410
rect 152536 217382 152872 217410
rect 153364 217382 153700 217410
rect 154192 217382 154528 217410
rect 155020 217382 155356 217410
rect 155848 217382 156184 217410
rect 156676 217382 157012 217410
rect 157504 217382 157840 217410
rect 158424 217382 158760 217410
rect 159252 217382 159588 217410
rect 160080 217382 160416 217410
rect 160908 217382 161244 217410
rect 161736 217382 162072 217410
rect 162564 217382 162808 217410
rect 163392 217382 163728 217410
rect 164312 217382 164648 217410
rect 165140 217382 165476 217410
rect 165968 217382 166304 217410
rect 166796 217382 167132 217410
rect 167624 217382 167960 217410
rect 168452 217382 168788 217410
rect 169280 217382 169616 217410
rect 170200 217382 170536 217410
rect 171028 217382 171088 217410
rect 171856 217382 172192 217410
rect 172684 217382 173020 217410
rect 173512 217382 173756 217410
rect 174340 217382 174676 217410
rect 175168 217382 175504 217410
rect 176088 217382 176424 217410
rect 176916 217382 177252 217410
rect 177744 217382 178080 217410
rect 178572 217382 178908 217410
rect 179400 217382 179736 217410
rect 180228 217382 180564 217410
rect 181056 217382 181392 217410
rect 181976 217382 182128 217410
rect 182804 217382 183140 217410
rect 183632 217382 183968 217410
rect 184460 217382 184796 217410
rect 185288 217382 185624 217410
rect 186116 217382 186452 217410
rect 186944 217382 187280 217410
rect 187864 217382 188200 217410
rect 188692 217382 189028 217410
rect 189520 217382 189856 217410
rect 190348 217382 190408 217410
rect 191176 217382 191512 217410
rect 192004 217382 192340 217410
rect 192832 217382 193076 217410
rect 193752 217382 194088 217410
rect 194580 217382 194916 217410
rect 195408 217382 195744 217410
rect 196236 217382 196572 217410
rect 197064 217382 197400 217410
rect 197892 217382 198228 217410
rect 198720 217382 199056 217410
rect 199640 217382 199976 217410
rect 200468 217382 200804 217410
rect 201296 217382 201356 217410
rect 202124 217382 202460 217410
rect 202952 217382 203288 217410
rect 203780 217382 204208 217410
rect 204608 217382 204944 217410
rect 205528 217382 205864 217410
rect 206356 217382 206692 217410
rect 207184 217382 207428 217410
rect 208012 217382 208348 217410
rect 208840 217382 209176 217410
rect 209668 217382 209728 217410
rect 210496 217382 210832 217410
rect 211416 217382 211752 217410
rect 212244 217382 212396 217410
rect 213072 217382 213408 217410
rect 213900 217382 214236 217410
rect 214728 217382 215064 217410
rect 215556 217382 215892 217410
rect 216384 217382 216720 217410
rect 217304 217382 217732 217410
rect 218132 217382 218376 217410
rect 218960 217382 219296 217410
rect 219788 217382 220124 217410
rect 220616 217382 220768 217410
rect 221444 217382 221780 217410
rect 222272 217382 222608 217410
rect 223192 217382 223528 217410
rect 224020 217382 224356 217410
rect 224848 217382 225184 217410
rect 225676 217382 226104 217410
rect 226504 217382 226840 217410
rect 227332 217382 227668 217410
rect 228160 217382 228496 217410
rect 229080 217382 229416 217410
rect 229908 217382 230244 217410
rect 230736 217382 231072 217410
rect 231564 217382 231808 217410
rect 232392 217382 232728 217410
rect 233220 217382 233556 217410
rect 234048 217382 234384 217410
rect 234968 217382 235304 217410
rect 235796 217382 236132 217410
rect 236624 217382 236960 217410
rect 237452 217382 237788 217410
rect 238280 217382 238616 217410
rect 239108 217382 239444 217410
rect 239936 217382 240088 217410
rect 240856 217382 241192 217410
rect 241684 217382 242020 217410
rect 242512 217382 242756 217410
rect 243340 217382 243676 217410
rect 244168 217382 244504 217410
rect 244996 217382 245424 217410
rect 245824 217382 246160 217410
rect 246744 217382 247080 217410
rect 247572 217382 247908 217410
rect 248400 217382 248736 217410
rect 249228 217382 249564 217410
rect 250056 217382 250392 217410
rect 250884 217382 251036 217410
rect 251712 217382 252048 217410
rect 252632 217382 252968 217410
rect 253460 217382 253888 217410
rect 254288 217382 254624 217410
rect 255116 217382 255452 217410
rect 255944 217382 256280 217410
rect 256772 217382 257108 217410
rect 257600 217382 257936 217410
rect 258520 217382 258856 217410
rect 259348 217382 259408 217410
rect 260176 217382 260512 217410
rect 261004 217382 261340 217410
rect 261832 217382 262168 217410
rect 262660 217382 262996 217410
rect 263488 217382 263824 217410
rect 264408 217382 264836 217410
rect 265236 217382 265572 217410
rect 266064 217382 266400 217410
rect 266892 217382 267320 217410
rect 267720 217382 268056 217410
rect 268548 217382 268884 217410
rect 269376 217382 269712 217410
rect 270296 217382 270448 217410
rect 271124 217382 271460 217410
rect 271952 217382 272288 217410
rect 272780 217382 273116 217410
rect 273608 217382 273944 217410
rect 274436 217382 274772 217410
rect 275264 217382 275600 217410
rect 276184 217382 276520 217410
rect 277012 217382 277348 217410
rect 277840 217382 278176 217410
rect 278668 217382 278728 217410
rect 279496 217382 279832 217410
rect 280324 217382 280660 217410
rect 281152 217382 281488 217410
rect 282072 217382 282408 217410
rect 282900 217382 283236 217410
rect 283728 217382 283972 217410
rect 284556 217382 284892 217410
rect 285384 217382 285720 217410
rect 286212 217382 286548 217410
rect 287040 217382 287376 217410
rect 287960 217382 288296 217410
rect 288788 217382 289124 217410
rect 289616 217382 289768 217410
rect 290016 217410 290044 217518
rect 291580 217410 291608 220934
rect 292408 217410 292436 221274
rect 290016 217382 290444 217410
rect 291272 217382 291608 217410
rect 292100 217382 292436 217410
rect 292592 217410 292620 234670
rect 292672 234660 292724 234666
rect 292672 234602 292724 234608
rect 292684 219586 292712 234602
rect 292764 233028 292816 233034
rect 292764 232970 292816 232976
rect 292776 220998 292804 232970
rect 292868 221202 292896 239686
rect 292960 239686 293158 239714
rect 293236 239686 293526 239714
rect 292960 221406 292988 239686
rect 292948 221400 293000 221406
rect 292948 221342 293000 221348
rect 293236 221338 293264 239686
rect 293880 234666 293908 239700
rect 293972 239686 294262 239714
rect 293868 234660 293920 234666
rect 293868 234602 293920 234608
rect 293972 233034 294000 239686
rect 294616 234734 294644 239700
rect 294604 234728 294656 234734
rect 294604 234670 294656 234676
rect 294984 234666 295012 239700
rect 295260 234734 295288 239700
rect 295352 239686 295642 239714
rect 295720 239686 296010 239714
rect 295248 234728 295300 234734
rect 295248 234670 295300 234676
rect 294972 234660 295024 234666
rect 294972 234602 295024 234608
rect 293960 233028 294012 233034
rect 293960 232970 294012 232976
rect 293224 221332 293276 221338
rect 293224 221274 293276 221280
rect 292856 221196 292908 221202
rect 292856 221138 292908 221144
rect 292764 220992 292816 220998
rect 295352 220946 295380 239686
rect 295432 234660 295484 234666
rect 295432 234602 295484 234608
rect 292764 220934 292816 220940
rect 295076 220918 295380 220946
rect 292684 219558 293448 219586
rect 293420 217410 293448 219558
rect 295076 217410 295104 220918
rect 292592 217382 292928 217410
rect 293420 217382 293848 217410
rect 294676 217382 295104 217410
rect 295444 217410 295472 234602
rect 295720 233050 295748 239686
rect 296364 234802 296392 239700
rect 296352 234796 296404 234802
rect 296352 234738 296404 234744
rect 296732 234734 296760 239700
rect 295892 234728 295944 234734
rect 295892 234670 295944 234676
rect 296720 234728 296772 234734
rect 296720 234670 296772 234676
rect 295800 234660 295852 234666
rect 295800 234602 295852 234608
rect 295628 233022 295748 233050
rect 295628 226334 295656 233022
rect 295628 226306 295748 226334
rect 295720 219722 295748 226306
rect 295812 221338 295840 234602
rect 295904 226334 295932 234670
rect 297100 234666 297128 239700
rect 297482 239686 297772 239714
rect 297744 234682 297772 239686
rect 297836 234870 297864 239700
rect 298112 236026 298140 239700
rect 298100 236020 298152 236026
rect 298100 235962 298152 235968
rect 297824 234864 297876 234870
rect 297824 234806 297876 234812
rect 298192 234796 298244 234802
rect 298192 234738 298244 234744
rect 297088 234660 297140 234666
rect 297744 234654 298140 234682
rect 297088 234602 297140 234608
rect 295904 226306 296760 226334
rect 295800 221332 295852 221338
rect 295800 221274 295852 221280
rect 295720 219694 295932 219722
rect 295904 217410 295932 219694
rect 296732 217410 296760 226306
rect 298112 221406 298140 234654
rect 298100 221400 298152 221406
rect 298100 221342 298152 221348
rect 297640 221332 297692 221338
rect 297640 221274 297692 221280
rect 297652 217410 297680 221274
rect 298204 217410 298232 234738
rect 298480 234734 298508 239700
rect 298284 234728 298336 234734
rect 298284 234670 298336 234676
rect 298468 234728 298520 234734
rect 298468 234670 298520 234676
rect 298296 221338 298324 234670
rect 298848 234666 298876 239700
rect 299216 235754 299244 239700
rect 299204 235748 299256 235754
rect 299204 235690 299256 235696
rect 299584 235618 299612 239700
rect 299952 235890 299980 239700
rect 299940 235884 299992 235890
rect 299940 235826 299992 235832
rect 299572 235612 299624 235618
rect 299572 235554 299624 235560
rect 300320 235550 300348 239700
rect 300308 235544 300360 235550
rect 300308 235486 300360 235492
rect 300688 235074 300716 239700
rect 300964 236094 300992 239700
rect 300952 236088 301004 236094
rect 300952 236030 301004 236036
rect 301332 235686 301360 239700
rect 301700 236978 301728 239700
rect 301688 236972 301740 236978
rect 301688 236914 301740 236920
rect 302068 236434 302096 239700
rect 302436 237182 302464 239700
rect 302424 237176 302476 237182
rect 302424 237118 302476 237124
rect 302804 237046 302832 239700
rect 302792 237040 302844 237046
rect 302792 236982 302844 236988
rect 303172 236706 303200 239700
rect 303160 236700 303212 236706
rect 303160 236642 303212 236648
rect 302056 236428 302108 236434
rect 302056 236370 302108 236376
rect 303540 236366 303568 239700
rect 303528 236360 303580 236366
rect 303528 236302 303580 236308
rect 303816 236230 303844 239700
rect 303804 236224 303856 236230
rect 303804 236166 303856 236172
rect 303804 236020 303856 236026
rect 303804 235962 303856 235968
rect 303712 235748 303764 235754
rect 303712 235690 303764 235696
rect 301320 235680 301372 235686
rect 301320 235622 301372 235628
rect 300676 235068 300728 235074
rect 300676 235010 300728 235016
rect 300860 234864 300912 234870
rect 300860 234806 300912 234812
rect 298836 234660 298888 234666
rect 298836 234602 298888 234608
rect 299388 221400 299440 221406
rect 299388 221342 299440 221348
rect 298284 221332 298336 221338
rect 298284 221274 298336 221280
rect 299400 217410 299428 221342
rect 300872 221338 300900 234806
rect 301044 234728 301096 234734
rect 301044 234670 301096 234676
rect 300952 234660 301004 234666
rect 300952 234602 301004 234608
rect 300964 221406 300992 234602
rect 300952 221400 301004 221406
rect 300952 221342 301004 221348
rect 300216 221332 300268 221338
rect 300216 221274 300268 221280
rect 300860 221332 300912 221338
rect 300860 221274 300912 221280
rect 300228 217410 300256 221274
rect 301056 217410 301084 234670
rect 302700 221400 302752 221406
rect 302700 221342 302752 221348
rect 301872 221332 301924 221338
rect 301872 221274 301924 221280
rect 301884 217410 301912 221274
rect 302712 217410 302740 221342
rect 303724 221338 303752 235690
rect 303712 221332 303764 221338
rect 303712 221274 303764 221280
rect 303816 217410 303844 235962
rect 304080 235884 304132 235890
rect 304080 235826 304132 235832
rect 304092 226334 304120 235826
rect 304184 235006 304212 239700
rect 304172 235000 304224 235006
rect 304172 234942 304224 234948
rect 304552 234938 304580 239700
rect 304920 235278 304948 239700
rect 304908 235272 304960 235278
rect 304908 235214 304960 235220
rect 304540 234932 304592 234938
rect 304540 234874 304592 234880
rect 305288 234666 305316 239700
rect 305656 235142 305684 239700
rect 306024 235210 306052 239700
rect 306392 235346 306420 239700
rect 306668 235686 306696 239700
rect 306656 235680 306708 235686
rect 306656 235622 306708 235628
rect 306656 235544 306708 235550
rect 306656 235486 306708 235492
rect 306380 235340 306432 235346
rect 306380 235282 306432 235288
rect 306012 235204 306064 235210
rect 306012 235146 306064 235152
rect 305644 235136 305696 235142
rect 305644 235078 305696 235084
rect 305276 234660 305328 234666
rect 305276 234602 305328 234608
rect 306288 234660 306340 234666
rect 306288 234602 306340 234608
rect 304092 226306 304304 226334
rect 304276 217410 304304 226306
rect 305276 221332 305328 221338
rect 305276 221274 305328 221280
rect 305288 217410 305316 221274
rect 306300 221066 306328 234602
rect 306288 221060 306340 221066
rect 306288 221002 306340 221008
rect 306668 217410 306696 235486
rect 307036 235074 307064 239700
rect 307300 235748 307352 235754
rect 307300 235690 307352 235696
rect 307208 235612 307260 235618
rect 307208 235554 307260 235560
rect 306748 235068 306800 235074
rect 306748 235010 306800 235016
rect 307024 235068 307076 235074
rect 307024 235010 307076 235016
rect 306760 221338 306788 235010
rect 306748 221332 306800 221338
rect 306748 221274 306800 221280
rect 295444 217382 295504 217410
rect 295904 217382 296332 217410
rect 296732 217382 297160 217410
rect 297652 217382 297988 217410
rect 298204 217382 298816 217410
rect 299400 217382 299736 217410
rect 300228 217382 300564 217410
rect 301056 217382 301392 217410
rect 301884 217382 302220 217410
rect 302712 217382 303048 217410
rect 303816 217382 303876 217410
rect 304276 217382 304704 217410
rect 305288 217382 305624 217410
rect 306452 217382 306696 217410
rect 307220 217410 307248 235554
rect 307312 226334 307340 235690
rect 307404 234802 307432 239700
rect 307392 234796 307444 234802
rect 307392 234738 307444 234744
rect 307772 234666 307800 239700
rect 308140 234734 308168 239700
rect 308522 239686 308720 239714
rect 308890 239686 309088 239714
rect 308128 234728 308180 234734
rect 308128 234670 308180 234676
rect 307760 234660 307812 234666
rect 307760 234602 307812 234608
rect 308496 234660 308548 234666
rect 308496 234602 308548 234608
rect 307312 226306 307708 226334
rect 307680 217410 307708 226306
rect 308508 222630 308536 234602
rect 308692 222834 308720 239686
rect 308772 235680 308824 235686
rect 308772 235622 308824 235628
rect 308784 223038 308812 235622
rect 308956 234796 309008 234802
rect 308956 234738 309008 234744
rect 308864 234728 308916 234734
rect 308864 234670 308916 234676
rect 308772 223032 308824 223038
rect 308772 222974 308824 222980
rect 308680 222828 308732 222834
rect 308680 222770 308732 222776
rect 308876 222766 308904 234670
rect 308968 223174 308996 234738
rect 308956 223168 309008 223174
rect 308956 223110 309008 223116
rect 309060 222902 309088 239686
rect 309244 236162 309272 239700
rect 309232 236156 309284 236162
rect 309232 236098 309284 236104
rect 309416 236088 309468 236094
rect 309416 236030 309468 236036
rect 309048 222896 309100 222902
rect 309048 222838 309100 222844
rect 308864 222760 308916 222766
rect 308864 222702 308916 222708
rect 308496 222624 308548 222630
rect 308496 222566 308548 222572
rect 309428 221338 309456 236030
rect 309520 234870 309548 239700
rect 309784 237040 309836 237046
rect 309784 236982 309836 236988
rect 309508 234864 309560 234870
rect 309508 234806 309560 234812
rect 309796 221406 309824 236982
rect 309888 234802 309916 239700
rect 309968 236972 310020 236978
rect 309968 236914 310020 236920
rect 309876 234796 309928 234802
rect 309876 234738 309928 234744
rect 309784 221400 309836 221406
rect 309784 221342 309836 221348
rect 308588 221332 308640 221338
rect 308588 221274 308640 221280
rect 309416 221332 309468 221338
rect 309416 221274 309468 221280
rect 308600 217410 308628 221274
rect 309980 217410 310008 236914
rect 310256 234734 310284 239700
rect 310624 235958 310652 239700
rect 310612 235952 310664 235958
rect 310612 235894 310664 235900
rect 310244 234728 310296 234734
rect 310244 234670 310296 234676
rect 310992 234666 311020 239700
rect 310980 234660 311032 234666
rect 310980 234602 311032 234608
rect 311360 222494 311388 239700
rect 311544 239686 311742 239714
rect 311440 234728 311492 234734
rect 311440 234670 311492 234676
rect 311452 222698 311480 234670
rect 311440 222692 311492 222698
rect 311440 222634 311492 222640
rect 311544 222562 311572 239686
rect 312096 237250 312124 239700
rect 312084 237244 312136 237250
rect 312084 237186 312136 237192
rect 312268 236428 312320 236434
rect 312268 236370 312320 236376
rect 311716 234864 311768 234870
rect 311716 234806 311768 234812
rect 311624 234660 311676 234666
rect 311624 234602 311676 234608
rect 311532 222556 311584 222562
rect 311532 222498 311584 222504
rect 311348 222488 311400 222494
rect 311348 222430 311400 222436
rect 311636 222358 311664 234602
rect 311728 223106 311756 234806
rect 311808 234796 311860 234802
rect 311808 234738 311860 234744
rect 311716 223100 311768 223106
rect 311716 223042 311768 223048
rect 311624 222352 311676 222358
rect 311624 222294 311676 222300
rect 311164 221400 311216 221406
rect 311164 221342 311216 221348
rect 310244 221332 310296 221338
rect 310244 221274 310296 221280
rect 307220 217382 307280 217410
rect 307680 217382 308108 217410
rect 308600 217382 308936 217410
rect 309764 217382 310008 217410
rect 310256 217410 310284 221274
rect 311176 217410 311204 221342
rect 311820 220998 311848 234738
rect 311808 220992 311860 220998
rect 311808 220934 311860 220940
rect 312280 217410 312308 236370
rect 312372 234870 312400 239700
rect 312636 236700 312688 236706
rect 312636 236642 312688 236648
rect 312360 234864 312412 234870
rect 312360 234806 312412 234812
rect 312648 226334 312676 236642
rect 312740 234734 312768 239700
rect 312820 237176 312872 237182
rect 312820 237118 312872 237124
rect 312728 234728 312780 234734
rect 312728 234670 312780 234676
rect 312832 226334 312860 237118
rect 313108 234802 313136 239700
rect 313476 236026 313504 239700
rect 313464 236020 313516 236026
rect 313464 235962 313516 235968
rect 313096 234796 313148 234802
rect 313096 234738 313148 234744
rect 313844 234666 313872 239700
rect 314226 239686 314332 239714
rect 314016 234864 314068 234870
rect 314016 234806 314068 234812
rect 313832 234660 313884 234666
rect 313832 234602 313884 234608
rect 314028 232966 314056 234806
rect 314108 234728 314160 234734
rect 314108 234670 314160 234676
rect 314200 234728 314252 234734
rect 314200 234670 314252 234676
rect 314016 232960 314068 232966
rect 314016 232902 314068 232908
rect 312648 226306 312768 226334
rect 312832 226306 313596 226334
rect 312740 217410 312768 226306
rect 313568 217410 313596 226306
rect 314120 222426 314148 234670
rect 314212 223446 314240 234670
rect 314200 223440 314252 223446
rect 314200 223382 314252 223388
rect 314108 222420 314160 222426
rect 314108 222362 314160 222368
rect 314304 222290 314332 239686
rect 314476 234796 314528 234802
rect 314476 234738 314528 234744
rect 314384 234660 314436 234666
rect 314384 234602 314436 234608
rect 314292 222284 314344 222290
rect 314292 222226 314344 222232
rect 314396 221542 314424 234602
rect 314488 233050 314516 234738
rect 314580 234734 314608 239700
rect 314948 237318 314976 239700
rect 314936 237312 314988 237318
rect 314936 237254 314988 237260
rect 315028 236360 315080 236366
rect 315028 236302 315080 236308
rect 314568 234728 314620 234734
rect 314568 234670 314620 234676
rect 314488 233022 314608 233050
rect 314476 232960 314528 232966
rect 314476 232902 314528 232908
rect 314384 221536 314436 221542
rect 314384 221478 314436 221484
rect 314488 221202 314516 232902
rect 314476 221196 314528 221202
rect 314476 221138 314528 221144
rect 314580 221134 314608 233022
rect 315040 221406 315068 236302
rect 315224 234870 315252 239700
rect 315396 235000 315448 235006
rect 315396 234942 315448 234948
rect 315304 234932 315356 234938
rect 315304 234874 315356 234880
rect 315212 234864 315264 234870
rect 315212 234806 315264 234812
rect 315028 221400 315080 221406
rect 315028 221342 315080 221348
rect 315316 221338 315344 234874
rect 315304 221332 315356 221338
rect 315304 221274 315356 221280
rect 314568 221128 314620 221134
rect 314568 221070 314620 221076
rect 315408 217546 315436 234942
rect 315592 234666 315620 239700
rect 315960 234802 315988 239700
rect 316328 236434 316356 239700
rect 316316 236428 316368 236434
rect 316316 236370 316368 236376
rect 315948 234796 316000 234802
rect 315948 234738 316000 234744
rect 316696 234734 316724 239700
rect 316684 234728 316736 234734
rect 316684 234670 316736 234676
rect 315580 234660 315632 234666
rect 315580 234602 315632 234608
rect 316960 234660 317012 234666
rect 316960 234602 317012 234608
rect 315488 221400 315540 221406
rect 315488 221342 315540 221348
rect 315132 217518 315436 217546
rect 315132 217410 315160 217518
rect 310256 217382 310592 217410
rect 311176 217382 311512 217410
rect 312280 217382 312340 217410
rect 312740 217382 313168 217410
rect 313568 217382 313996 217410
rect 314824 217382 315160 217410
rect 315500 217410 315528 221342
rect 316132 221332 316184 221338
rect 316132 221274 316184 221280
rect 316144 217410 316172 221274
rect 316972 221270 317000 234602
rect 317064 222222 317092 239700
rect 317432 237182 317460 239700
rect 317420 237176 317472 237182
rect 317420 237118 317472 237124
rect 317800 236502 317828 239700
rect 317788 236496 317840 236502
rect 317788 236438 317840 236444
rect 317972 236224 318024 236230
rect 317972 236166 318024 236172
rect 317880 235272 317932 235278
rect 317880 235214 317932 235220
rect 317788 235204 317840 235210
rect 317788 235146 317840 235152
rect 317696 235136 317748 235142
rect 317696 235078 317748 235084
rect 317144 234864 317196 234870
rect 317144 234806 317196 234812
rect 317052 222216 317104 222222
rect 317052 222158 317104 222164
rect 317156 221814 317184 234806
rect 317328 234796 317380 234802
rect 317328 234738 317380 234744
rect 317236 234728 317288 234734
rect 317236 234670 317288 234676
rect 317248 222970 317276 234670
rect 317236 222964 317288 222970
rect 317236 222906 317288 222912
rect 317144 221808 317196 221814
rect 317144 221750 317196 221756
rect 317340 221474 317368 234738
rect 317328 221468 317380 221474
rect 317328 221410 317380 221416
rect 317604 221332 317656 221338
rect 317604 221274 317656 221280
rect 316960 221264 317012 221270
rect 316960 221206 317012 221212
rect 317616 217410 317644 221274
rect 315500 217382 315652 217410
rect 316144 217382 316480 217410
rect 317400 217382 317644 217410
rect 317708 217410 317736 235078
rect 317800 221406 317828 235146
rect 317788 221400 317840 221406
rect 317788 221342 317840 221348
rect 317892 220538 317920 235214
rect 317984 221338 318012 236166
rect 318076 234802 318104 239700
rect 318064 234796 318116 234802
rect 318064 234738 318116 234744
rect 318444 234734 318472 239700
rect 318812 236910 318840 239700
rect 318800 236904 318852 236910
rect 318800 236846 318852 236852
rect 319180 236366 319208 239700
rect 319168 236360 319220 236366
rect 319168 236302 319220 236308
rect 318432 234728 318484 234734
rect 318432 234670 318484 234676
rect 319548 234666 319576 239700
rect 319824 239686 319930 239714
rect 319536 234660 319588 234666
rect 319536 234602 319588 234608
rect 319824 221678 319852 239686
rect 320284 236842 320312 239700
rect 320272 236836 320324 236842
rect 320272 236778 320324 236784
rect 320652 236298 320680 239700
rect 320640 236292 320692 236298
rect 320640 236234 320692 236240
rect 320824 235068 320876 235074
rect 320824 235010 320876 235016
rect 320088 234796 320140 234802
rect 320088 234738 320140 234744
rect 319904 234728 319956 234734
rect 319904 234670 319956 234676
rect 319812 221672 319864 221678
rect 319812 221614 319864 221620
rect 319916 221474 319944 234670
rect 319996 234660 320048 234666
rect 319996 234602 320048 234608
rect 320008 221950 320036 234602
rect 319996 221944 320048 221950
rect 319996 221886 320048 221892
rect 320100 221610 320128 234738
rect 320836 226334 320864 235010
rect 320928 234870 320956 239700
rect 321008 235340 321060 235346
rect 321008 235282 321060 235288
rect 320916 234864 320968 234870
rect 320916 234806 320968 234812
rect 321020 226334 321048 235282
rect 321296 234734 321324 239700
rect 321664 234802 321692 239700
rect 322032 236230 322060 239700
rect 322020 236224 322072 236230
rect 322020 236166 322072 236172
rect 321652 234796 321704 234802
rect 321652 234738 321704 234744
rect 321284 234728 321336 234734
rect 321284 234670 321336 234676
rect 322400 234666 322428 239700
rect 322584 239686 322782 239714
rect 322480 234728 322532 234734
rect 322480 234670 322532 234676
rect 322388 234660 322440 234666
rect 322388 234602 322440 234608
rect 320836 226306 320956 226334
rect 321020 226306 321968 226334
rect 320088 221604 320140 221610
rect 320088 221546 320140 221552
rect 319904 221468 319956 221474
rect 319904 221410 319956 221416
rect 319536 221400 319588 221406
rect 319536 221342 319588 221348
rect 320928 221354 320956 226306
rect 317972 221332 318024 221338
rect 317972 221274 318024 221280
rect 317892 220510 318656 220538
rect 318628 217410 318656 220510
rect 319548 217410 319576 221342
rect 320928 221326 321140 221354
rect 320364 221060 320416 221066
rect 320364 221002 320416 221008
rect 320376 217410 320404 221002
rect 321112 217410 321140 221326
rect 321940 217410 321968 226306
rect 322492 221746 322520 234670
rect 322584 222086 322612 239686
rect 323136 235006 323164 239700
rect 323124 235000 323176 235006
rect 323124 234942 323176 234948
rect 322848 234864 322900 234870
rect 322848 234806 322900 234812
rect 322756 234796 322808 234802
rect 322756 234738 322808 234744
rect 322664 234660 322716 234666
rect 322664 234602 322716 234608
rect 322676 222154 322704 234602
rect 322664 222148 322716 222154
rect 322664 222090 322716 222096
rect 322572 222080 322624 222086
rect 322572 222022 322624 222028
rect 322768 222018 322796 234738
rect 322756 222012 322808 222018
rect 322756 221954 322808 221960
rect 322860 221882 322888 234806
rect 323504 234666 323532 239700
rect 323780 234734 323808 239700
rect 324148 234870 324176 239700
rect 324516 236774 324544 239700
rect 324504 236768 324556 236774
rect 324504 236710 324556 236716
rect 324136 234864 324188 234870
rect 324136 234806 324188 234812
rect 324884 234802 324912 239700
rect 324872 234796 324924 234802
rect 324872 234738 324924 234744
rect 323768 234728 323820 234734
rect 323768 234670 323820 234676
rect 323492 234660 323544 234666
rect 323492 234602 323544 234608
rect 325148 234660 325200 234666
rect 325148 234602 325200 234608
rect 325160 223514 325188 234602
rect 325148 223508 325200 223514
rect 325148 223450 325200 223456
rect 323124 223168 323176 223174
rect 323124 223110 323176 223116
rect 322848 221876 322900 221882
rect 322848 221818 322900 221824
rect 322480 221740 322532 221746
rect 322480 221682 322532 221688
rect 323136 217410 323164 223110
rect 323768 223032 323820 223038
rect 323768 222974 323820 222980
rect 323780 217410 323808 222974
rect 325252 222834 325280 239700
rect 325436 239686 325634 239714
rect 325332 234728 325384 234734
rect 325332 234670 325384 234676
rect 325344 223038 325372 234670
rect 325436 223174 325464 239686
rect 325988 236978 326016 239700
rect 325976 236972 326028 236978
rect 325976 236914 326028 236920
rect 326356 234870 326384 239700
rect 325516 234864 325568 234870
rect 325516 234806 325568 234812
rect 326344 234864 326396 234870
rect 326344 234806 326396 234812
rect 325528 223582 325556 234806
rect 325608 234796 325660 234802
rect 325608 234738 325660 234744
rect 325516 223576 325568 223582
rect 325516 223518 325568 223524
rect 325620 223242 325648 234738
rect 326632 234666 326660 239700
rect 327000 234802 327028 239700
rect 326988 234796 327040 234802
rect 326988 234738 327040 234744
rect 327368 234734 327396 239700
rect 327750 239686 328040 239714
rect 327356 234728 327408 234734
rect 327356 234670 327408 234676
rect 326620 234660 326672 234666
rect 326620 234602 326672 234608
rect 327908 234660 327960 234666
rect 327908 234602 327960 234608
rect 325608 223236 325660 223242
rect 325608 223178 325660 223184
rect 325424 223168 325476 223174
rect 325424 223110 325476 223116
rect 325332 223032 325384 223038
rect 325332 222974 325384 222980
rect 326252 222896 326304 222902
rect 326252 222838 326304 222844
rect 324596 222828 324648 222834
rect 324596 222770 324648 222776
rect 325240 222828 325292 222834
rect 325240 222770 325292 222776
rect 324608 217410 324636 222770
rect 325700 222624 325752 222630
rect 325700 222566 325752 222572
rect 325712 217410 325740 222566
rect 326264 217410 326292 222838
rect 327920 222766 327948 234602
rect 327080 222760 327132 222766
rect 327080 222702 327132 222708
rect 327908 222760 327960 222766
rect 327908 222702 327960 222708
rect 327092 217410 327120 222702
rect 328012 222630 328040 239686
rect 328104 222873 328132 239700
rect 328472 234870 328500 239700
rect 328644 236156 328696 236162
rect 328644 236098 328696 236104
rect 328184 234864 328236 234870
rect 328184 234806 328236 234812
rect 328460 234864 328512 234870
rect 328460 234806 328512 234812
rect 328196 223378 328224 234806
rect 328276 234796 328328 234802
rect 328276 234738 328328 234744
rect 328184 223372 328236 223378
rect 328184 223314 328236 223320
rect 328288 223310 328316 234738
rect 328368 234728 328420 234734
rect 328368 234670 328420 234676
rect 328276 223304 328328 223310
rect 328276 223246 328328 223252
rect 328380 222902 328408 234670
rect 328656 226334 328684 236098
rect 328840 235074 328868 239700
rect 329208 237386 329236 239700
rect 329196 237380 329248 237386
rect 329196 237322 329248 237328
rect 328828 235068 328880 235074
rect 328828 235010 328880 235016
rect 329484 234802 329512 239700
rect 329748 237176 329800 237182
rect 329748 237118 329800 237124
rect 329472 234796 329524 234802
rect 329472 234738 329524 234744
rect 328656 226306 328776 226334
rect 328368 222896 328420 222902
rect 328090 222864 328146 222873
rect 328368 222838 328420 222844
rect 328090 222799 328146 222808
rect 328000 222624 328052 222630
rect 328000 222566 328052 222572
rect 327908 220992 327960 220998
rect 327908 220934 327960 220940
rect 327920 217410 327948 220934
rect 328748 217410 328776 226306
rect 329656 222692 329708 222698
rect 329656 222634 329708 222640
rect 329668 217410 329696 222634
rect 329760 221066 329788 237118
rect 329852 234666 329880 239700
rect 330220 234734 330248 239700
rect 330588 236094 330616 239700
rect 330576 236088 330628 236094
rect 330576 236030 330628 236036
rect 330852 234864 330904 234870
rect 330852 234806 330904 234812
rect 330208 234728 330260 234734
rect 330208 234670 330260 234676
rect 329840 234660 329892 234666
rect 329840 234602 329892 234608
rect 330760 234660 330812 234666
rect 330760 234602 330812 234608
rect 330484 223100 330536 223106
rect 330484 223042 330536 223048
rect 329748 221060 329800 221066
rect 329748 221002 329800 221008
rect 330496 217410 330524 223042
rect 330772 222737 330800 234602
rect 330864 223106 330892 234806
rect 330852 223100 330904 223106
rect 330852 223042 330904 223048
rect 330758 222728 330814 222737
rect 330758 222663 330814 222672
rect 330956 222601 330984 239700
rect 331324 234870 331352 239700
rect 331692 235618 331720 239700
rect 331772 235952 331824 235958
rect 331772 235894 331824 235900
rect 331680 235612 331732 235618
rect 331680 235554 331732 235560
rect 331312 234864 331364 234870
rect 331312 234806 331364 234812
rect 331128 234796 331180 234802
rect 331128 234738 331180 234744
rect 331036 234728 331088 234734
rect 331036 234670 331088 234676
rect 331048 223145 331076 234670
rect 331034 223136 331090 223145
rect 331034 223071 331090 223080
rect 331140 223009 331168 234738
rect 331784 226334 331812 235894
rect 332060 234734 332088 239700
rect 332048 234728 332100 234734
rect 332048 234670 332100 234676
rect 332336 234666 332364 239700
rect 332704 234802 332732 239700
rect 333072 235414 333100 239700
rect 333060 235408 333112 235414
rect 333060 235350 333112 235356
rect 332692 234796 332744 234802
rect 332692 234738 332744 234744
rect 332324 234660 332376 234666
rect 332324 234602 332376 234608
rect 331784 226306 332088 226334
rect 331126 223000 331182 223009
rect 331126 222935 331182 222944
rect 330942 222592 330998 222601
rect 330942 222527 330998 222536
rect 331312 222488 331364 222494
rect 331312 222430 331364 222436
rect 331324 217410 331352 222430
rect 332060 217410 332088 226306
rect 333440 223990 333468 239700
rect 333716 239686 333822 239714
rect 333520 234728 333572 234734
rect 333520 234670 333572 234676
rect 333428 223984 333480 223990
rect 333428 223926 333480 223932
rect 333532 223922 333560 234670
rect 333612 234660 333664 234666
rect 333612 234602 333664 234608
rect 333520 223916 333572 223922
rect 333520 223858 333572 223864
rect 332968 222556 333020 222562
rect 332968 222498 333020 222504
rect 332980 217410 333008 222498
rect 333624 222465 333652 234602
rect 333610 222456 333666 222465
rect 333610 222391 333666 222400
rect 333716 222329 333744 239686
rect 333796 234864 333848 234870
rect 333796 234806 333848 234812
rect 333808 222698 333836 234806
rect 333888 234796 333940 234802
rect 333888 234738 333940 234744
rect 333796 222692 333848 222698
rect 333796 222634 333848 222640
rect 333900 222562 333928 234738
rect 334176 234734 334204 239700
rect 334440 237244 334492 237250
rect 334440 237186 334492 237192
rect 334164 234728 334216 234734
rect 334164 234670 334216 234676
rect 334452 226334 334480 237186
rect 334544 235958 334572 239700
rect 334532 235952 334584 235958
rect 334532 235894 334584 235900
rect 334912 230722 334940 239700
rect 335202 239686 335492 239714
rect 335464 232966 335492 239686
rect 335556 234666 335584 239700
rect 335938 239686 336228 239714
rect 336096 234728 336148 234734
rect 336096 234670 336148 234676
rect 335544 234660 335596 234666
rect 335544 234602 335596 234608
rect 335452 232960 335504 232966
rect 335452 232902 335504 232908
rect 334900 230716 334952 230722
rect 334900 230658 334952 230664
rect 334452 226306 335492 226334
rect 333888 222556 333940 222562
rect 333888 222498 333940 222504
rect 334716 222420 334768 222426
rect 334716 222362 334768 222368
rect 333980 222352 334032 222358
rect 333702 222320 333758 222329
rect 333980 222294 334032 222300
rect 333702 222255 333758 222264
rect 333992 217410 334020 222294
rect 334728 217410 334756 222362
rect 335464 217410 335492 226306
rect 336108 222494 336136 234670
rect 336096 222488 336148 222494
rect 336096 222430 336148 222436
rect 336200 222057 336228 239686
rect 336292 234938 336320 239700
rect 336384 239686 336674 239714
rect 336280 234932 336332 234938
rect 336280 234874 336332 234880
rect 336384 233050 336412 239686
rect 336648 234932 336700 234938
rect 336648 234874 336700 234880
rect 336464 234660 336516 234666
rect 336464 234602 336516 234608
rect 336292 233022 336412 233050
rect 336292 224262 336320 233022
rect 336372 232960 336424 232966
rect 336372 232902 336424 232908
rect 336280 224256 336332 224262
rect 336280 224198 336332 224204
rect 336384 224058 336412 232902
rect 336372 224052 336424 224058
rect 336372 223994 336424 224000
rect 336476 222426 336504 234602
rect 336660 230654 336688 234874
rect 337028 234802 337056 239700
rect 337108 236020 337160 236026
rect 337108 235962 337160 235968
rect 337016 234796 337068 234802
rect 337016 234738 337068 234744
rect 336648 230648 336700 230654
rect 336648 230590 336700 230596
rect 336464 222420 336516 222426
rect 336464 222362 336516 222368
rect 336186 222048 336242 222057
rect 336186 221983 336242 221992
rect 337120 221338 337148 235962
rect 337396 234734 337424 239700
rect 337384 234728 337436 234734
rect 337384 234670 337436 234676
rect 337764 230586 337792 239700
rect 338040 234666 338068 239700
rect 338120 236904 338172 236910
rect 338120 236846 338172 236852
rect 338028 234660 338080 234666
rect 338028 234602 338080 234608
rect 337752 230580 337804 230586
rect 337752 230522 337804 230528
rect 338028 222284 338080 222290
rect 338028 222226 338080 222232
rect 337108 221332 337160 221338
rect 337108 221274 337160 221280
rect 336740 221196 336792 221202
rect 336740 221138 336792 221144
rect 336752 217410 336780 221138
rect 337200 221128 337252 221134
rect 337200 221070 337252 221076
rect 317708 217382 318228 217410
rect 318628 217382 319056 217410
rect 319548 217382 319884 217410
rect 320376 217382 320712 217410
rect 321112 217382 321540 217410
rect 321940 217382 322368 217410
rect 323136 217382 323288 217410
rect 323780 217382 324116 217410
rect 324608 217382 324944 217410
rect 325712 217382 325772 217410
rect 326264 217382 326600 217410
rect 327092 217382 327428 217410
rect 327920 217382 328256 217410
rect 328748 217382 329176 217410
rect 329668 217382 330004 217410
rect 330496 217382 330832 217410
rect 331324 217382 331660 217410
rect 332060 217382 332488 217410
rect 332980 217382 333316 217410
rect 333992 217382 334144 217410
rect 334728 217382 335064 217410
rect 335464 217382 335892 217410
rect 336720 217382 336780 217410
rect 337212 217410 337240 221070
rect 338040 217410 338068 222226
rect 338132 221134 338160 236846
rect 338408 236026 338436 239700
rect 338790 239686 339080 239714
rect 339158 239686 339448 239714
rect 338396 236020 338448 236026
rect 338396 235962 338448 235968
rect 339052 234954 339080 239686
rect 339052 234926 339356 234954
rect 339224 234796 339276 234802
rect 339224 234738 339276 234744
rect 338856 234728 338908 234734
rect 338856 234670 338908 234676
rect 338868 222358 338896 234670
rect 338948 234660 339000 234666
rect 338948 234602 339000 234608
rect 338960 232914 338988 234602
rect 338960 232886 339172 232914
rect 339144 224194 339172 232886
rect 339132 224188 339184 224194
rect 339132 224130 339184 224136
rect 338856 222352 338908 222358
rect 338856 222294 338908 222300
rect 339236 222290 339264 234738
rect 339328 223553 339356 234926
rect 339420 230382 339448 239686
rect 339512 234802 339540 239700
rect 339500 234796 339552 234802
rect 339500 234738 339552 234744
rect 339408 230376 339460 230382
rect 339408 230318 339460 230324
rect 339880 226710 339908 239700
rect 340248 234666 340276 239700
rect 340616 234734 340644 239700
rect 340906 239686 341196 239714
rect 340880 236836 340932 236842
rect 340880 236778 340932 236784
rect 340788 235000 340840 235006
rect 340788 234942 340840 234948
rect 340604 234728 340656 234734
rect 340604 234670 340656 234676
rect 340236 234660 340288 234666
rect 340236 234602 340288 234608
rect 339868 226704 339920 226710
rect 339868 226646 339920 226652
rect 339314 223544 339370 223553
rect 339314 223479 339370 223488
rect 339684 223440 339736 223446
rect 339684 223382 339736 223388
rect 339224 222284 339276 222290
rect 339224 222226 339276 222232
rect 338856 221332 338908 221338
rect 338856 221274 338908 221280
rect 338120 221128 338172 221134
rect 338120 221070 338172 221076
rect 338868 217410 338896 221274
rect 339696 217410 339724 223382
rect 340604 221536 340656 221542
rect 340604 221478 340656 221484
rect 340616 217410 340644 221478
rect 340800 221338 340828 234942
rect 340788 221332 340840 221338
rect 340788 221274 340840 221280
rect 340892 221270 340920 236778
rect 341168 224398 341196 239686
rect 341260 226778 341288 239700
rect 341642 239686 341748 239714
rect 341616 234660 341668 234666
rect 341616 234602 341668 234608
rect 341248 226772 341300 226778
rect 341248 226714 341300 226720
rect 341156 224392 341208 224398
rect 341156 224334 341208 224340
rect 341628 222193 341656 234602
rect 341720 231810 341748 239686
rect 341904 239686 342010 239714
rect 341800 234796 341852 234802
rect 341800 234738 341852 234744
rect 341708 231804 341760 231810
rect 341708 231746 341760 231752
rect 341812 224126 341840 234738
rect 341904 224534 341932 239686
rect 342364 234802 342392 239700
rect 342746 239686 343036 239714
rect 342720 237312 342772 237318
rect 342720 237254 342772 237260
rect 342352 234796 342404 234802
rect 342352 234738 342404 234744
rect 341984 234728 342036 234734
rect 341984 234670 342036 234676
rect 341892 224528 341944 224534
rect 341892 224470 341944 224476
rect 341996 224466 342024 234670
rect 341984 224460 342036 224466
rect 341984 224402 342036 224408
rect 341800 224120 341852 224126
rect 341800 224062 341852 224068
rect 341614 222184 341670 222193
rect 341614 222119 341670 222128
rect 340880 221264 340932 221270
rect 340880 221206 340932 221212
rect 341432 221196 341484 221202
rect 341432 221138 341484 221144
rect 341444 217410 341472 221138
rect 342732 217410 342760 237254
rect 343008 226846 343036 239686
rect 343100 234870 343128 239700
rect 343364 236972 343416 236978
rect 343364 236914 343416 236920
rect 343272 236768 343324 236774
rect 343272 236710 343324 236716
rect 343088 234864 343140 234870
rect 343088 234806 343140 234812
rect 342996 226840 343048 226846
rect 342996 226782 343048 226788
rect 343088 221400 343140 221406
rect 343088 221342 343140 221348
rect 337212 217382 337548 217410
rect 338040 217382 338376 217410
rect 338868 217382 339204 217410
rect 339696 217382 340032 217410
rect 340616 217382 340952 217410
rect 341444 217382 341780 217410
rect 342608 217382 342760 217410
rect 343100 217410 343128 221342
rect 343284 220998 343312 236710
rect 343376 231792 343404 236914
rect 343468 234734 343496 239700
rect 343640 235068 343692 235074
rect 343640 235010 343692 235016
rect 343456 234728 343508 234734
rect 343456 234670 343508 234676
rect 343652 234546 343680 235010
rect 343744 234666 343772 239700
rect 343732 234660 343784 234666
rect 343732 234602 343784 234608
rect 343652 234518 343772 234546
rect 343376 231764 343680 231792
rect 343652 221406 343680 231764
rect 343744 221542 343772 234518
rect 344112 226914 344140 239700
rect 344376 234796 344428 234802
rect 344376 234738 344428 234744
rect 344100 226908 344152 226914
rect 344100 226850 344152 226856
rect 344388 224330 344416 234738
rect 344480 227050 344508 239700
rect 344756 239686 344862 239714
rect 344652 234728 344704 234734
rect 344652 234670 344704 234676
rect 344468 227044 344520 227050
rect 344468 226986 344520 226992
rect 344664 224602 344692 234670
rect 344756 224738 344784 239686
rect 345216 234802 345244 239700
rect 345388 236428 345440 236434
rect 345388 236370 345440 236376
rect 345204 234796 345256 234802
rect 345204 234738 345256 234744
rect 344836 234660 344888 234666
rect 344836 234602 344888 234608
rect 344848 224806 344876 234602
rect 345400 226334 345428 236370
rect 345584 226982 345612 239700
rect 345952 227254 345980 239700
rect 346216 235408 346268 235414
rect 346216 235350 346268 235356
rect 345940 227248 345992 227254
rect 345940 227190 345992 227196
rect 345572 226976 345624 226982
rect 345572 226918 345624 226924
rect 345400 226306 345520 226334
rect 344836 224800 344888 224806
rect 344836 224742 344888 224748
rect 344744 224732 344796 224738
rect 344744 224674 344796 224680
rect 344652 224596 344704 224602
rect 344652 224538 344704 224544
rect 344376 224324 344428 224330
rect 344376 224266 344428 224272
rect 345020 222216 345072 222222
rect 345020 222158 345072 222164
rect 343916 221808 343968 221814
rect 343916 221750 343968 221756
rect 343732 221536 343784 221542
rect 343732 221478 343784 221484
rect 343640 221400 343692 221406
rect 343640 221342 343692 221348
rect 343272 220992 343324 220998
rect 343272 220934 343324 220940
rect 343928 217410 343956 221750
rect 345032 217410 345060 222158
rect 345492 217410 345520 226306
rect 346228 223446 346256 235350
rect 346320 234734 346348 239700
rect 346492 235952 346544 235958
rect 346492 235894 346544 235900
rect 346400 235612 346452 235618
rect 346400 235554 346452 235560
rect 346308 234728 346360 234734
rect 346308 234670 346360 234676
rect 346216 223440 346268 223446
rect 346216 223382 346268 223388
rect 346412 221814 346440 235554
rect 346504 224516 346532 235894
rect 346596 234666 346624 239700
rect 346584 234660 346636 234666
rect 346584 234602 346636 234608
rect 346964 227118 346992 239700
rect 347044 234932 347096 234938
rect 347044 234874 347096 234880
rect 346952 227112 347004 227118
rect 346952 227054 347004 227060
rect 347056 226166 347084 234874
rect 347332 234802 347360 239700
rect 347700 234938 347728 239700
rect 347688 234932 347740 234938
rect 347688 234874 347740 234880
rect 348068 234802 348096 239700
rect 348148 236496 348200 236502
rect 348148 236438 348200 236444
rect 347136 234796 347188 234802
rect 347136 234738 347188 234744
rect 347320 234796 347372 234802
rect 347320 234738 347372 234744
rect 347688 234796 347740 234802
rect 347688 234738 347740 234744
rect 348056 234796 348108 234802
rect 348056 234738 348108 234744
rect 347044 226160 347096 226166
rect 347044 226102 347096 226108
rect 347148 224670 347176 234738
rect 347596 234728 347648 234734
rect 347596 234670 347648 234676
rect 347504 234660 347556 234666
rect 347504 234602 347556 234608
rect 347516 232914 347544 234602
rect 347424 232886 347544 232914
rect 347424 226234 347452 232886
rect 347412 226228 347464 226234
rect 347412 226170 347464 226176
rect 347608 224874 347636 234670
rect 347700 227322 347728 234738
rect 347688 227316 347740 227322
rect 347688 227258 347740 227264
rect 348160 226334 348188 236438
rect 348436 227186 348464 239700
rect 348804 227390 348832 239700
rect 349068 234864 349120 234870
rect 349068 234806 349120 234812
rect 348792 227384 348844 227390
rect 348792 227326 348844 227332
rect 348424 227180 348476 227186
rect 348424 227122 348476 227128
rect 348160 226306 348924 226334
rect 347596 224868 347648 224874
rect 347596 224810 347648 224816
rect 347136 224664 347188 224670
rect 347136 224606 347188 224612
rect 346504 224488 347452 224516
rect 347424 222970 347452 224488
rect 347320 222964 347372 222970
rect 347320 222906 347372 222912
rect 347412 222964 347464 222970
rect 347412 222906 347464 222912
rect 346400 221808 346452 221814
rect 346400 221750 346452 221756
rect 346492 221060 346544 221066
rect 346492 221002 346544 221008
rect 346504 217410 346532 221002
rect 347332 217410 347360 222906
rect 348148 221468 348200 221474
rect 348148 221410 348200 221416
rect 348160 217410 348188 221410
rect 348896 217410 348924 226306
rect 349080 222222 349108 234806
rect 349172 234734 349200 239700
rect 349160 234728 349212 234734
rect 349160 234670 349212 234676
rect 349448 234666 349476 239700
rect 349436 234660 349488 234666
rect 349436 234602 349488 234608
rect 349816 227662 349844 239700
rect 349896 234796 349948 234802
rect 349896 234738 349948 234744
rect 349804 227656 349856 227662
rect 349804 227598 349856 227604
rect 349908 226302 349936 234738
rect 350184 227526 350212 239700
rect 350552 234734 350580 239700
rect 350920 234802 350948 239700
rect 351092 236360 351144 236366
rect 351092 236302 351144 236308
rect 350908 234796 350960 234802
rect 350908 234738 350960 234744
rect 350264 234728 350316 234734
rect 350264 234670 350316 234676
rect 350540 234728 350592 234734
rect 350540 234670 350592 234676
rect 350172 227520 350224 227526
rect 350172 227462 350224 227468
rect 349896 226296 349948 226302
rect 349896 226238 349948 226244
rect 350276 226030 350304 234670
rect 350356 234660 350408 234666
rect 350356 234602 350408 234608
rect 350264 226024 350316 226030
rect 350264 225966 350316 225972
rect 350368 225826 350396 234602
rect 350356 225820 350408 225826
rect 350356 225762 350408 225768
rect 349068 222216 349120 222222
rect 349068 222158 349120 222164
rect 350632 221604 350684 221610
rect 350632 221546 350684 221552
rect 349804 221128 349856 221134
rect 349804 221070 349856 221076
rect 349816 217410 349844 221070
rect 350644 217410 350672 221546
rect 351104 221338 351132 236302
rect 351288 227458 351316 239700
rect 351656 227594 351684 239700
rect 352024 234666 352052 239700
rect 352314 239686 352604 239714
rect 352682 239686 352972 239714
rect 353050 239686 353248 239714
rect 352576 234818 352604 239686
rect 352944 234920 352972 239686
rect 352944 234892 353156 234920
rect 352576 234790 352972 234818
rect 352564 234728 352616 234734
rect 352564 234670 352616 234676
rect 352012 234660 352064 234666
rect 352012 234602 352064 234608
rect 351644 227588 351696 227594
rect 351644 227530 351696 227536
rect 351276 227452 351328 227458
rect 351276 227394 351328 227400
rect 352576 226098 352604 234670
rect 352656 234660 352708 234666
rect 352656 234602 352708 234608
rect 352564 226092 352616 226098
rect 352564 226034 352616 226040
rect 352668 225962 352696 234602
rect 352656 225956 352708 225962
rect 352656 225898 352708 225904
rect 352944 225622 352972 234790
rect 353024 234796 353076 234802
rect 353024 234738 353076 234744
rect 353036 225894 353064 234738
rect 353128 229090 353156 234892
rect 353116 229084 353168 229090
rect 353116 229026 353168 229032
rect 353220 228818 353248 239686
rect 353404 234802 353432 239700
rect 353392 234796 353444 234802
rect 353392 234738 353444 234744
rect 353772 234734 353800 239700
rect 353760 234728 353812 234734
rect 353760 234670 353812 234676
rect 354140 229022 354168 239700
rect 354128 229016 354180 229022
rect 354128 228958 354180 228964
rect 354508 228886 354536 239700
rect 354876 234666 354904 239700
rect 355166 239686 355364 239714
rect 354864 234660 354916 234666
rect 354864 234602 354916 234608
rect 354496 228880 354548 228886
rect 354496 228822 354548 228828
rect 353208 228812 353260 228818
rect 353208 228754 353260 228760
rect 353024 225888 353076 225894
rect 353024 225830 353076 225836
rect 352932 225616 352984 225622
rect 352932 225558 352984 225564
rect 355336 225554 355364 239686
rect 355416 234728 355468 234734
rect 355416 234670 355468 234676
rect 355428 225690 355456 234670
rect 355520 228954 355548 239700
rect 355784 234796 355836 234802
rect 355784 234738 355836 234744
rect 355692 234660 355744 234666
rect 355692 234602 355744 234608
rect 355508 228948 355560 228954
rect 355508 228890 355560 228896
rect 355416 225684 355468 225690
rect 355416 225626 355468 225632
rect 355324 225548 355376 225554
rect 355324 225490 355376 225496
rect 355704 225418 355732 234602
rect 355796 225758 355824 234738
rect 355888 228682 355916 239700
rect 356256 234802 356284 239700
rect 356428 236292 356480 236298
rect 356428 236234 356480 236240
rect 356244 234796 356296 234802
rect 356244 234738 356296 234744
rect 355876 228676 355928 228682
rect 355876 228618 355928 228624
rect 355784 225752 355836 225758
rect 355784 225694 355836 225700
rect 355692 225412 355744 225418
rect 355692 225354 355744 225360
rect 354036 221944 354088 221950
rect 354036 221886 354088 221892
rect 351460 221672 351512 221678
rect 351460 221614 351512 221620
rect 351092 221332 351144 221338
rect 351092 221274 351144 221280
rect 351472 217410 351500 221614
rect 352380 221332 352432 221338
rect 352380 221274 352432 221280
rect 352392 217410 352420 221274
rect 353300 221196 353352 221202
rect 353300 221138 353352 221144
rect 353312 217410 353340 221138
rect 354048 217410 354076 221886
rect 354864 221740 354916 221746
rect 354864 221682 354916 221688
rect 354876 217410 354904 221682
rect 356440 217410 356468 236234
rect 356624 234734 356652 239700
rect 356612 234728 356664 234734
rect 356612 234670 356664 234676
rect 356992 228614 357020 239700
rect 357360 228750 357388 239700
rect 357728 234666 357756 239700
rect 358018 239686 358216 239714
rect 358084 234728 358136 234734
rect 358084 234670 358136 234676
rect 357716 234660 357768 234666
rect 357716 234602 357768 234608
rect 357348 228744 357400 228750
rect 357348 228686 357400 228692
rect 356980 228608 357032 228614
rect 356980 228550 357032 228556
rect 358096 225350 358124 234670
rect 358084 225344 358136 225350
rect 358084 225286 358136 225292
rect 358188 225146 358216 239686
rect 358372 228546 358400 239700
rect 358544 234796 358596 234802
rect 358544 234738 358596 234744
rect 358452 234660 358504 234666
rect 358452 234602 358504 234608
rect 358360 228540 358412 228546
rect 358360 228482 358412 228488
rect 358464 225214 358492 234602
rect 358556 225486 358584 234738
rect 358740 228410 358768 239700
rect 359108 234802 359136 239700
rect 359188 236224 359240 236230
rect 359188 236166 359240 236172
rect 359096 234796 359148 234802
rect 359096 234738 359148 234744
rect 358728 228404 358780 228410
rect 358728 228346 358780 228352
rect 358544 225480 358596 225486
rect 358544 225422 358596 225428
rect 358452 225208 358504 225214
rect 358452 225150 358504 225156
rect 358176 225140 358228 225146
rect 358176 225082 358228 225088
rect 358268 222080 358320 222086
rect 358268 222022 358320 222028
rect 356520 222012 356572 222018
rect 356520 221954 356572 221960
rect 343100 217382 343436 217410
rect 343928 217382 344264 217410
rect 345032 217382 345092 217410
rect 345492 217382 345920 217410
rect 346504 217382 346840 217410
rect 347332 217382 347668 217410
rect 348160 217382 348496 217410
rect 348896 217382 349324 217410
rect 349816 217382 350152 217410
rect 350644 217382 350980 217410
rect 351472 217382 351808 217410
rect 352392 217382 352728 217410
rect 353312 217382 353556 217410
rect 354048 217382 354384 217410
rect 354876 217382 355212 217410
rect 356040 217382 356468 217410
rect 356532 217410 356560 221954
rect 357348 221876 357400 221882
rect 357348 221818 357400 221824
rect 357360 217410 357388 221818
rect 358280 217410 358308 222022
rect 359200 217410 359228 236166
rect 359476 234734 359504 239700
rect 359464 234728 359516 234734
rect 359464 234670 359516 234676
rect 359844 228478 359872 239700
rect 359832 228472 359884 228478
rect 359832 228414 359884 228420
rect 360212 228342 360240 239700
rect 360580 234666 360608 239700
rect 360870 239686 360976 239714
rect 361238 239686 361528 239714
rect 360568 234660 360620 234666
rect 360568 234602 360620 234608
rect 360200 228336 360252 228342
rect 360200 228278 360252 228284
rect 360948 226137 360976 239686
rect 361212 234796 361264 234802
rect 361212 234738 361264 234744
rect 360934 226128 360990 226137
rect 360934 226063 360990 226072
rect 361224 225282 361252 234738
rect 361396 234728 361448 234734
rect 361396 234670 361448 234676
rect 361304 234660 361356 234666
rect 361304 234602 361356 234608
rect 361212 225276 361264 225282
rect 361212 225218 361264 225224
rect 361316 224942 361344 234602
rect 361408 225078 361436 234670
rect 361500 228274 361528 239686
rect 361488 228268 361540 228274
rect 361488 228210 361540 228216
rect 361592 228206 361620 239700
rect 361960 234666 361988 239700
rect 362328 234734 362356 239700
rect 362316 234728 362368 234734
rect 362316 234670 362368 234676
rect 361948 234660 362000 234666
rect 361948 234602 362000 234608
rect 361580 228200 361632 228206
rect 361580 228142 361632 228148
rect 362696 228138 362724 239700
rect 363064 231742 363092 239700
rect 363446 239686 363644 239714
rect 363722 239686 364012 239714
rect 364090 239686 364288 239714
rect 363512 234660 363564 234666
rect 363512 234602 363564 234608
rect 363052 231736 363104 231742
rect 363052 231678 363104 231684
rect 362684 228132 362736 228138
rect 362684 228074 362736 228080
rect 361396 225072 361448 225078
rect 361396 225014 361448 225020
rect 363524 225010 363552 234602
rect 363616 233050 363644 239686
rect 363616 233022 363736 233050
rect 363708 225729 363736 233022
rect 363984 227934 364012 239686
rect 364064 234728 364116 234734
rect 364064 234670 364116 234676
rect 363972 227928 364024 227934
rect 363972 227870 364024 227876
rect 364076 226001 364104 234670
rect 364260 228002 364288 239686
rect 364444 231674 364472 239700
rect 364812 234666 364840 239700
rect 364800 234660 364852 234666
rect 364800 234602 364852 234608
rect 364432 231668 364484 231674
rect 364432 231610 364484 231616
rect 364248 227996 364300 228002
rect 364248 227938 364300 227944
rect 365180 227798 365208 239700
rect 365548 228070 365576 239700
rect 365916 231538 365944 239700
rect 366298 239686 366404 239714
rect 365904 231532 365956 231538
rect 365904 231474 365956 231480
rect 365536 228064 365588 228070
rect 365536 228006 365588 228012
rect 365168 227792 365220 227798
rect 365168 227734 365220 227740
rect 364062 225992 364118 226001
rect 364062 225927 364118 225936
rect 363694 225720 363750 225729
rect 363694 225655 363750 225664
rect 366376 225593 366404 239686
rect 366560 228857 366588 239700
rect 366546 228848 366602 228857
rect 366546 228783 366602 228792
rect 366928 227730 366956 239700
rect 367008 234660 367060 234666
rect 367008 234602 367060 234608
rect 366916 227724 366968 227730
rect 366916 227666 366968 227672
rect 367020 225865 367048 234602
rect 367296 231606 367324 239700
rect 367664 234666 367692 239700
rect 367652 234660 367704 234666
rect 367652 234602 367704 234608
rect 367284 231600 367336 231606
rect 367284 231542 367336 231548
rect 368032 228721 368060 239700
rect 368018 228712 368074 228721
rect 368018 228647 368074 228656
rect 368400 227866 368428 239700
rect 368768 231402 368796 239700
rect 369150 239686 369256 239714
rect 369124 234660 369176 234666
rect 369124 234602 369176 234608
rect 368756 231396 368808 231402
rect 368756 231338 368808 231344
rect 368388 227860 368440 227866
rect 368388 227802 368440 227808
rect 367006 225856 367062 225865
rect 367006 225791 367062 225800
rect 366362 225584 366418 225593
rect 366362 225519 366418 225528
rect 369136 225457 369164 234602
rect 369122 225448 369178 225457
rect 369122 225383 369178 225392
rect 369228 225185 369256 239686
rect 369412 228041 369440 239700
rect 369780 228449 369808 239700
rect 370148 231470 370176 239700
rect 370516 234666 370544 239700
rect 370504 234660 370556 234666
rect 370504 234602 370556 234608
rect 370136 231464 370188 231470
rect 370136 231406 370188 231412
rect 369766 228440 369822 228449
rect 369766 228375 369822 228384
rect 370884 228177 370912 239700
rect 371252 228585 371280 239700
rect 371620 231334 371648 239700
rect 372002 239686 372108 239714
rect 371976 234660 372028 234666
rect 371976 234602 372028 234608
rect 371608 231328 371660 231334
rect 371608 231270 371660 231276
rect 371238 228576 371294 228585
rect 371238 228511 371294 228520
rect 370870 228168 370926 228177
rect 370870 228103 370926 228112
rect 369398 228032 369454 228041
rect 369398 227967 369454 227976
rect 371988 225321 372016 234602
rect 371974 225312 372030 225321
rect 371974 225247 372030 225256
rect 369214 225176 369270 225185
rect 369214 225111 369270 225120
rect 372080 225049 372108 239686
rect 372264 227633 372292 239700
rect 372632 228313 372660 239700
rect 373000 231266 373028 239700
rect 373368 234666 373396 239700
rect 373356 234660 373408 234666
rect 373356 234602 373408 234608
rect 372988 231260 373040 231266
rect 372988 231202 373040 231208
rect 372618 228304 372674 228313
rect 372618 228239 372674 228248
rect 373736 227769 373764 239700
rect 374104 227905 374132 239700
rect 374472 231198 374500 239700
rect 374564 239686 374854 239714
rect 374932 239686 375130 239714
rect 374460 231192 374512 231198
rect 374460 231134 374512 231140
rect 374564 231130 374592 239686
rect 374932 234784 374960 239686
rect 374656 234756 374960 234784
rect 374552 231124 374604 231130
rect 374552 231066 374604 231072
rect 374090 227896 374146 227905
rect 374090 227831 374146 227840
rect 373722 227760 373778 227769
rect 373722 227695 373778 227704
rect 372250 227624 372306 227633
rect 372250 227559 372306 227568
rect 372066 225040 372122 225049
rect 363512 225004 363564 225010
rect 372066 224975 372122 224984
rect 363512 224946 363564 224952
rect 361304 224936 361356 224942
rect 361304 224878 361356 224884
rect 361764 223576 361816 223582
rect 361764 223518 361816 223524
rect 360752 222148 360804 222154
rect 360752 222090 360804 222096
rect 359924 221264 359976 221270
rect 359924 221206 359976 221212
rect 359936 217410 359964 221206
rect 360764 217410 360792 222090
rect 361776 217410 361804 223518
rect 362408 223508 362460 223514
rect 362408 223450 362460 223456
rect 362420 217410 362448 223450
rect 374656 223417 374684 234756
rect 375484 234734 375512 239700
rect 375748 237380 375800 237386
rect 375748 237322 375800 237328
rect 375472 234728 375524 234734
rect 375472 234670 375524 234676
rect 374736 234660 374788 234666
rect 374736 234602 374788 234608
rect 374748 224913 374776 234602
rect 375760 226334 375788 237322
rect 375852 237153 375880 239700
rect 375838 237144 375894 237153
rect 375838 237079 375894 237088
rect 376220 231062 376248 239700
rect 376588 235006 376616 239700
rect 376576 235000 376628 235006
rect 376576 234942 376628 234948
rect 376956 234666 376984 239700
rect 377338 239686 377628 239714
rect 376944 234660 376996 234666
rect 376944 234602 376996 234608
rect 376208 231056 376260 231062
rect 376208 230998 376260 231004
rect 375760 226306 375880 226334
rect 374734 224904 374790 224913
rect 374734 224839 374790 224848
rect 374642 223408 374698 223417
rect 369124 223372 369176 223378
rect 374642 223343 374698 223352
rect 369124 223314 369176 223320
rect 368296 223304 368348 223310
rect 368296 223246 368348 223252
rect 365812 223236 365864 223242
rect 365812 223178 365864 223184
rect 364984 223168 365036 223174
rect 364984 223110 365036 223116
rect 364340 223032 364392 223038
rect 364340 222974 364392 222980
rect 363236 220992 363288 220998
rect 363236 220934 363288 220940
rect 363248 217410 363276 220934
rect 364352 217410 364380 222974
rect 364996 217410 365024 223110
rect 365824 217410 365852 223178
rect 367468 222828 367520 222834
rect 367468 222770 367520 222776
rect 366640 221400 366692 221406
rect 366640 221342 366692 221348
rect 366652 217410 366680 221342
rect 367480 217410 367508 222770
rect 368308 217410 368336 223246
rect 369136 217410 369164 223314
rect 371700 223100 371752 223106
rect 371700 223042 371752 223048
rect 370044 222896 370096 222902
rect 370044 222838 370096 222844
rect 370056 217410 370084 222838
rect 370872 222760 370924 222766
rect 370872 222702 370924 222708
rect 370884 217410 370912 222702
rect 371712 217410 371740 223042
rect 374182 222864 374238 222873
rect 374182 222799 374238 222808
rect 372620 222624 372672 222630
rect 372620 222566 372672 222572
rect 372632 217410 372660 222566
rect 373356 221536 373408 221542
rect 373356 221478 373408 221484
rect 373368 217410 373396 221478
rect 374196 217410 374224 222799
rect 375378 222728 375434 222737
rect 375378 222663 375434 222672
rect 375392 217410 375420 222663
rect 356532 217382 356868 217410
rect 357360 217382 357696 217410
rect 358280 217382 358616 217410
rect 359200 217382 359444 217410
rect 359936 217382 360272 217410
rect 360764 217382 361100 217410
rect 361776 217382 361928 217410
rect 362420 217382 362756 217410
rect 363248 217382 363584 217410
rect 364352 217382 364504 217410
rect 364996 217382 365332 217410
rect 365824 217382 366160 217410
rect 366652 217382 366988 217410
rect 367480 217382 367816 217410
rect 368308 217382 368644 217410
rect 369136 217382 369472 217410
rect 370056 217382 370392 217410
rect 370884 217382 371220 217410
rect 371712 217382 372048 217410
rect 372632 217382 372876 217410
rect 373368 217382 373704 217410
rect 374196 217382 374532 217410
rect 375360 217382 375420 217410
rect 375852 217410 375880 226306
rect 377600 223281 377628 239686
rect 377692 233510 377720 239700
rect 377968 236162 377996 239700
rect 378336 237017 378364 239700
rect 378322 237008 378378 237017
rect 378322 236943 378378 236952
rect 378704 236881 378732 239700
rect 378690 236872 378746 236881
rect 378690 236807 378746 236816
rect 377956 236156 378008 236162
rect 377956 236098 378008 236104
rect 378508 236088 378560 236094
rect 378508 236030 378560 236036
rect 377956 234660 378008 234666
rect 377956 234602 378008 234608
rect 377680 233504 377732 233510
rect 377680 233446 377732 233452
rect 377586 223272 377642 223281
rect 377586 223207 377642 223216
rect 377968 223145 377996 234602
rect 378520 226334 378548 236030
rect 379072 235142 379100 239700
rect 379440 236230 379468 239700
rect 379428 236224 379480 236230
rect 379428 236166 379480 236172
rect 379060 235136 379112 235142
rect 379060 235078 379112 235084
rect 379428 234728 379480 234734
rect 379428 234670 379480 234676
rect 378520 226306 379192 226334
rect 376758 223136 376814 223145
rect 376758 223071 376814 223080
rect 377954 223136 378010 223145
rect 377954 223071 378010 223080
rect 376772 217410 376800 223071
rect 377586 223000 377642 223009
rect 377586 222935 377642 222944
rect 377600 217410 377628 222935
rect 378416 222692 378468 222698
rect 378416 222634 378468 222640
rect 378428 217410 378456 222634
rect 379164 217410 379192 226306
rect 379440 221474 379468 234670
rect 379808 234666 379836 239700
rect 380190 239686 380480 239714
rect 380558 239686 380756 239714
rect 379796 234660 379848 234666
rect 379796 234602 379848 234608
rect 380452 222873 380480 239686
rect 380624 234660 380676 234666
rect 380624 234602 380676 234608
rect 380636 229514 380664 234602
rect 380728 229650 380756 239686
rect 380820 235074 380848 239700
rect 381188 236745 381216 239700
rect 381174 236736 381230 236745
rect 381174 236671 381230 236680
rect 381556 236473 381584 239700
rect 381542 236464 381598 236473
rect 381542 236399 381598 236408
rect 381924 235210 381952 239700
rect 381912 235204 381964 235210
rect 381912 235146 381964 235152
rect 380808 235068 380860 235074
rect 380808 235010 380860 235016
rect 382292 234666 382320 239700
rect 382674 239686 382964 239714
rect 383042 239686 383332 239714
rect 382280 234660 382332 234666
rect 382280 234602 382332 234608
rect 380728 229622 380848 229650
rect 380636 229486 380756 229514
rect 380728 223009 380756 229486
rect 380714 223000 380770 223009
rect 380714 222935 380770 222944
rect 380438 222864 380494 222873
rect 380438 222799 380494 222808
rect 380072 221808 380124 221814
rect 380072 221750 380124 221756
rect 379428 221468 379480 221474
rect 379428 221410 379480 221416
rect 380084 217410 380112 221750
rect 380820 221610 380848 229622
rect 382648 223916 382700 223922
rect 382648 223858 382700 223864
rect 381082 222592 381138 222601
rect 381082 222527 381138 222536
rect 381820 222556 381872 222562
rect 380808 221604 380860 221610
rect 380808 221546 380860 221552
rect 381096 217410 381124 222527
rect 381820 222498 381872 222504
rect 381832 217410 381860 222498
rect 382660 217410 382688 223858
rect 382936 222601 382964 239686
rect 383304 233050 383332 239686
rect 383396 235278 383424 239700
rect 383672 236609 383700 239700
rect 383658 236600 383714 236609
rect 383658 236535 383714 236544
rect 384040 235346 384068 239700
rect 384028 235340 384080 235346
rect 384028 235282 384080 235288
rect 383384 235272 383436 235278
rect 383384 235214 383436 235220
rect 384408 234802 384436 239700
rect 384396 234796 384448 234802
rect 384396 234738 384448 234744
rect 384776 234734 384804 239700
rect 384764 234728 384816 234734
rect 384764 234670 384816 234676
rect 385144 234666 385172 239700
rect 385512 235414 385540 239700
rect 385880 236337 385908 239700
rect 385866 236328 385922 236337
rect 385866 236263 385922 236272
rect 386248 235618 386276 239700
rect 386236 235612 386288 235618
rect 386236 235554 386288 235560
rect 385500 235408 385552 235414
rect 385500 235350 385552 235356
rect 386524 234870 386552 239700
rect 386512 234864 386564 234870
rect 386512 234806 386564 234812
rect 386236 234728 386288 234734
rect 386236 234670 386288 234676
rect 384948 234660 385000 234666
rect 384948 234602 385000 234608
rect 385132 234660 385184 234666
rect 385132 234602 385184 234608
rect 383304 233022 383608 233050
rect 382922 222592 382978 222601
rect 382922 222527 382978 222536
rect 383580 221882 383608 233022
rect 383660 223440 383712 223446
rect 383660 223382 383712 223388
rect 383568 221876 383620 221882
rect 383568 221818 383620 221824
rect 383672 217410 383700 223382
rect 384302 222456 384358 222465
rect 384302 222391 384358 222400
rect 384316 217410 384344 222391
rect 384960 221542 384988 234602
rect 385960 223984 386012 223990
rect 385960 223926 386012 223932
rect 385132 222488 385184 222494
rect 385132 222430 385184 222436
rect 384948 221536 385000 221542
rect 384948 221478 385000 221484
rect 385144 217410 385172 222430
rect 385972 217410 386000 223926
rect 386248 222737 386276 234670
rect 386892 234666 386920 239700
rect 387260 234734 387288 239700
rect 387628 236298 387656 239700
rect 387616 236292 387668 236298
rect 387616 236234 387668 236240
rect 387996 236201 388024 239700
rect 387982 236192 388038 236201
rect 387616 236156 387668 236162
rect 387982 236127 388038 236136
rect 387616 236098 387668 236104
rect 387248 234728 387300 234734
rect 387248 234670 387300 234676
rect 386328 234660 386380 234666
rect 386328 234602 386380 234608
rect 386880 234660 386932 234666
rect 386880 234602 386932 234608
rect 386234 222728 386290 222737
rect 386234 222663 386290 222672
rect 386340 222018 386368 234602
rect 386788 222964 386840 222970
rect 386788 222906 386840 222912
rect 386328 222012 386380 222018
rect 386328 221954 386380 221960
rect 386800 217410 386828 222906
rect 387628 221406 387656 236098
rect 387800 234796 387852 234802
rect 387800 234738 387852 234744
rect 387706 222320 387762 222329
rect 387706 222255 387762 222264
rect 387616 221400 387668 221406
rect 387616 221342 387668 221348
rect 387720 217410 387748 222255
rect 387812 221678 387840 234738
rect 388364 230314 388392 239700
rect 388732 235482 388760 239700
rect 389100 236065 389128 239700
rect 389086 236056 389142 236065
rect 389086 235991 389142 236000
rect 388720 235476 388772 235482
rect 388720 235418 388772 235424
rect 389088 234728 389140 234734
rect 389088 234670 389140 234676
rect 388996 234660 389048 234666
rect 388996 234602 389048 234608
rect 388352 230308 388404 230314
rect 388352 230250 388404 230256
rect 389008 222465 389036 234602
rect 388994 222456 389050 222465
rect 388536 222420 388588 222426
rect 388994 222391 389050 222400
rect 388536 222362 388588 222368
rect 387800 221672 387852 221678
rect 387800 221614 387852 221620
rect 388548 217410 388576 222362
rect 389100 222086 389128 234670
rect 389376 230994 389404 239700
rect 389744 233782 389772 239700
rect 390112 234666 390140 239700
rect 390376 236224 390428 236230
rect 390376 236166 390428 236172
rect 390100 234660 390152 234666
rect 390100 234602 390152 234608
rect 389732 233776 389784 233782
rect 389732 233718 389784 233724
rect 389364 230988 389416 230994
rect 389364 230930 389416 230936
rect 389364 230716 389416 230722
rect 389364 230658 389416 230664
rect 389088 222080 389140 222086
rect 389088 222022 389140 222028
rect 389376 217410 389404 230658
rect 390190 222048 390246 222057
rect 390190 221983 390246 221992
rect 390204 217410 390232 221983
rect 390388 221338 390416 236166
rect 390480 230926 390508 239700
rect 390848 236162 390876 239700
rect 390836 236156 390888 236162
rect 390836 236098 390888 236104
rect 391216 235929 391244 239700
rect 391202 235920 391258 235929
rect 391202 235855 391258 235864
rect 390560 234864 390612 234870
rect 390560 234806 390612 234812
rect 390468 230920 390520 230926
rect 390468 230862 390520 230868
rect 390572 221950 390600 234806
rect 391584 230858 391612 239700
rect 391952 234666 391980 239700
rect 391848 234660 391900 234666
rect 391848 234602 391900 234608
rect 391940 234660 391992 234666
rect 391940 234602 391992 234608
rect 391572 230852 391624 230858
rect 391572 230794 391624 230800
rect 391020 224052 391072 224058
rect 391020 223994 391072 224000
rect 390560 221944 390612 221950
rect 390560 221886 390612 221892
rect 390376 221332 390428 221338
rect 390376 221274 390428 221280
rect 391032 217410 391060 223994
rect 391860 222329 391888 234602
rect 391846 222320 391902 222329
rect 391846 222255 391902 222264
rect 391940 222284 391992 222290
rect 391940 222226 391992 222232
rect 391952 217410 391980 222226
rect 392228 220930 392256 239700
rect 392596 230722 392624 239700
rect 392964 235754 392992 239700
rect 393332 235890 393360 239700
rect 393320 235884 393372 235890
rect 393320 235826 393372 235832
rect 392952 235748 393004 235754
rect 392952 235690 393004 235696
rect 393700 233442 393728 239700
rect 393780 235612 393832 235618
rect 393964 235612 394016 235618
rect 393832 235572 393964 235600
rect 393780 235554 393832 235560
rect 393964 235554 394016 235560
rect 394068 235550 394096 239700
rect 394450 239686 394556 239714
rect 394056 235544 394108 235550
rect 394056 235486 394108 235492
rect 393688 233436 393740 233442
rect 393688 233378 393740 233384
rect 392584 230716 392636 230722
rect 392584 230658 392636 230664
rect 392676 230648 392728 230654
rect 392676 230590 392728 230596
rect 392216 220924 392268 220930
rect 392216 220866 392268 220872
rect 392688 217410 392716 230590
rect 394528 223310 394556 239686
rect 394804 230654 394832 239700
rect 395080 235822 395108 239700
rect 395448 237386 395476 239700
rect 395436 237380 395488 237386
rect 395436 237322 395488 237328
rect 395160 236020 395212 236026
rect 395160 235962 395212 235968
rect 395068 235816 395120 235822
rect 395068 235758 395120 235764
rect 394792 230648 394844 230654
rect 394792 230590 394844 230596
rect 394700 224256 394752 224262
rect 394700 224198 394752 224204
rect 394516 223304 394568 223310
rect 394516 223246 394568 223252
rect 393596 222352 393648 222358
rect 393596 222294 393648 222300
rect 393608 217410 393636 222294
rect 394712 217410 394740 224198
rect 395172 217410 395200 235962
rect 395816 230586 395844 239700
rect 396184 236366 396212 239700
rect 396566 239686 396856 239714
rect 396172 236360 396224 236366
rect 396172 236302 396224 236308
rect 395712 230580 395764 230586
rect 395712 230522 395764 230528
rect 395804 230580 395856 230586
rect 395804 230522 395856 230528
rect 395724 218054 395752 230522
rect 396828 220998 396856 239686
rect 396920 233374 396948 239700
rect 397288 237318 397316 239700
rect 397276 237312 397328 237318
rect 397276 237254 397328 237260
rect 397656 235958 397684 239700
rect 397644 235952 397696 235958
rect 397644 235894 397696 235900
rect 396908 233368 396960 233374
rect 396908 233310 396960 233316
rect 397932 233306 397960 239700
rect 398300 234734 398328 239700
rect 398288 234728 398340 234734
rect 398288 234670 398340 234676
rect 397920 233300 397972 233306
rect 397920 233242 397972 233248
rect 398564 226704 398616 226710
rect 398564 226646 398616 226652
rect 397736 224188 397788 224194
rect 397736 224130 397788 224136
rect 396906 223544 396962 223553
rect 396906 223479 396962 223488
rect 396816 220992 396868 220998
rect 396816 220934 396868 220940
rect 395724 218026 396120 218054
rect 396092 217410 396120 218026
rect 396920 217410 396948 223479
rect 397748 217410 397776 224130
rect 398576 217410 398604 226646
rect 398668 223242 398696 239700
rect 399036 236978 399064 239700
rect 399404 237250 399432 239700
rect 399786 239686 400076 239714
rect 399392 237244 399444 237250
rect 399392 237186 399444 237192
rect 399024 236972 399076 236978
rect 399024 236914 399076 236920
rect 399300 236360 399352 236366
rect 399300 236302 399352 236308
rect 398656 223236 398708 223242
rect 398656 223178 398708 223184
rect 399312 221066 399340 236302
rect 399484 230376 399536 230382
rect 399484 230318 399536 230324
rect 399300 221060 399352 221066
rect 399300 221002 399352 221008
rect 399496 217410 399524 230318
rect 400048 223106 400076 239686
rect 400140 233238 400168 239700
rect 400508 237182 400536 239700
rect 400496 237176 400548 237182
rect 400496 237118 400548 237124
rect 400784 236230 400812 239700
rect 401152 237114 401180 239700
rect 401140 237108 401192 237114
rect 401140 237050 401192 237056
rect 401520 236434 401548 239700
rect 401508 236428 401560 236434
rect 401508 236370 401560 236376
rect 401508 236292 401560 236298
rect 401508 236234 401560 236240
rect 400772 236224 400824 236230
rect 400772 236166 400824 236172
rect 401520 235550 401548 236234
rect 401600 236156 401652 236162
rect 401600 236098 401652 236104
rect 401612 235686 401640 236098
rect 401600 235680 401652 235686
rect 401600 235622 401652 235628
rect 401416 235544 401468 235550
rect 401416 235486 401468 235492
rect 401508 235544 401560 235550
rect 401508 235486 401560 235492
rect 401324 233776 401376 233782
rect 401324 233718 401376 233724
rect 400128 233232 400180 233238
rect 400128 233174 400180 233180
rect 401140 224120 401192 224126
rect 401140 224062 401192 224068
rect 400036 223100 400088 223106
rect 400036 223042 400088 223048
rect 400402 222184 400458 222193
rect 400402 222119 400458 222128
rect 400416 217410 400444 222119
rect 401152 217410 401180 224062
rect 401336 221746 401364 233718
rect 401428 222154 401456 235486
rect 401600 230988 401652 230994
rect 401600 230930 401652 230936
rect 401612 230314 401640 230930
rect 401600 230308 401652 230314
rect 401600 230250 401652 230256
rect 401888 223038 401916 239700
rect 402270 239686 402560 239714
rect 401968 226772 402020 226778
rect 401968 226714 402020 226720
rect 401876 223032 401928 223038
rect 401876 222974 401928 222980
rect 401416 222148 401468 222154
rect 401416 222090 401468 222096
rect 401324 221740 401376 221746
rect 401324 221682 401376 221688
rect 401980 217410 402008 226714
rect 402532 222970 402560 239686
rect 402624 234938 402652 239700
rect 402992 236910 403020 239700
rect 402980 236904 403032 236910
rect 402980 236846 403032 236852
rect 403360 236842 403388 239700
rect 403348 236836 403400 236842
rect 403348 236778 403400 236784
rect 402612 234932 402664 234938
rect 402612 234874 402664 234880
rect 403636 234666 403664 239700
rect 403808 234728 403860 234734
rect 403808 234670 403860 234676
rect 403072 234660 403124 234666
rect 403072 234602 403124 234608
rect 403624 234660 403676 234666
rect 403624 234602 403676 234608
rect 402980 224460 403032 224466
rect 402980 224402 403032 224408
rect 402520 222964 402572 222970
rect 402520 222906 402572 222912
rect 402992 217410 403020 224402
rect 403084 221814 403112 234602
rect 403624 231804 403676 231810
rect 403624 231746 403676 231752
rect 403072 221808 403124 221814
rect 403072 221750 403124 221756
rect 403636 217410 403664 231746
rect 403820 223446 403848 234670
rect 403808 223440 403860 223446
rect 403808 223382 403860 223388
rect 404004 222698 404032 239700
rect 404372 222766 404400 239700
rect 404740 236706 404768 239700
rect 405108 237046 405136 239700
rect 405096 237040 405148 237046
rect 405096 236982 405148 236988
rect 405476 236774 405504 239700
rect 405464 236768 405516 236774
rect 405464 236710 405516 236716
rect 404728 236700 404780 236706
rect 404728 236642 404780 236648
rect 405740 226840 405792 226846
rect 405740 226782 405792 226788
rect 404452 224392 404504 224398
rect 404452 224334 404504 224340
rect 404360 222760 404412 222766
rect 404360 222702 404412 222708
rect 403992 222692 404044 222698
rect 403992 222634 404044 222640
rect 404464 217410 404492 224334
rect 405752 217410 405780 226782
rect 405844 222834 405872 239700
rect 406212 237374 406240 239700
rect 406212 237346 406332 237374
rect 406200 224528 406252 224534
rect 406200 224470 406252 224476
rect 405832 222828 405884 222834
rect 405832 222770 405884 222776
rect 375852 217382 376280 217410
rect 376772 217382 377108 217410
rect 377600 217382 377936 217410
rect 378428 217382 378764 217410
rect 379164 217382 379592 217410
rect 380084 217382 380420 217410
rect 381096 217382 381248 217410
rect 381832 217382 382168 217410
rect 382660 217382 382996 217410
rect 383672 217382 383824 217410
rect 384316 217382 384652 217410
rect 385144 217382 385480 217410
rect 385972 217382 386308 217410
rect 386800 217382 387136 217410
rect 387720 217382 388056 217410
rect 388548 217382 388884 217410
rect 389376 217382 389712 217410
rect 390204 217382 390540 217410
rect 391032 217382 391368 217410
rect 391952 217382 392196 217410
rect 392688 217382 393024 217410
rect 393608 217382 393944 217410
rect 394712 217382 394772 217410
rect 395172 217382 395600 217410
rect 396092 217382 396428 217410
rect 396920 217382 397256 217410
rect 397748 217382 398084 217410
rect 398576 217382 398912 217410
rect 399496 217382 399832 217410
rect 400416 217382 400660 217410
rect 401152 217382 401488 217410
rect 401980 217382 402316 217410
rect 402992 217382 403144 217410
rect 403636 217382 403972 217410
rect 404464 217382 404800 217410
rect 405720 217382 405780 217410
rect 406212 217410 406240 224470
rect 406304 222630 406332 237346
rect 406384 236428 406436 236434
rect 406384 236370 406436 236376
rect 406396 223174 406424 236370
rect 406384 223168 406436 223174
rect 406384 223110 406436 223116
rect 406292 222624 406344 222630
rect 406292 222566 406344 222572
rect 406488 222562 406516 239700
rect 406856 236638 406884 239700
rect 406844 236632 406896 236638
rect 406844 236574 406896 236580
rect 407224 236570 407252 239700
rect 407212 236564 407264 236570
rect 407212 236506 407264 236512
rect 407592 236502 407620 239700
rect 407974 239686 408172 239714
rect 407580 236496 407632 236502
rect 407580 236438 407632 236444
rect 407396 234660 407448 234666
rect 407396 234602 407448 234608
rect 407408 222902 407436 234602
rect 407856 224324 407908 224330
rect 407856 224266 407908 224272
rect 407396 222896 407448 222902
rect 407396 222838 407448 222844
rect 406476 222556 406528 222562
rect 406476 222498 406528 222504
rect 407028 222216 407080 222222
rect 407028 222158 407080 222164
rect 407040 217410 407068 222158
rect 407868 217410 407896 224266
rect 408144 222426 408172 239686
rect 408236 239686 408342 239714
rect 408132 222420 408184 222426
rect 408132 222362 408184 222368
rect 408236 222358 408264 239686
rect 408696 237374 408724 239700
rect 408696 237346 408816 237374
rect 408684 226908 408736 226914
rect 408684 226850 408736 226856
rect 408224 222352 408276 222358
rect 408224 222294 408276 222300
rect 408696 217410 408724 226850
rect 408788 222494 408816 237346
rect 409064 236434 409092 239700
rect 409052 236428 409104 236434
rect 409052 236370 409104 236376
rect 409340 236366 409368 239700
rect 409328 236360 409380 236366
rect 409328 236302 409380 236308
rect 409512 224596 409564 224602
rect 409512 224538 409564 224544
rect 408776 222488 408828 222494
rect 408776 222430 408828 222436
rect 409524 217410 409552 224538
rect 409708 222222 409736 239700
rect 410076 236162 410104 239700
rect 410064 236156 410116 236162
rect 410064 236098 410116 236104
rect 410444 236094 410472 239700
rect 410432 236088 410484 236094
rect 410432 236030 410484 236036
rect 410812 236026 410840 239700
rect 410800 236020 410852 236026
rect 410800 235962 410852 235968
rect 410340 227044 410392 227050
rect 410340 226986 410392 226992
rect 409696 222216 409748 222222
rect 409696 222158 409748 222164
rect 410352 217410 410380 226986
rect 411180 222193 411208 239700
rect 411548 234734 411576 239700
rect 411536 234728 411588 234734
rect 411536 234670 411588 234676
rect 411916 234666 411944 239700
rect 413296 237102 413600 237130
rect 413296 236230 413324 237102
rect 413572 237046 413600 237102
rect 413468 237040 413520 237046
rect 413468 236982 413520 236988
rect 413560 237040 413612 237046
rect 413560 236982 413612 236988
rect 413480 236570 413508 236982
rect 413652 236768 413704 236774
rect 413652 236710 413704 236716
rect 413744 236768 413796 236774
rect 413744 236710 413796 236716
rect 413376 236564 413428 236570
rect 413376 236506 413428 236512
rect 413468 236564 413520 236570
rect 413468 236506 413520 236512
rect 413388 236298 413416 236506
rect 413664 236502 413692 236710
rect 413560 236496 413612 236502
rect 413560 236438 413612 236444
rect 413652 236496 413704 236502
rect 413652 236438 413704 236444
rect 413376 236292 413428 236298
rect 413376 236234 413428 236240
rect 413572 236230 413600 236438
rect 413284 236224 413336 236230
rect 413284 236166 413336 236172
rect 413560 236224 413612 236230
rect 413560 236166 413612 236172
rect 413756 234938 413784 236710
rect 413744 234932 413796 234938
rect 413744 234874 413796 234880
rect 413836 234728 413888 234734
rect 413836 234670 413888 234676
rect 411904 234660 411956 234666
rect 411904 234602 411956 234608
rect 412088 226976 412140 226982
rect 412088 226918 412140 226924
rect 411260 224800 411312 224806
rect 411260 224742 411312 224748
rect 411166 222184 411222 222193
rect 411166 222119 411222 222128
rect 411272 217410 411300 224742
rect 412100 217410 412128 226918
rect 412916 224732 412968 224738
rect 412916 224674 412968 224680
rect 412928 217410 412956 224674
rect 413848 222290 413876 234670
rect 413928 234660 413980 234666
rect 413928 234602 413980 234608
rect 413836 222284 413888 222290
rect 413836 222226 413888 222232
rect 413940 221270 413968 234602
rect 417148 227316 417200 227322
rect 417148 227258 417200 227264
rect 414020 227248 414072 227254
rect 414020 227190 414072 227196
rect 413928 221264 413980 221270
rect 413928 221206 413980 221212
rect 414032 217410 414060 227190
rect 415400 227112 415452 227118
rect 415400 227054 415452 227060
rect 414572 224664 414624 224670
rect 414572 224606 414624 224612
rect 414584 217410 414612 224606
rect 415412 217410 415440 227054
rect 416228 224868 416280 224874
rect 416228 224810 416280 224816
rect 416240 217410 416268 224810
rect 417160 217410 417188 227258
rect 406212 217382 406548 217410
rect 407040 217382 407376 217410
rect 407868 217382 408204 217410
rect 408696 217382 409032 217410
rect 409524 217382 409860 217410
rect 410352 217382 410688 217410
rect 411272 217382 411608 217410
rect 412100 217382 412436 217410
rect 412928 217382 413264 217410
rect 414032 217382 414092 217410
rect 414584 217382 414920 217410
rect 415412 217382 415748 217410
rect 416240 217382 416576 217410
rect 417160 217382 417496 217410
rect 418080 216714 418108 248231
rect 418434 245984 418490 245993
rect 418434 245919 418490 245928
rect 418158 243536 418214 243545
rect 418158 243471 418214 243480
rect 59452 216708 59504 216714
rect 59452 216650 59504 216656
rect 418068 216708 418120 216714
rect 418068 216650 418120 216656
rect 418172 216646 418200 243471
rect 418252 226228 418304 226234
rect 418252 226170 418304 226176
rect 418264 217410 418292 226170
rect 418264 217382 418324 217410
rect 418448 216782 418476 245919
rect 418526 241224 418582 241233
rect 418526 241159 418582 241168
rect 418540 216918 418568 241159
rect 533988 237380 534040 237386
rect 533988 237322 534040 237328
rect 486422 237144 486478 237153
rect 486422 237079 486478 237088
rect 481548 235000 481600 235006
rect 481548 234942 481600 234948
rect 454132 231736 454184 231742
rect 454132 231678 454184 231684
rect 428924 229084 428976 229090
rect 428924 229026 428976 229032
rect 422300 227656 422352 227662
rect 422300 227598 422352 227604
rect 420460 227384 420512 227390
rect 420460 227326 420512 227332
rect 418804 227180 418856 227186
rect 418804 227122 418856 227128
rect 418816 217410 418844 227122
rect 419724 226160 419776 226166
rect 419724 226102 419776 226108
rect 419736 217410 419764 226102
rect 420472 217410 420500 227326
rect 421288 226296 421340 226302
rect 421288 226238 421340 226244
rect 421300 217410 421328 226238
rect 422312 217410 422340 227598
rect 427176 227588 427228 227594
rect 427176 227530 427228 227536
rect 423864 227520 423916 227526
rect 423864 227462 423916 227468
rect 423036 226024 423088 226030
rect 423036 225966 423088 225972
rect 423048 217410 423076 225966
rect 423876 217410 423904 227462
rect 425520 227452 425572 227458
rect 425520 227394 425572 227400
rect 425060 225820 425112 225826
rect 425060 225762 425112 225768
rect 425072 217410 425100 225762
rect 418816 217382 419152 217410
rect 419736 217382 419980 217410
rect 420472 217382 420808 217410
rect 421300 217382 421636 217410
rect 422312 217382 422464 217410
rect 423048 217382 423384 217410
rect 423876 217382 424212 217410
rect 425040 217382 425100 217410
rect 425532 217410 425560 227394
rect 426348 226092 426400 226098
rect 426348 226034 426400 226040
rect 426360 217410 426388 226034
rect 427188 217410 427216 227530
rect 428004 225888 428056 225894
rect 428004 225830 428056 225836
rect 428016 217410 428044 225830
rect 428936 217410 428964 229026
rect 432236 229016 432288 229022
rect 432236 228958 432288 228964
rect 430580 228812 430632 228818
rect 430580 228754 430632 228760
rect 429752 225956 429804 225962
rect 429752 225898 429804 225904
rect 429764 217410 429792 225898
rect 430592 217410 430620 228754
rect 431408 225616 431460 225622
rect 431408 225558 431460 225564
rect 431420 217410 431448 225558
rect 432248 217410 432276 228958
rect 435640 228948 435692 228954
rect 435640 228890 435692 228896
rect 433892 228880 433944 228886
rect 433892 228822 433944 228828
rect 433340 225752 433392 225758
rect 433340 225694 433392 225700
rect 433352 217410 433380 225694
rect 433904 217410 433932 228822
rect 434812 225684 434864 225690
rect 434812 225626 434864 225632
rect 434824 217410 434852 225626
rect 435652 217410 435680 228890
rect 440700 228744 440752 228750
rect 440700 228686 440752 228692
rect 437296 228676 437348 228682
rect 437296 228618 437348 228624
rect 436468 225412 436520 225418
rect 436468 225354 436520 225360
rect 436480 217410 436508 225354
rect 437308 217410 437336 228618
rect 438952 228608 439004 228614
rect 438952 228550 439004 228556
rect 438124 225548 438176 225554
rect 438124 225490 438176 225496
rect 438136 217410 438164 225490
rect 438964 217410 438992 228550
rect 439780 225480 439832 225486
rect 439780 225422 439832 225428
rect 439792 217410 439820 225422
rect 440712 217410 440740 228686
rect 442356 228540 442408 228546
rect 442356 228482 442408 228488
rect 441620 225344 441672 225350
rect 441620 225286 441672 225292
rect 441632 217410 441660 225286
rect 442368 217410 442396 228482
rect 445668 228472 445720 228478
rect 445668 228414 445720 228420
rect 444380 228404 444432 228410
rect 444380 228346 444432 228352
rect 443184 225208 443236 225214
rect 443184 225150 443236 225156
rect 443196 217410 443224 225150
rect 444392 217410 444420 228346
rect 444840 225140 444892 225146
rect 444840 225082 444892 225088
rect 425532 217382 425868 217410
rect 426360 217382 426696 217410
rect 427188 217382 427524 217410
rect 428016 217382 428352 217410
rect 428936 217382 429272 217410
rect 429764 217382 430100 217410
rect 430592 217382 430928 217410
rect 431420 217382 431756 217410
rect 432248 217382 432584 217410
rect 433352 217382 433412 217410
rect 433904 217382 434240 217410
rect 434824 217382 435160 217410
rect 435652 217382 435988 217410
rect 436480 217382 436816 217410
rect 437308 217382 437644 217410
rect 438136 217382 438472 217410
rect 438964 217382 439300 217410
rect 439792 217382 440128 217410
rect 440712 217382 441048 217410
rect 441632 217382 441876 217410
rect 442368 217382 442704 217410
rect 443196 217382 443532 217410
rect 444360 217382 444420 217410
rect 444852 217410 444880 225082
rect 445680 217410 445708 228414
rect 447416 228336 447468 228342
rect 447416 228278 447468 228284
rect 446588 225276 446640 225282
rect 446588 225218 446640 225224
rect 446600 217410 446628 225218
rect 447428 217410 447456 228278
rect 449072 228268 449124 228274
rect 449072 228210 449124 228216
rect 448244 225072 448296 225078
rect 448244 225014 448296 225020
rect 448256 217410 448284 225014
rect 449084 217410 449112 228210
rect 450728 228200 450780 228206
rect 450728 228142 450780 228148
rect 449900 224936 449952 224942
rect 449900 224878 449952 224884
rect 449912 217410 449940 224878
rect 450740 217410 450768 228142
rect 452660 228132 452712 228138
rect 452660 228074 452712 228080
rect 451554 226128 451610 226137
rect 451554 226063 451610 226072
rect 451568 217410 451596 226063
rect 452672 217410 452700 228074
rect 453304 225004 453356 225010
rect 453304 224946 453356 224952
rect 453316 217410 453344 224946
rect 454144 217410 454172 231678
rect 457444 231668 457496 231674
rect 457444 231610 457496 231616
rect 455788 227996 455840 228002
rect 455788 227938 455840 227944
rect 454958 225992 455014 226001
rect 454958 225927 455014 225936
rect 454972 217410 455000 225927
rect 455800 217410 455828 227938
rect 456614 225720 456670 225729
rect 456614 225655 456670 225664
rect 456628 217410 456656 225655
rect 457456 217410 457484 231610
rect 464252 231600 464304 231606
rect 464252 231542 464304 231548
rect 460940 231532 460992 231538
rect 460940 231474 460992 231480
rect 459192 228064 459244 228070
rect 459192 228006 459244 228012
rect 458364 227928 458416 227934
rect 458364 227870 458416 227876
rect 458376 217410 458404 227870
rect 459204 217410 459232 228006
rect 460018 225856 460074 225865
rect 460018 225791 460074 225800
rect 460032 217410 460060 225791
rect 460952 217410 460980 231474
rect 461676 227792 461728 227798
rect 461676 227734 461728 227740
rect 461688 217410 461716 227734
rect 462504 227724 462556 227730
rect 462504 227666 462556 227672
rect 462516 217410 462544 227666
rect 463698 225584 463754 225593
rect 463698 225519 463754 225528
rect 463712 217410 463740 225519
rect 444852 217382 445188 217410
rect 445680 217382 446016 217410
rect 446600 217382 446936 217410
rect 447428 217382 447764 217410
rect 448256 217382 448592 217410
rect 449084 217382 449420 217410
rect 449912 217382 450248 217410
rect 450740 217382 451076 217410
rect 451568 217382 451904 217410
rect 452672 217382 452824 217410
rect 453316 217382 453652 217410
rect 454144 217382 454480 217410
rect 454972 217382 455308 217410
rect 455800 217382 456136 217410
rect 456628 217382 456964 217410
rect 457456 217382 457792 217410
rect 458376 217382 458712 217410
rect 459204 217382 459540 217410
rect 460032 217382 460368 217410
rect 460952 217382 461196 217410
rect 461688 217382 462024 217410
rect 462516 217382 462852 217410
rect 463680 217382 463740 217410
rect 464264 217410 464292 231542
rect 470968 231464 471020 231470
rect 470968 231406 471020 231412
rect 467564 231396 467616 231402
rect 467564 231338 467616 231344
rect 465078 228848 465134 228857
rect 465078 228783 465134 228792
rect 465092 217410 465120 228783
rect 465908 227860 465960 227866
rect 465908 227802 465960 227808
rect 465920 217410 465948 227802
rect 466734 225448 466790 225457
rect 466734 225383 466790 225392
rect 466748 217410 466776 225383
rect 467576 217410 467604 231338
rect 468390 228712 468446 228721
rect 468390 228647 468446 228656
rect 468404 217410 468432 228647
rect 469218 228440 469274 228449
rect 469218 228375 469274 228384
rect 469232 217410 469260 228375
rect 470138 225176 470194 225185
rect 470138 225111 470194 225120
rect 470152 217410 470180 225111
rect 470980 217410 471008 231406
rect 474280 231328 474332 231334
rect 474280 231270 474332 231276
rect 472622 228576 472678 228585
rect 472622 228511 472678 228520
rect 471978 228032 472034 228041
rect 471978 227967 472034 227976
rect 471992 217410 472020 227967
rect 472636 217410 472664 228511
rect 473450 225312 473506 225321
rect 473450 225247 473506 225256
rect 473464 217410 473492 225247
rect 474292 217410 474320 231270
rect 477684 231260 477736 231266
rect 477684 231202 477736 231208
rect 476026 228304 476082 228313
rect 476026 228239 476082 228248
rect 475106 228168 475162 228177
rect 475106 228103 475162 228112
rect 475120 217410 475148 228103
rect 476040 217410 476068 228239
rect 476854 225040 476910 225049
rect 476854 224975 476910 224984
rect 476868 217410 476896 224975
rect 477696 217410 477724 231202
rect 480996 231192 481048 231198
rect 480996 231134 481048 231140
rect 479338 227896 479394 227905
rect 479338 227831 479394 227840
rect 478510 227624 478566 227633
rect 478510 227559 478566 227568
rect 478524 217410 478552 227559
rect 479352 217410 479380 227831
rect 480258 224904 480314 224913
rect 480258 224839 480314 224848
rect 480272 217410 480300 224839
rect 481008 217410 481036 231134
rect 481560 221270 481588 234942
rect 483020 231124 483072 231130
rect 483020 231066 483072 231072
rect 481914 227760 481970 227769
rect 481914 227695 481970 227704
rect 481548 221264 481600 221270
rect 481548 221206 481600 221212
rect 481928 217410 481956 227695
rect 483032 217410 483060 231066
rect 483846 223408 483902 223417
rect 483846 223343 483902 223352
rect 483860 217410 483888 223343
rect 484400 221468 484452 221474
rect 484400 221410 484452 221416
rect 484412 217410 484440 221410
rect 485228 221196 485280 221202
rect 485228 221138 485280 221144
rect 485240 217410 485268 221138
rect 464264 217382 464600 217410
rect 465092 217382 465428 217410
rect 465920 217382 466256 217410
rect 466748 217382 467084 217410
rect 467576 217382 467912 217410
rect 468404 217382 468740 217410
rect 469232 217382 469568 217410
rect 470152 217382 470488 217410
rect 470980 217382 471316 217410
rect 471992 217382 472144 217410
rect 472636 217382 472972 217410
rect 473464 217382 473800 217410
rect 474292 217382 474628 217410
rect 475120 217382 475456 217410
rect 476040 217382 476376 217410
rect 476868 217382 477204 217410
rect 477696 217382 478032 217410
rect 478524 217382 478860 217410
rect 479352 217382 479688 217410
rect 480272 217382 480516 217410
rect 481008 217382 481344 217410
rect 481928 217382 482264 217410
rect 483032 217382 483092 217410
rect 483860 217382 484256 217410
rect 484412 217382 484748 217410
rect 485240 217382 485576 217410
rect 418528 216912 418580 216918
rect 418528 216854 418580 216860
rect 418436 216776 418488 216782
rect 418436 216718 418488 216724
rect 59268 216640 59320 216646
rect 59268 216582 59320 216588
rect 418160 216640 418212 216646
rect 418160 216582 418212 216588
rect 484228 216442 484256 217382
rect 486436 216458 486464 237079
rect 492310 237008 492366 237017
rect 492310 236943 492366 236952
rect 489828 235068 489880 235074
rect 489828 235010 489880 235016
rect 487160 231056 487212 231062
rect 487160 230998 487212 231004
rect 487172 218142 487200 230998
rect 489458 223272 489514 223281
rect 489458 223207 489514 223216
rect 488630 223136 488686 223145
rect 488630 223071 488686 223080
rect 487804 221264 487856 221270
rect 488644 221241 488672 223071
rect 487804 221206 487856 221212
rect 488630 221232 488686 221241
rect 487160 218136 487212 218142
rect 487160 218078 487212 218084
rect 487172 217410 487200 218078
rect 487816 217410 487844 221206
rect 488630 221167 488686 221176
rect 488644 217410 488672 221167
rect 487172 217382 487232 217410
rect 487816 217382 488152 217410
rect 488644 217382 488980 217410
rect 489472 216458 489500 223207
rect 489840 221270 489868 235010
rect 489920 233504 489972 233510
rect 489920 233446 489972 233452
rect 489932 226334 489960 233446
rect 489932 226306 490236 226334
rect 489828 221264 489880 221270
rect 489828 221206 489880 221212
rect 490208 220862 490236 226306
rect 491300 221400 491352 221406
rect 491300 221342 491352 221348
rect 490196 220856 490248 220862
rect 490196 220798 490248 220804
rect 490208 217410 490236 220798
rect 491312 217410 491340 221342
rect 492324 217410 492352 236943
rect 492586 236872 492642 236881
rect 492586 236807 492642 236816
rect 492600 226334 492628 236807
rect 497002 236736 497058 236745
rect 497002 236671 497058 236680
rect 495348 235136 495400 235142
rect 495348 235078 495400 235084
rect 492600 226306 492720 226334
rect 492692 220969 492720 226306
rect 495360 223582 495388 235078
rect 494336 223576 494388 223582
rect 494336 223518 494388 223524
rect 495348 223576 495400 223582
rect 495348 223518 495400 223524
rect 494058 222864 494114 222873
rect 494058 222799 494114 222808
rect 494072 221105 494100 222799
rect 494058 221096 494114 221105
rect 494058 221031 494114 221040
rect 492678 220960 492734 220969
rect 492678 220895 492734 220904
rect 492692 217410 492720 220895
rect 494348 217410 494376 223518
rect 495346 223000 495402 223009
rect 495346 222935 495402 222944
rect 494520 221332 494572 221338
rect 494520 221274 494572 221280
rect 490208 217382 490636 217410
rect 491312 217382 491464 217410
rect 492292 217394 492628 217410
rect 492292 217388 492640 217394
rect 492292 217382 492588 217388
rect 492692 217382 493120 217410
rect 494040 217382 494376 217410
rect 494532 217410 494560 221274
rect 494532 217382 494868 217410
rect 492588 217330 492640 217336
rect 495360 216594 495388 222935
rect 496450 221096 496506 221105
rect 496450 221031 496506 221040
rect 496464 217410 496492 221031
rect 496464 217382 496524 217410
rect 495360 216578 496032 216594
rect 495360 216572 496044 216578
rect 495360 216566 495992 216572
rect 495992 216514 496044 216520
rect 497016 216510 497044 236671
rect 502706 236600 502762 236609
rect 502706 236535 502762 236544
rect 499946 236464 500002 236473
rect 499946 236399 500002 236408
rect 499488 223508 499540 223514
rect 499488 223450 499540 223456
rect 499500 221610 499528 223450
rect 497372 221604 497424 221610
rect 497372 221546 497424 221552
rect 499488 221604 499540 221610
rect 499488 221546 499540 221552
rect 497384 217410 497412 221546
rect 497832 221264 497884 221270
rect 497832 221206 497884 221212
rect 497352 217382 497412 217410
rect 497844 217410 497872 221206
rect 499960 217410 499988 236399
rect 500868 235204 500920 235210
rect 500868 235146 500920 235152
rect 500880 223378 500908 235146
rect 500868 223372 500920 223378
rect 500868 223314 500920 223320
rect 500880 217410 500908 223314
rect 502614 222592 502670 222601
rect 502614 222527 502670 222536
rect 501236 221536 501288 221542
rect 502628 221513 502656 222527
rect 501236 221478 501288 221484
rect 502614 221504 502670 221513
rect 497844 217382 498180 217410
rect 499928 217382 500264 217410
rect 497004 216504 497056 216510
rect 486404 216442 486740 216458
rect 489472 216442 490144 216458
rect 499304 216504 499356 216510
rect 497004 216446 497056 216452
rect 499008 216452 499304 216458
rect 499008 216446 499356 216452
rect 484216 216436 484268 216442
rect 486404 216436 486752 216442
rect 486404 216430 486700 216436
rect 484216 216378 484268 216384
rect 489472 216436 490156 216442
rect 489472 216430 490104 216436
rect 486700 216378 486752 216384
rect 499008 216430 499344 216446
rect 500236 216442 500264 217382
rect 500316 217388 500368 217394
rect 500756 217382 500908 217410
rect 501248 217410 501276 221478
rect 502614 221439 502670 221448
rect 502628 217410 502656 221439
rect 502720 217530 502748 236535
rect 507858 236328 507914 236337
rect 507858 236263 507914 236272
rect 506388 235340 506440 235346
rect 506388 235282 506440 235288
rect 502800 235272 502852 235278
rect 502800 235214 502852 235220
rect 502812 226334 502840 235214
rect 506400 226334 506428 235282
rect 502812 226306 503668 226334
rect 503536 221876 503588 221882
rect 503536 221818 503588 221824
rect 503548 221134 503576 221818
rect 503536 221128 503588 221134
rect 503536 221070 503588 221076
rect 502708 217524 502760 217530
rect 502708 217466 502760 217472
rect 503548 217410 503576 221070
rect 501248 217382 501584 217410
rect 502412 217382 502656 217410
rect 503240 217382 503576 217410
rect 503640 217410 503668 226306
rect 506124 226306 506428 226334
rect 506124 221202 506152 226306
rect 507122 222728 507178 222737
rect 507122 222663 507178 222672
rect 506296 221672 506348 221678
rect 506296 221614 506348 221620
rect 506112 221196 506164 221202
rect 506112 221138 506164 221144
rect 504870 217524 504922 217530
rect 504870 217466 504922 217472
rect 504882 217410 504910 217466
rect 506124 217410 506152 221138
rect 503640 217382 504068 217410
rect 504882 217396 505048 217410
rect 504896 217382 505048 217396
rect 505816 217382 506152 217410
rect 506308 217410 506336 221614
rect 507136 221377 507164 222663
rect 507122 221368 507178 221377
rect 507122 221303 507178 221312
rect 507136 217410 507164 221303
rect 507872 217666 507900 236263
rect 513746 236192 513802 236201
rect 513746 236127 513802 236136
rect 512000 235612 512052 235618
rect 512000 235554 512052 235560
rect 511908 235476 511960 235482
rect 511908 235418 511960 235424
rect 507952 235408 508004 235414
rect 507952 235350 508004 235356
rect 507964 226334 507992 235350
rect 507964 226306 508728 226334
rect 507952 222012 508004 222018
rect 507952 221954 508004 221960
rect 507964 221406 507992 221954
rect 507952 221400 508004 221406
rect 507952 221342 508004 221348
rect 507860 217660 507912 217666
rect 507860 217602 507912 217608
rect 507964 217410 507992 221342
rect 508700 217410 508728 226306
rect 510618 222456 510674 222465
rect 510618 222391 510674 222400
rect 510632 221649 510660 222391
rect 511356 221944 511408 221950
rect 511356 221886 511408 221892
rect 510618 221640 510674 221649
rect 510618 221575 510674 221584
rect 511080 221264 511132 221270
rect 511080 221206 511132 221212
rect 509930 217660 509982 217666
rect 509930 217602 509982 217608
rect 509942 217410 509970 217602
rect 511092 217410 511120 221206
rect 506308 217382 506644 217410
rect 507136 217382 507472 217410
rect 507964 217382 508300 217410
rect 508700 217382 509128 217410
rect 509942 217396 510292 217410
rect 509956 217382 510292 217396
rect 510784 217382 511120 217410
rect 511368 217410 511396 221886
rect 511920 221338 511948 235418
rect 511908 221332 511960 221338
rect 511908 221274 511960 221280
rect 512012 221270 512040 235554
rect 513472 235544 513524 235550
rect 513472 235486 513524 235492
rect 513484 226334 513512 235486
rect 513760 226334 513788 236127
rect 517426 236056 517482 236065
rect 517426 235991 517482 236000
rect 515496 230988 515548 230994
rect 515496 230930 515548 230936
rect 513484 226306 513696 226334
rect 513760 226306 513880 226334
rect 513380 222080 513432 222086
rect 513380 222022 513432 222028
rect 512458 221640 512514 221649
rect 512458 221575 512514 221584
rect 512000 221264 512052 221270
rect 512000 221206 512052 221212
rect 512472 217410 512500 221575
rect 513392 221474 513420 222022
rect 513380 221468 513432 221474
rect 513380 221410 513432 221416
rect 513392 217410 513420 221410
rect 513668 220538 513696 226306
rect 513668 220510 513788 220538
rect 511368 217382 511704 217410
rect 512472 217382 512532 217410
rect 513360 217382 513420 217410
rect 513760 217410 513788 220510
rect 513852 217666 513880 226306
rect 515508 218210 515536 230930
rect 517440 222329 517468 235991
rect 522946 235920 523002 235929
rect 522946 235855 523002 235864
rect 528468 235884 528520 235890
rect 520188 235680 520240 235686
rect 520188 235622 520240 235628
rect 518072 230920 518124 230926
rect 518072 230862 518124 230868
rect 517426 222320 517482 222329
rect 517426 222255 517482 222264
rect 517886 222320 517942 222329
rect 517886 222255 517942 222264
rect 516416 221332 516468 221338
rect 516416 221274 516468 221280
rect 515496 218204 515548 218210
rect 515496 218146 515548 218152
rect 513840 217660 513892 217666
rect 513840 217602 513892 217608
rect 514990 217660 515042 217666
rect 514990 217602 515042 217608
rect 515002 217410 515030 217602
rect 515508 217410 515536 218146
rect 516428 217410 516456 221274
rect 517900 217410 517928 222255
rect 518084 218278 518112 230862
rect 518992 230852 519044 230858
rect 518992 230794 519044 230800
rect 518900 221740 518952 221746
rect 518900 221682 518952 221688
rect 518072 218272 518124 218278
rect 518072 218214 518124 218220
rect 518624 218272 518676 218278
rect 518624 218214 518676 218220
rect 518636 217410 518664 218214
rect 513760 217382 514188 217410
rect 515002 217396 515168 217410
rect 515016 217382 515168 217396
rect 515508 217382 515844 217410
rect 516428 217382 516672 217410
rect 517592 217382 517928 217410
rect 518420 217382 518664 217410
rect 518912 217410 518940 221682
rect 519004 218346 519032 230794
rect 519726 222456 519782 222465
rect 519726 222391 519782 222400
rect 518992 218340 519044 218346
rect 518992 218282 519044 218288
rect 518912 217382 519248 217410
rect 500316 217330 500368 217336
rect 500328 216442 500356 217330
rect 505020 216578 505048 217382
rect 505008 216572 505060 216578
rect 505008 216514 505060 216520
rect 510264 216510 510292 217382
rect 515140 216578 515168 217382
rect 519740 216866 519768 222391
rect 520200 221338 520228 235622
rect 522960 221921 522988 235855
rect 528468 235826 528520 235832
rect 524420 235748 524472 235754
rect 524420 235690 524472 235696
rect 523408 230784 523460 230790
rect 523408 230726 523460 230732
rect 522946 221912 523002 221921
rect 522946 221847 523002 221856
rect 520188 221332 520240 221338
rect 520188 221274 520240 221280
rect 521660 221332 521712 221338
rect 521660 221274 521712 221280
rect 521200 218340 521252 218346
rect 521200 218282 521252 218288
rect 521212 217410 521240 218282
rect 520904 217382 521240 217410
rect 521672 217410 521700 221274
rect 522960 217410 522988 221847
rect 523420 218414 523448 230726
rect 523960 221808 524012 221814
rect 523960 221750 524012 221756
rect 523408 218408 523460 218414
rect 523408 218350 523460 218356
rect 523776 218408 523828 218414
rect 523776 218350 523828 218356
rect 523788 217410 523816 218350
rect 521672 217382 521732 217410
rect 522560 217382 522988 217410
rect 523480 217382 523816 217410
rect 523972 217410 524000 221750
rect 524432 221338 524460 235690
rect 525892 230716 525944 230722
rect 525892 230658 525944 230664
rect 525904 221678 525932 230658
rect 528480 222057 528508 235826
rect 529940 235816 529992 235822
rect 529940 235758 529992 235764
rect 528560 233436 528612 233442
rect 528560 233378 528612 233384
rect 528466 222048 528522 222057
rect 528466 221983 528522 221992
rect 528480 221785 528508 221983
rect 528572 221814 528600 233378
rect 528650 222320 528706 222329
rect 528650 222255 528706 222264
rect 528560 221808 528612 221814
rect 527914 221776 527970 221785
rect 527914 221711 527970 221720
rect 528466 221776 528522 221785
rect 528664 221785 528692 222255
rect 529020 222148 529072 222154
rect 529020 222090 529072 222096
rect 528560 221750 528612 221756
rect 528650 221776 528706 221785
rect 528466 221711 528522 221720
rect 525892 221672 525944 221678
rect 525892 221614 525944 221620
rect 524420 221332 524472 221338
rect 524420 221274 524472 221280
rect 525064 220924 525116 220930
rect 525064 220866 525116 220872
rect 525076 217410 525104 220866
rect 525904 217410 525932 221614
rect 526444 221332 526496 221338
rect 526444 221274 526496 221280
rect 526456 217410 526484 221274
rect 527928 217410 527956 221711
rect 528572 217410 528600 221750
rect 528650 221711 528706 221720
rect 523972 217382 524308 217410
rect 525076 217382 525472 217410
rect 525904 217382 525964 217410
rect 526456 217382 526792 217410
rect 527620 217382 527956 217410
rect 528448 217382 528600 217410
rect 529032 217410 529060 222090
rect 529952 221338 529980 235758
rect 530952 230648 531004 230654
rect 530952 230590 531004 230596
rect 530032 223304 530084 223310
rect 530032 223246 530084 223252
rect 529940 221332 529992 221338
rect 529940 221274 529992 221280
rect 530044 217410 530072 223246
rect 530964 221950 530992 230590
rect 533160 230580 533212 230586
rect 533160 230522 533212 230528
rect 533172 222018 533200 230522
rect 533160 222012 533212 222018
rect 533160 221954 533212 221960
rect 533804 222012 533856 222018
rect 533804 221954 533856 221960
rect 530952 221944 531004 221950
rect 530952 221886 531004 221892
rect 530964 217410 530992 221886
rect 532976 221468 533028 221474
rect 532976 221410 533028 221416
rect 531504 221332 531556 221338
rect 531504 221274 531556 221280
rect 531516 217410 531544 221274
rect 532988 217410 533016 221410
rect 533816 217410 533844 221954
rect 534000 221474 534028 237322
rect 535460 237312 535512 237318
rect 535460 237254 535512 237260
rect 535472 226334 535500 237254
rect 539508 237244 539560 237250
rect 539508 237186 539560 237192
rect 536748 235952 536800 235958
rect 536748 235894 536800 235900
rect 535472 226306 536512 226334
rect 536288 222964 536340 222970
rect 536288 222906 536340 222912
rect 536380 222964 536432 222970
rect 536380 222906 536432 222912
rect 536300 222154 536328 222906
rect 536288 222148 536340 222154
rect 536288 222090 536340 222096
rect 533988 221468 534040 221474
rect 533988 221410 534040 221416
rect 533988 221060 534040 221066
rect 533988 221002 534040 221008
rect 529032 217382 529368 217410
rect 530044 217382 530348 217410
rect 530964 217382 531024 217410
rect 531516 217382 531852 217410
rect 532680 217382 533016 217410
rect 533508 217382 533844 217410
rect 534000 217410 534028 221002
rect 534908 220992 534960 220998
rect 534908 220934 534960 220940
rect 534920 217410 534948 220934
rect 536392 217410 536420 222906
rect 534000 217382 534336 217410
rect 534920 217382 535408 217410
rect 536084 217382 536420 217410
rect 536484 217410 536512 226306
rect 536760 221610 536788 235894
rect 536840 233368 536892 233374
rect 536840 233310 536892 233316
rect 536852 222970 536880 233310
rect 539048 223440 539100 223446
rect 539048 223382 539100 223388
rect 538864 223304 538916 223310
rect 538864 223246 538916 223252
rect 536840 222964 536892 222970
rect 536840 222906 536892 222912
rect 536748 221604 536800 221610
rect 536748 221546 536800 221552
rect 538036 221604 538088 221610
rect 538036 221546 538088 221552
rect 538048 217410 538076 221546
rect 538876 217410 538904 223246
rect 536484 217382 536912 217410
rect 537740 217382 538076 217410
rect 538568 217382 538904 217410
rect 539060 217410 539088 223382
rect 539520 221542 539548 237186
rect 542268 237176 542320 237182
rect 542268 237118 542320 237124
rect 539600 233300 539652 233306
rect 539600 233242 539652 233248
rect 539612 223310 539640 233242
rect 539600 223304 539652 223310
rect 539600 223246 539652 223252
rect 539876 223236 539928 223242
rect 539876 223178 539928 223184
rect 539508 221536 539560 221542
rect 539508 221478 539560 221484
rect 539060 217382 539396 217410
rect 525444 216986 525472 217382
rect 530320 217122 530348 217382
rect 530308 217116 530360 217122
rect 530308 217058 530360 217064
rect 535380 217054 535408 217382
rect 539888 217138 539916 223178
rect 542176 223100 542228 223106
rect 542176 223042 542228 223048
rect 541440 221876 541492 221882
rect 541440 221818 541492 221824
rect 541452 217410 541480 221818
rect 541624 221536 541676 221542
rect 541624 221478 541676 221484
rect 541144 217382 541480 217410
rect 541636 217410 541664 221478
rect 542188 221066 542216 223042
rect 542280 221542 542308 237118
rect 545120 237108 545172 237114
rect 545120 237050 545172 237056
rect 545028 237040 545080 237046
rect 545028 236982 545080 236988
rect 542360 236972 542412 236978
rect 542360 236914 542412 236920
rect 542372 223106 542400 236914
rect 542452 233232 542504 233238
rect 542452 233174 542504 233180
rect 542464 223242 542492 233174
rect 542452 223236 542504 223242
rect 542452 223178 542504 223184
rect 543648 223236 543700 223242
rect 543648 223178 543700 223184
rect 542360 223100 542412 223106
rect 542360 223042 542412 223048
rect 542372 221882 542400 223042
rect 542360 221876 542412 221882
rect 542360 221818 542412 221824
rect 542268 221536 542320 221542
rect 542268 221478 542320 221484
rect 542176 221060 542228 221066
rect 542176 221002 542228 221008
rect 543096 221060 543148 221066
rect 543096 221002 543148 221008
rect 543108 217410 543136 221002
rect 543660 217410 543688 223178
rect 544936 223032 544988 223038
rect 544936 222974 544988 222980
rect 544948 222086 544976 222974
rect 544936 222080 544988 222086
rect 544936 222022 544988 222028
rect 545040 221746 545068 236982
rect 545132 223038 545160 237050
rect 550364 236904 550416 236910
rect 550364 236846 550416 236852
rect 547788 236768 547840 236774
rect 547788 236710 547840 236716
rect 546040 223440 546092 223446
rect 546040 223382 546092 223388
rect 546052 223038 546080 223382
rect 546960 223304 547012 223310
rect 546960 223246 547012 223252
rect 546684 223168 546736 223174
rect 546684 223110 546736 223116
rect 545120 223032 545172 223038
rect 545120 222974 545172 222980
rect 546040 223032 546092 223038
rect 546040 222974 546092 222980
rect 545028 221740 545080 221746
rect 545028 221682 545080 221688
rect 544108 221536 544160 221542
rect 544108 221478 544160 221484
rect 541636 217382 541972 217410
rect 542800 217382 543136 217410
rect 543628 217382 543688 217410
rect 544120 217410 544148 221478
rect 545040 217410 545068 221682
rect 546052 217410 546080 222974
rect 546696 217410 546724 223110
rect 546972 222970 547000 223246
rect 546960 222964 547012 222970
rect 546960 222906 547012 222912
rect 547512 222080 547564 222086
rect 547512 222022 547564 222028
rect 547524 221882 547552 222022
rect 547512 221876 547564 221882
rect 547512 221818 547564 221824
rect 547524 217410 547552 221818
rect 547800 221542 547828 236710
rect 548340 222148 548392 222154
rect 548340 222090 548392 222096
rect 547788 221536 547840 221542
rect 547788 221478 547840 221484
rect 548352 220930 548380 222090
rect 549260 221536 549312 221542
rect 549260 221478 549312 221484
rect 548340 220924 548392 220930
rect 548340 220866 548392 220872
rect 548352 217410 548380 220866
rect 549272 217410 549300 221478
rect 550376 217410 550404 236846
rect 550548 236836 550600 236842
rect 550548 236778 550600 236784
rect 550560 222970 550588 236778
rect 552296 236700 552348 236706
rect 552296 236642 552348 236648
rect 550548 222964 550600 222970
rect 550548 222906 550600 222912
rect 551468 222964 551520 222970
rect 551468 222906 551520 222912
rect 551480 217410 551508 222906
rect 552020 222896 552072 222902
rect 552020 222838 552072 222844
rect 552032 217410 552060 222838
rect 552204 222760 552256 222766
rect 552204 222702 552256 222708
rect 552112 222692 552164 222698
rect 552112 222634 552164 222640
rect 552124 222086 552152 222634
rect 552112 222080 552164 222086
rect 552112 222022 552164 222028
rect 552216 220998 552244 222702
rect 552308 221542 552336 236642
rect 557540 236632 557592 236638
rect 557540 236574 557592 236580
rect 556160 236564 556212 236570
rect 556160 236506 556212 236512
rect 556068 236496 556120 236502
rect 556068 236438 556120 236444
rect 555056 222760 555108 222766
rect 555056 222702 555108 222708
rect 552848 222080 552900 222086
rect 552848 222022 552900 222028
rect 552296 221536 552348 221542
rect 552296 221478 552348 221484
rect 552204 220992 552256 220998
rect 552204 220934 552256 220940
rect 544120 217382 544456 217410
rect 545040 217382 545284 217410
rect 546052 217382 546112 217410
rect 546696 217382 547032 217410
rect 547524 217382 547860 217410
rect 548352 217382 548688 217410
rect 549272 217382 549516 217410
rect 550344 217382 550680 217410
rect 551172 217382 551508 217410
rect 552000 217382 552060 217410
rect 552860 217410 552888 222022
rect 554412 221604 554464 221610
rect 554412 221546 554464 221552
rect 554228 221536 554280 221542
rect 554228 221478 554280 221484
rect 553676 220992 553728 220998
rect 553676 220934 553728 220940
rect 553688 217410 553716 220934
rect 554240 217410 554268 221478
rect 554424 221066 554452 221546
rect 555068 221066 555096 222702
rect 556080 222698 556108 236438
rect 556068 222692 556120 222698
rect 556068 222634 556120 222640
rect 555424 222488 555476 222494
rect 555424 222430 555476 222436
rect 555436 222358 555464 222430
rect 555424 222352 555476 222358
rect 555424 222294 555476 222300
rect 555700 222216 555752 222222
rect 555700 222158 555752 222164
rect 554412 221060 554464 221066
rect 554412 221002 554464 221008
rect 555056 221060 555108 221066
rect 555056 221002 555108 221008
rect 555712 217410 555740 222158
rect 552860 217382 552920 217410
rect 553688 217382 553748 217410
rect 554240 217382 554576 217410
rect 555404 217382 555740 217410
rect 556080 217410 556108 222634
rect 556172 222222 556200 236506
rect 556160 222216 556212 222222
rect 556160 222158 556212 222164
rect 557552 221066 557580 236574
rect 563152 236428 563204 236434
rect 563152 236370 563204 236376
rect 561588 236292 561640 236298
rect 561588 236234 561640 236240
rect 557908 222896 557960 222902
rect 557908 222838 557960 222844
rect 556804 221060 556856 221066
rect 556804 221002 556856 221008
rect 557540 221060 557592 221066
rect 557540 221002 557592 221008
rect 556816 217410 556844 221002
rect 557920 217410 557948 222838
rect 559104 222828 559156 222834
rect 559104 222770 559156 222776
rect 559116 217410 559144 222770
rect 561600 222562 561628 236234
rect 561680 236224 561732 236230
rect 561680 236166 561732 236172
rect 561692 222766 561720 236166
rect 561680 222760 561732 222766
rect 561680 222702 561732 222708
rect 561588 222556 561640 222562
rect 561588 222498 561640 222504
rect 561600 222154 561628 222498
rect 560760 222148 560812 222154
rect 560760 222090 560812 222096
rect 561588 222148 561640 222154
rect 561588 222090 561640 222096
rect 559288 221060 559340 221066
rect 559288 221002 559340 221008
rect 556080 217382 556232 217410
rect 556816 217382 557060 217410
rect 557888 217382 557948 217410
rect 558808 217382 559144 217410
rect 559300 217410 559328 221002
rect 560772 217410 560800 222090
rect 561692 217410 561720 222702
rect 562876 222488 562928 222494
rect 562876 222430 562928 222436
rect 561772 222420 561824 222426
rect 561772 222362 561824 222368
rect 559300 217382 559636 217410
rect 560464 217382 560800 217410
rect 561292 217382 561720 217410
rect 561784 217410 561812 222362
rect 562888 217410 562916 222430
rect 563164 221066 563192 236370
rect 565544 236360 565596 236366
rect 565544 236302 565596 236308
rect 564072 222896 564124 222902
rect 564072 222838 564124 222844
rect 564084 222630 564112 222838
rect 563980 222624 564032 222630
rect 563980 222566 564032 222572
rect 564072 222624 564124 222630
rect 564072 222566 564124 222572
rect 563992 222494 564020 222566
rect 563980 222488 564032 222494
rect 563980 222430 564032 222436
rect 563152 221060 563204 221066
rect 563152 221002 563204 221008
rect 563992 217410 564020 222430
rect 564348 221060 564400 221066
rect 564348 221002 564400 221008
rect 561784 217382 562120 217410
rect 562888 217382 563100 217410
rect 563776 217382 564020 217410
rect 564360 217410 564388 221002
rect 565556 217410 565584 236302
rect 565820 236156 565872 236162
rect 565820 236098 565872 236104
rect 565832 226334 565860 236098
rect 568028 236088 568080 236094
rect 568028 236030 568080 236036
rect 565832 226306 566780 226334
rect 566004 222284 566056 222290
rect 566004 222226 566056 222232
rect 566016 217410 566044 222226
rect 566752 217410 566780 226306
rect 568040 217410 568068 236030
rect 569880 222193 569908 248406
rect 569960 236020 570012 236026
rect 569960 235962 570012 235968
rect 569972 222358 570000 235962
rect 570236 222420 570288 222426
rect 570236 222362 570288 222368
rect 569960 222352 570012 222358
rect 569960 222294 570012 222300
rect 569314 222184 569370 222193
rect 569132 222148 569184 222154
rect 569314 222119 569370 222128
rect 569866 222184 569922 222193
rect 569972 222154 570000 222294
rect 569866 222119 569922 222128
rect 569960 222148 570012 222154
rect 569132 222090 569184 222096
rect 568304 217456 568356 217462
rect 564360 217382 564696 217410
rect 565524 217394 565768 217410
rect 565524 217388 565780 217394
rect 565524 217382 565728 217388
rect 550652 217258 550680 217382
rect 563072 217326 563100 217382
rect 566016 217382 566352 217410
rect 566752 217382 567180 217410
rect 568008 217404 568304 217410
rect 569144 217410 569172 222090
rect 568008 217398 568356 217404
rect 568008 217382 568344 217398
rect 568836 217382 569172 217410
rect 569328 217410 569356 222119
rect 569960 222090 570012 222096
rect 570248 217410 570276 222362
rect 570558 217524 570610 217530
rect 570558 217466 570610 217472
rect 570570 217410 570598 217466
rect 571536 217410 571564 256702
rect 571720 221066 571748 262210
rect 571800 259480 571852 259486
rect 571800 259422 571852 259428
rect 571708 221060 571760 221066
rect 571708 221002 571760 221008
rect 569328 217382 569664 217410
rect 570248 217396 570598 217410
rect 570248 217382 570584 217396
rect 571412 217382 571564 217410
rect 571812 217410 571840 259422
rect 574100 253972 574152 253978
rect 574100 253914 574152 253920
rect 572628 251252 572680 251258
rect 572628 251194 572680 251200
rect 572640 222601 572668 251194
rect 574112 226334 574140 253914
rect 574112 226306 575152 226334
rect 572812 222828 572864 222834
rect 572812 222770 572864 222776
rect 572626 222592 572682 222601
rect 572626 222527 572682 222536
rect 572824 221066 572852 222770
rect 574374 222592 574430 222601
rect 574374 222527 574430 222536
rect 573546 222184 573602 222193
rect 573546 222119 573602 222128
rect 572720 221060 572772 221066
rect 572720 221002 572772 221008
rect 572812 221060 572864 221066
rect 572812 221002 572864 221008
rect 572732 217410 572760 221002
rect 573560 217410 573588 222119
rect 574388 217410 574416 222527
rect 575124 217410 575152 226306
rect 607588 223576 607640 223582
rect 607588 223518 607640 223524
rect 607128 220856 607180 220862
rect 607128 220798 607180 220804
rect 606668 218136 606720 218142
rect 606668 218078 606720 218084
rect 571812 217382 572240 217410
rect 572732 217382 573068 217410
rect 573560 217382 573896 217410
rect 574388 217382 574724 217410
rect 575124 217382 575552 217410
rect 565728 217330 565780 217336
rect 563060 217320 563112 217326
rect 563060 217262 563112 217268
rect 550640 217252 550692 217258
rect 550640 217194 550692 217200
rect 540520 217184 540572 217190
rect 539888 217132 540520 217138
rect 539888 217126 540572 217132
rect 539888 217110 540560 217126
rect 535368 217048 535420 217054
rect 535368 216990 535420 216996
rect 525432 216980 525484 216986
rect 525432 216922 525484 216928
rect 519740 216850 520412 216866
rect 519740 216844 520424 216850
rect 519740 216838 520372 216844
rect 520372 216786 520424 216792
rect 515128 216572 515180 216578
rect 515128 216514 515180 216520
rect 502524 216504 502576 216510
rect 510252 216504 510304 216510
rect 502576 216452 502748 216458
rect 502524 216446 502748 216452
rect 510252 216446 510304 216452
rect 502536 216442 502748 216446
rect 500224 216436 500276 216442
rect 490104 216378 490156 216384
rect 500224 216378 500276 216384
rect 500316 216436 500368 216442
rect 502536 216436 502760 216442
rect 502536 216430 502708 216436
rect 500316 216378 500368 216384
rect 502708 216378 502760 216384
rect 579710 216200 579766 216209
rect 579710 216135 579766 216144
rect 579724 215694 579752 216135
rect 579712 215688 579764 215694
rect 579712 215630 579764 215636
rect 599768 215688 599820 215694
rect 599768 215630 599820 215636
rect 582286 214704 582342 214713
rect 582286 214639 582342 214648
rect 580262 213208 580318 213217
rect 580262 213143 580318 213152
rect 580276 212566 580304 213143
rect 582300 212634 582328 214639
rect 582288 212628 582340 212634
rect 582288 212570 582340 212576
rect 580264 212560 580316 212566
rect 580264 212502 580316 212508
rect 581642 211712 581698 211721
rect 581642 211647 581698 211656
rect 580538 210216 580594 210225
rect 580538 210151 580594 210160
rect 580552 209846 580580 210151
rect 581656 209914 581684 211647
rect 581644 209908 581696 209914
rect 581644 209850 581696 209856
rect 580540 209840 580592 209846
rect 580540 209782 580592 209788
rect 599124 209840 599176 209846
rect 599124 209782 599176 209788
rect 581458 208720 581514 208729
rect 581458 208655 581514 208664
rect 581472 207058 581500 208655
rect 582288 207120 582340 207126
rect 582286 207088 582288 207097
rect 582340 207088 582342 207097
rect 581460 207052 581512 207058
rect 582286 207023 582342 207032
rect 581460 206994 581512 207000
rect 582286 205592 582342 205601
rect 582286 205527 582342 205536
rect 582300 204338 582328 205527
rect 599136 205465 599164 209782
rect 599780 209545 599808 215630
rect 599952 212628 600004 212634
rect 599952 212570 600004 212576
rect 599860 212560 599912 212566
rect 599860 212502 599912 212508
rect 599766 209536 599822 209545
rect 599766 209471 599822 209480
rect 599872 207505 599900 212502
rect 599964 208593 599992 212570
rect 606680 210202 606708 218078
rect 607140 210202 607168 220798
rect 607600 210202 607628 223518
rect 608048 223508 608100 223514
rect 608048 223450 608100 223456
rect 608060 210202 608088 223450
rect 616880 223440 616932 223446
rect 616880 223382 616932 223388
rect 608508 223372 608560 223378
rect 608508 223314 608560 223320
rect 608520 210202 608548 223314
rect 615040 223304 615092 223310
rect 615040 223246 615092 223252
rect 614580 222012 614632 222018
rect 614580 221954 614632 221960
rect 614028 221944 614080 221950
rect 614028 221886 614080 221892
rect 613568 221808 613620 221814
rect 613568 221750 613620 221756
rect 613108 221672 613160 221678
rect 613108 221614 613160 221620
rect 610808 221400 610860 221406
rect 610808 221342 610860 221348
rect 609888 221332 609940 221338
rect 609888 221274 609940 221280
rect 609428 221196 609480 221202
rect 609428 221138 609480 221144
rect 608968 221128 609020 221134
rect 608968 221070 609020 221076
rect 608980 210202 609008 221070
rect 609440 210202 609468 221138
rect 609900 210202 609928 221274
rect 610348 221264 610400 221270
rect 610348 221206 610400 221212
rect 610360 210202 610388 221206
rect 610820 210202 610848 221342
rect 612648 218408 612700 218414
rect 612648 218350 612700 218356
rect 612188 218340 612240 218346
rect 612188 218282 612240 218288
rect 611728 218272 611780 218278
rect 611728 218214 611780 218220
rect 611268 218204 611320 218210
rect 611268 218146 611320 218152
rect 611280 210202 611308 218146
rect 611740 210202 611768 218214
rect 612200 210202 612228 218282
rect 612660 210202 612688 218350
rect 613120 210202 613148 221614
rect 613580 210202 613608 221750
rect 614040 210202 614068 221886
rect 614592 210202 614620 221954
rect 615052 210202 615080 223246
rect 615500 223236 615552 223242
rect 615500 223178 615552 223184
rect 615512 210202 615540 223178
rect 616420 223168 616472 223174
rect 616420 223110 616472 223116
rect 615960 223100 616012 223106
rect 615960 223042 616012 223048
rect 615972 210202 616000 223042
rect 616432 210202 616460 223110
rect 616892 210202 616920 223382
rect 617800 222964 617852 222970
rect 617800 222906 617852 222912
rect 617340 220924 617392 220930
rect 617340 220866 617392 220872
rect 617352 210202 617380 220866
rect 617812 210202 617840 222906
rect 619640 222760 619692 222766
rect 619640 222702 619692 222708
rect 618720 222692 618772 222698
rect 618720 222634 618772 222640
rect 618260 220992 618312 220998
rect 618260 220934 618312 220940
rect 618272 210202 618300 220934
rect 618732 210202 618760 222634
rect 619180 221060 619232 221066
rect 619180 221002 619232 221008
rect 619192 210202 619220 221002
rect 619652 210202 619680 222702
rect 633624 222624 633676 222630
rect 633624 222566 633676 222572
rect 620100 222488 620152 222494
rect 620100 222430 620152 222436
rect 620112 210202 620140 222430
rect 621020 222352 621072 222358
rect 621020 222294 621072 222300
rect 620560 222216 620612 222222
rect 620560 222158 620612 222164
rect 620572 210202 620600 222158
rect 621032 210202 621060 222294
rect 633164 222148 633216 222154
rect 633164 222090 633216 222096
rect 632704 222080 632756 222086
rect 628010 222048 628066 222057
rect 632704 222022 632756 222028
rect 628010 221983 628066 221992
rect 627090 221912 627146 221921
rect 627090 221847 627146 221856
rect 626170 221776 626226 221785
rect 626170 221711 626226 221720
rect 625250 221640 625306 221649
rect 625250 221575 625306 221584
rect 623410 221504 623466 221513
rect 623410 221439 623466 221448
rect 621478 221232 621534 221241
rect 621478 221167 621534 221176
rect 621492 210202 621520 221167
rect 622952 216368 623004 216374
rect 622952 216310 623004 216316
rect 622492 216300 622544 216306
rect 622492 216242 622544 216248
rect 622032 216232 622084 216238
rect 622032 216174 622084 216180
rect 622044 210202 622072 216174
rect 622504 210202 622532 216242
rect 622964 210202 622992 216310
rect 623424 210202 623452 221439
rect 624330 221368 624386 221377
rect 624330 221303 624386 221312
rect 623872 216436 623924 216442
rect 623872 216378 623924 216384
rect 623884 210202 623912 216378
rect 624344 210202 624372 221303
rect 624792 216504 624844 216510
rect 624792 216446 624844 216452
rect 624804 210202 624832 216446
rect 625264 210202 625292 221575
rect 625712 216572 625764 216578
rect 625712 216514 625764 216520
rect 625724 210202 625752 216514
rect 626184 210202 626212 221711
rect 626632 216844 626684 216850
rect 626632 216786 626684 216792
rect 626644 210202 626672 216786
rect 627104 210202 627132 221847
rect 627552 216980 627604 216986
rect 627552 216922 627604 216928
rect 627564 210202 627592 216922
rect 628024 210202 628052 221983
rect 631784 221876 631836 221882
rect 631784 221818 631836 221824
rect 631324 221740 631376 221746
rect 631324 221682 631376 221688
rect 630864 221604 630916 221610
rect 630864 221546 630916 221552
rect 629944 221536 629996 221542
rect 629944 221478 629996 221484
rect 628932 221468 628984 221474
rect 628932 221410 628984 221416
rect 628472 217116 628524 217122
rect 628472 217058 628524 217064
rect 628484 210202 628512 217058
rect 628944 210202 628972 221410
rect 629484 217048 629536 217054
rect 629484 216990 629536 216996
rect 629496 210202 629524 216990
rect 629956 210202 629984 221478
rect 630404 217184 630456 217190
rect 630404 217126 630456 217132
rect 630416 210202 630444 217126
rect 630876 210202 630904 221546
rect 631336 210202 631364 221682
rect 631796 210202 631824 221818
rect 632244 217252 632296 217258
rect 632244 217194 632296 217200
rect 632256 210202 632284 217194
rect 632716 210202 632744 222022
rect 633176 210202 633204 222090
rect 633636 210202 633664 222566
rect 634084 222556 634136 222562
rect 634084 222498 634136 222504
rect 634096 210202 634124 222498
rect 637394 221096 637450 221105
rect 637394 221031 637450 221040
rect 636934 220960 636990 220969
rect 636934 220895 636990 220904
rect 635924 217524 635976 217530
rect 635924 217466 635976 217472
rect 635464 217456 635516 217462
rect 635464 217398 635516 217404
rect 635004 217388 635056 217394
rect 635004 217330 635056 217336
rect 634544 217320 634596 217326
rect 634544 217262 634596 217268
rect 634556 210202 634584 217262
rect 635016 210202 635044 217330
rect 635476 210202 635504 217398
rect 635936 210202 635964 217466
rect 636384 216096 636436 216102
rect 636384 216038 636436 216044
rect 636396 210202 636424 216038
rect 636948 210202 636976 220895
rect 637408 210202 637436 221031
rect 647148 220380 647200 220386
rect 647148 220322 647200 220328
rect 646964 218000 647016 218006
rect 646964 217942 647016 217948
rect 644112 217932 644164 217938
rect 644112 217874 644164 217880
rect 639696 216912 639748 216918
rect 639696 216854 639748 216860
rect 637856 216164 637908 216170
rect 637856 216106 637908 216112
rect 637868 210202 637896 216106
rect 638316 216028 638368 216034
rect 638316 215970 638368 215976
rect 638328 210202 638356 215970
rect 638776 215960 638828 215966
rect 638776 215902 638828 215908
rect 638788 210202 638816 215902
rect 639708 210202 639736 216854
rect 640156 216776 640208 216782
rect 640156 216718 640208 216724
rect 640168 210202 640196 216718
rect 641076 216708 641128 216714
rect 641076 216650 641128 216656
rect 642732 216708 642784 216714
rect 642732 216650 642784 216656
rect 640616 216640 640668 216646
rect 640616 216582 640668 216588
rect 640628 210202 640656 216582
rect 641088 210202 641116 216650
rect 641824 210310 642128 210338
rect 641824 210202 641852 210310
rect 606648 210174 606708 210202
rect 607108 210174 607168 210202
rect 607568 210174 607628 210202
rect 608028 210174 608088 210202
rect 608488 210174 608548 210202
rect 608948 210174 609008 210202
rect 609408 210174 609468 210202
rect 609868 210174 609928 210202
rect 610328 210174 610388 210202
rect 610788 210174 610848 210202
rect 611248 210174 611308 210202
rect 611708 210174 611768 210202
rect 612168 210174 612228 210202
rect 612628 210174 612688 210202
rect 613088 210174 613148 210202
rect 613548 210174 613608 210202
rect 614008 210174 614068 210202
rect 614560 210174 614620 210202
rect 615020 210174 615080 210202
rect 615480 210174 615540 210202
rect 615940 210174 616000 210202
rect 616400 210174 616460 210202
rect 616860 210174 616920 210202
rect 617320 210174 617380 210202
rect 617780 210174 617840 210202
rect 618240 210174 618300 210202
rect 618700 210174 618760 210202
rect 619160 210174 619220 210202
rect 619620 210174 619680 210202
rect 620080 210174 620140 210202
rect 620540 210174 620600 210202
rect 621000 210174 621060 210202
rect 621460 210174 621520 210202
rect 622012 210174 622072 210202
rect 622472 210174 622532 210202
rect 622932 210174 622992 210202
rect 623392 210174 623452 210202
rect 623852 210174 623912 210202
rect 624312 210174 624372 210202
rect 624772 210174 624832 210202
rect 625232 210174 625292 210202
rect 625692 210174 625752 210202
rect 626152 210174 626212 210202
rect 626612 210174 626672 210202
rect 627072 210174 627132 210202
rect 627532 210174 627592 210202
rect 627992 210174 628052 210202
rect 628452 210174 628512 210202
rect 628912 210174 628972 210202
rect 629464 210174 629524 210202
rect 629924 210174 629984 210202
rect 630384 210174 630444 210202
rect 630844 210174 630904 210202
rect 631304 210174 631364 210202
rect 631764 210174 631824 210202
rect 632224 210174 632284 210202
rect 632684 210174 632744 210202
rect 633144 210174 633204 210202
rect 633604 210174 633664 210202
rect 634064 210174 634124 210202
rect 634524 210174 634584 210202
rect 634984 210174 635044 210202
rect 635444 210174 635504 210202
rect 635904 210174 635964 210202
rect 636364 210174 636424 210202
rect 636916 210174 636976 210202
rect 637376 210174 637436 210202
rect 637836 210174 637896 210202
rect 638296 210174 638356 210202
rect 638756 210174 638816 210202
rect 639676 210174 639736 210202
rect 640136 210174 640196 210202
rect 640596 210174 640656 210202
rect 641056 210174 641116 210202
rect 641516 210174 641852 210202
rect 642100 210066 642128 210310
rect 642744 210202 642772 216650
rect 643204 210310 643508 210338
rect 643204 210202 643232 210310
rect 642436 210188 642772 210202
rect 642422 210174 642772 210188
rect 642896 210174 643232 210202
rect 642422 210066 642450 210174
rect 642100 210052 642450 210066
rect 643480 210066 643508 210310
rect 644124 210202 644152 217874
rect 645584 216300 645636 216306
rect 645584 216242 645636 216248
rect 644676 210310 644980 210338
rect 644676 210202 644704 210310
rect 643816 210188 644152 210202
rect 643802 210174 644152 210188
rect 644368 210174 644704 210202
rect 643802 210066 643830 210174
rect 643480 210052 643830 210066
rect 644952 210066 644980 210310
rect 645596 210202 645624 216242
rect 646056 210310 646360 210338
rect 646056 210202 646084 210310
rect 645288 210188 645624 210202
rect 645274 210174 645624 210188
rect 645748 210174 646084 210202
rect 645274 210066 645302 210174
rect 644952 210052 645302 210066
rect 646332 210066 646360 210310
rect 646976 210202 647004 217942
rect 647160 210202 647188 220322
rect 649908 220312 649960 220318
rect 649908 220254 649960 220260
rect 648528 220244 648580 220250
rect 648528 220186 648580 220192
rect 647436 210310 647740 210338
rect 647436 210202 647464 210310
rect 646668 210188 647004 210202
rect 646654 210174 647004 210188
rect 647128 210174 647464 210202
rect 646654 210066 646682 210174
rect 646332 210052 646682 210066
rect 647712 210066 647740 210310
rect 648540 210202 648568 220186
rect 648816 210310 649120 210338
rect 648816 210202 648844 210310
rect 648508 210174 648844 210202
rect 649092 210066 649120 210310
rect 649920 210202 649948 220254
rect 651288 220176 651340 220182
rect 651288 220118 651340 220124
rect 651300 212498 651328 220118
rect 651392 216714 651420 987498
rect 652852 987488 652904 987494
rect 652852 987430 652904 987436
rect 652668 987420 652720 987426
rect 652668 987362 652720 987368
rect 651564 987216 651616 987222
rect 651564 987158 651616 987164
rect 651472 986944 651524 986950
rect 651472 986886 651524 986892
rect 651484 218006 651512 986886
rect 651472 218000 651524 218006
rect 651472 217942 651524 217948
rect 651576 217938 651604 987158
rect 651656 987012 651708 987018
rect 651656 986954 651708 986960
rect 651564 217932 651616 217938
rect 651564 217874 651616 217880
rect 651380 216708 651432 216714
rect 651380 216650 651432 216656
rect 651668 216306 651696 986954
rect 652680 220182 652708 987362
rect 652760 987284 652812 987290
rect 652760 987226 652812 987232
rect 652772 222034 652800 987226
rect 652864 222222 652892 987430
rect 658280 987148 658332 987154
rect 658280 987090 658332 987096
rect 658188 987080 658240 987086
rect 658188 987022 658240 987028
rect 652944 984564 652996 984570
rect 652944 984506 652996 984512
rect 652956 266354 652984 984506
rect 655428 984292 655480 984298
rect 655428 984234 655480 984240
rect 654690 922720 654746 922729
rect 654690 922655 654746 922664
rect 654704 922282 654732 922655
rect 654692 922276 654744 922282
rect 654692 922218 654744 922224
rect 654874 909528 654930 909537
rect 654874 909463 654930 909472
rect 654888 908138 654916 909463
rect 654876 908132 654928 908138
rect 654876 908074 654928 908080
rect 654690 896200 654746 896209
rect 654690 896135 654746 896144
rect 654704 895422 654732 896135
rect 654692 895416 654744 895422
rect 654692 895358 654744 895364
rect 655150 882872 655206 882881
rect 655150 882807 655206 882816
rect 655164 870806 655192 882807
rect 655152 870800 655204 870806
rect 655152 870742 655204 870748
rect 655242 856352 655298 856361
rect 655242 856287 655298 856296
rect 655256 855642 655284 856287
rect 655244 855636 655296 855642
rect 655244 855578 655296 855584
rect 654874 843024 654930 843033
rect 654874 842959 654930 842968
rect 654888 841838 654916 842959
rect 654876 841832 654928 841838
rect 654876 841774 654928 841780
rect 655058 816504 655114 816513
rect 655058 816439 655114 816448
rect 655072 815658 655100 816439
rect 655060 815652 655112 815658
rect 655060 815594 655112 815600
rect 655058 789984 655114 789993
rect 655058 789919 655114 789928
rect 655072 789410 655100 789919
rect 655060 789404 655112 789410
rect 655060 789346 655112 789352
rect 654690 763328 654746 763337
rect 654690 763263 654746 763272
rect 654704 761802 654732 763263
rect 654692 761796 654744 761802
rect 654692 761738 654744 761744
rect 654690 750136 654746 750145
rect 654690 750071 654746 750080
rect 654704 749018 654732 750071
rect 654692 749012 654744 749018
rect 654692 748954 654744 748960
rect 654138 736808 654194 736817
rect 654138 736743 654194 736752
rect 654152 736302 654180 736743
rect 654140 736296 654192 736302
rect 654140 736238 654192 736244
rect 654874 696960 654930 696969
rect 654874 696895 654930 696904
rect 654888 696454 654916 696895
rect 654876 696448 654928 696454
rect 654876 696390 654928 696396
rect 654138 683632 654194 683641
rect 654138 683567 654194 683576
rect 654152 683466 654180 683567
rect 654140 683460 654192 683466
rect 654140 683402 654192 683408
rect 654874 643784 654930 643793
rect 654874 643719 654930 643728
rect 654888 643142 654916 643719
rect 654876 643136 654928 643142
rect 654876 643078 654928 643084
rect 654138 630592 654194 630601
rect 654138 630527 654194 630536
rect 654152 629338 654180 630527
rect 654140 629332 654192 629338
rect 654140 629274 654192 629280
rect 654598 617264 654654 617273
rect 654598 617199 654654 617208
rect 654322 603936 654378 603945
rect 654322 603871 654378 603880
rect 654336 602206 654364 603871
rect 654612 603090 654640 617199
rect 654600 603084 654652 603090
rect 654600 603026 654652 603032
rect 654324 602200 654376 602206
rect 654324 602142 654376 602148
rect 654506 577416 654562 577425
rect 654506 577351 654562 577360
rect 654520 576910 654548 577351
rect 654508 576904 654560 576910
rect 654508 576846 654560 576852
rect 654322 564088 654378 564097
rect 654322 564023 654378 564032
rect 654336 556170 654364 564023
rect 654324 556164 654376 556170
rect 654324 556106 654376 556112
rect 655058 550896 655114 550905
rect 655058 550831 655114 550840
rect 655072 550254 655100 550831
rect 655060 550248 655112 550254
rect 655060 550190 655112 550196
rect 654690 537568 654746 537577
rect 654690 537503 654746 537512
rect 654704 536450 654732 537503
rect 654692 536444 654744 536450
rect 654692 536386 654744 536392
rect 654138 524240 654194 524249
rect 654138 524175 654194 524184
rect 654152 522510 654180 524175
rect 654140 522504 654192 522510
rect 654140 522446 654192 522452
rect 654782 511048 654838 511057
rect 654782 510983 654838 510992
rect 654796 510678 654824 510983
rect 654784 510672 654836 510678
rect 654784 510614 654836 510620
rect 655058 484392 655114 484401
rect 655058 484327 655114 484336
rect 655072 483342 655100 484327
rect 655060 483336 655112 483342
rect 655060 483278 655112 483284
rect 654874 471200 654930 471209
rect 654874 471135 654930 471144
rect 654888 470558 654916 471135
rect 654876 470552 654928 470558
rect 654876 470494 654928 470500
rect 654138 457872 654194 457881
rect 654138 457807 654194 457816
rect 654152 457366 654180 457807
rect 654140 457360 654192 457366
rect 654140 457302 654192 457308
rect 654874 431352 654930 431361
rect 654874 431287 654930 431296
rect 654888 430642 654916 431287
rect 654876 430636 654928 430642
rect 654876 430578 654928 430584
rect 655058 418024 655114 418033
rect 655058 417959 655114 417968
rect 655072 417518 655100 417959
rect 655060 417512 655112 417518
rect 655060 417454 655112 417460
rect 654874 404696 654930 404705
rect 654874 404631 654930 404640
rect 654888 404054 654916 404631
rect 654876 404048 654928 404054
rect 654876 403990 654928 403996
rect 654138 391504 654194 391513
rect 654138 391439 654194 391448
rect 654152 389842 654180 391439
rect 654140 389836 654192 389842
rect 654140 389778 654192 389784
rect 654874 351656 654930 351665
rect 654874 351591 654930 351600
rect 654888 350606 654916 351591
rect 654876 350600 654928 350606
rect 654876 350542 654928 350548
rect 654322 338328 654378 338337
rect 654322 338263 654378 338272
rect 654336 336870 654364 338263
rect 654324 336864 654376 336870
rect 654324 336806 654376 336812
rect 654322 325000 654378 325009
rect 654322 324935 654378 324944
rect 654336 323950 654364 324935
rect 654324 323944 654376 323950
rect 654324 323886 654376 323892
rect 654138 311808 654194 311817
rect 654138 311743 654194 311752
rect 654152 311710 654180 311743
rect 654140 311704 654192 311710
rect 654140 311646 654192 311652
rect 655440 310486 655468 984234
rect 655518 975896 655574 975905
rect 655518 975831 655574 975840
rect 655532 938602 655560 975831
rect 655702 962568 655758 962577
rect 655702 962503 655758 962512
rect 655612 960560 655664 960566
rect 655612 960502 655664 960508
rect 655520 938596 655572 938602
rect 655520 938538 655572 938544
rect 655624 936193 655652 960502
rect 655716 938738 655744 962503
rect 655794 949376 655850 949385
rect 655794 949311 655850 949320
rect 655808 938874 655836 949311
rect 655796 938868 655848 938874
rect 655796 938810 655848 938816
rect 655704 938732 655756 938738
rect 655704 938674 655756 938680
rect 655610 936184 655666 936193
rect 655610 936119 655666 936128
rect 656806 869680 656862 869689
rect 656806 869615 656808 869624
rect 656860 869615 656862 869624
rect 656808 869586 656860 869592
rect 655518 829832 655574 829841
rect 655518 829767 655574 829776
rect 655532 782474 655560 829767
rect 656162 803312 656218 803321
rect 656162 803247 656164 803256
rect 656216 803247 656218 803256
rect 656164 803218 656216 803224
rect 655520 782468 655572 782474
rect 655520 782410 655572 782416
rect 655518 776656 655574 776665
rect 655518 776591 655574 776600
rect 655532 738342 655560 776591
rect 655520 738336 655572 738342
rect 655520 738278 655572 738284
rect 655518 723480 655574 723489
rect 655518 723415 655574 723424
rect 655532 691422 655560 723415
rect 655978 710288 656034 710297
rect 655978 710223 656034 710232
rect 655992 709782 656020 710223
rect 655980 709776 656032 709782
rect 655980 709718 656032 709724
rect 655520 691416 655572 691422
rect 655520 691358 655572 691364
rect 655518 670440 655574 670449
rect 655518 670375 655574 670384
rect 655532 647222 655560 670375
rect 656806 657112 656862 657121
rect 656806 657047 656808 657056
rect 656860 657047 656862 657056
rect 656808 657018 656860 657024
rect 655520 647216 655572 647222
rect 655520 647158 655572 647164
rect 656806 590744 656862 590753
rect 656806 590679 656808 590688
rect 656860 590679 656862 590688
rect 656808 590650 656860 590656
rect 656806 497720 656862 497729
rect 656806 497655 656808 497664
rect 656860 497655 656862 497664
rect 656808 497626 656860 497632
rect 656806 444544 656862 444553
rect 656806 444479 656808 444488
rect 656860 444479 656862 444488
rect 656808 444450 656860 444456
rect 656808 378208 656860 378214
rect 656806 378176 656808 378185
rect 656860 378176 656862 378185
rect 656806 378111 656862 378120
rect 656806 364848 656862 364857
rect 656806 364783 656862 364792
rect 656820 364410 656848 364783
rect 656808 364404 656860 364410
rect 656808 364346 656860 364352
rect 655428 310480 655480 310486
rect 655428 310422 655480 310428
rect 656806 298480 656862 298489
rect 656806 298415 656808 298424
rect 656860 298415 656862 298424
rect 656808 298386 656860 298392
rect 655702 285288 655758 285297
rect 655702 285223 655758 285232
rect 655716 284782 655744 285223
rect 655704 284776 655756 284782
rect 655704 284718 655756 284724
rect 652944 266348 652996 266354
rect 652944 266290 652996 266296
rect 658200 262449 658228 987022
rect 658292 264994 658320 987090
rect 658464 984224 658516 984230
rect 658464 984166 658516 984172
rect 658372 984156 658424 984162
rect 658372 984098 658424 984104
rect 658384 311846 658412 984098
rect 658476 314634 658504 984166
rect 663800 908132 663852 908138
rect 663800 908074 663852 908080
rect 660948 895416 661000 895422
rect 660948 895358 661000 895364
rect 660960 759354 660988 895358
rect 663708 869644 663760 869650
rect 663708 869586 663760 869592
rect 661040 803276 661092 803282
rect 661040 803218 661092 803224
rect 660948 759348 661000 759354
rect 660948 759290 661000 759296
rect 660948 709776 661000 709782
rect 660948 709718 661000 709724
rect 660960 579834 660988 709718
rect 661052 670818 661080 803218
rect 661132 736296 661184 736302
rect 661132 736238 661184 736244
rect 661040 670812 661092 670818
rect 661040 670754 661092 670760
rect 661144 623898 661172 736238
rect 663720 716174 663748 869586
rect 663812 759490 663840 908074
rect 666468 855636 666520 855642
rect 666468 855578 666520 855584
rect 663892 789404 663944 789410
rect 663892 789346 663944 789352
rect 663800 759484 663852 759490
rect 663800 759426 663852 759432
rect 663708 716168 663760 716174
rect 663708 716110 663760 716116
rect 663800 696448 663852 696454
rect 663800 696390 663852 696396
rect 663708 657076 663760 657082
rect 663708 657018 663760 657024
rect 661132 623892 661184 623898
rect 661132 623834 661184 623840
rect 661040 602200 661092 602206
rect 661040 602142 661092 602148
rect 660948 579828 661000 579834
rect 660948 579770 661000 579776
rect 661052 491434 661080 602142
rect 663720 535634 663748 657018
rect 663812 579970 663840 696390
rect 663904 670614 663932 789346
rect 666480 716582 666508 855578
rect 666468 716576 666520 716582
rect 666468 716518 666520 716524
rect 663892 670608 663944 670614
rect 663892 670550 663944 670556
rect 666468 643136 666520 643142
rect 666468 643078 666520 643084
rect 663800 579964 663852 579970
rect 663800 579906 663852 579912
rect 663892 576904 663944 576910
rect 663892 576846 663944 576852
rect 663708 535628 663760 535634
rect 663708 535570 663760 535576
rect 661224 522504 661276 522510
rect 661224 522446 661276 522452
rect 661040 491428 661092 491434
rect 661040 491370 661092 491376
rect 661040 457360 661092 457366
rect 661040 457302 661092 457308
rect 660948 417512 661000 417518
rect 660948 417454 661000 417460
rect 658464 314628 658516 314634
rect 658464 314570 658516 314576
rect 658372 311840 658424 311846
rect 658372 311782 658424 311788
rect 660960 267782 660988 417454
rect 661052 312050 661080 457302
rect 661132 404048 661184 404054
rect 661132 403990 661184 403996
rect 661040 312044 661092 312050
rect 661040 311986 661092 311992
rect 661144 267986 661172 403990
rect 661236 403170 661264 522446
rect 663800 497684 663852 497690
rect 663800 497626 663852 497632
rect 663708 470552 663760 470558
rect 663708 470494 663760 470500
rect 661224 403164 661276 403170
rect 661224 403106 661276 403112
rect 663720 313342 663748 470494
rect 663812 356250 663840 497626
rect 663904 491570 663932 576846
rect 666480 535770 666508 643078
rect 666468 535764 666520 535770
rect 666468 535706 666520 535712
rect 663892 491564 663944 491570
rect 663892 491506 663944 491512
rect 663892 444508 663944 444514
rect 663892 444450 663944 444456
rect 663800 356244 663852 356250
rect 663800 356186 663852 356192
rect 663708 313336 663760 313342
rect 663708 313278 663760 313284
rect 663904 312934 663932 444450
rect 666468 430636 666520 430642
rect 666468 430578 666520 430584
rect 663892 312928 663944 312934
rect 663892 312870 663944 312876
rect 666480 268122 666508 430578
rect 666468 268116 666520 268122
rect 666468 268058 666520 268064
rect 661132 267980 661184 267986
rect 661132 267922 661184 267928
rect 660948 267776 661000 267782
rect 660948 267718 661000 267724
rect 658280 264988 658332 264994
rect 658280 264930 658332 264936
rect 658186 262440 658242 262449
rect 658186 262375 658242 262384
rect 662880 230512 662932 230518
rect 662880 230454 662932 230460
rect 662788 230444 662840 230450
rect 662788 230386 662840 230392
rect 652852 222216 652904 222222
rect 652852 222158 652904 222164
rect 652772 222006 652892 222034
rect 652668 220176 652720 220182
rect 652668 220118 652720 220124
rect 652864 220114 652892 222006
rect 652760 220108 652812 220114
rect 652760 220050 652812 220056
rect 652852 220108 652904 220114
rect 652852 220050 652904 220056
rect 651656 216300 651708 216306
rect 651656 216242 651708 216248
rect 651288 212492 651340 212498
rect 651288 212434 651340 212440
rect 651380 212492 651432 212498
rect 651380 212434 651432 212440
rect 651392 210338 651420 212434
rect 650196 210310 650500 210338
rect 650196 210202 650224 210310
rect 649888 210174 650224 210202
rect 650472 210066 650500 210310
rect 651392 210310 651972 210338
rect 651392 210202 651420 210310
rect 651268 210174 651420 210202
rect 651944 210066 651972 210310
rect 652772 210202 652800 220050
rect 655520 220040 655572 220046
rect 655520 219982 655572 219988
rect 654140 219972 654192 219978
rect 654140 219914 654192 219920
rect 653048 210310 653352 210338
rect 653048 210202 653076 210310
rect 652740 210174 653076 210202
rect 653324 210066 653352 210310
rect 654152 210202 654180 219914
rect 654428 210310 654732 210338
rect 654428 210202 654456 210310
rect 654120 210174 654456 210202
rect 654704 210066 654732 210310
rect 655532 210202 655560 219982
rect 656900 219904 656952 219910
rect 656900 219846 656952 219852
rect 655808 210310 656112 210338
rect 655808 210202 655836 210310
rect 655500 210174 655836 210202
rect 656084 210066 656112 210310
rect 656912 210202 656940 219846
rect 658280 219836 658332 219842
rect 658280 219778 658332 219784
rect 657188 210310 657492 210338
rect 657188 210202 657216 210310
rect 656880 210174 657216 210202
rect 657464 210066 657492 210310
rect 658292 210202 658320 219778
rect 659752 219768 659804 219774
rect 659752 219710 659804 219716
rect 658568 210310 658872 210338
rect 658568 210202 658596 210310
rect 658260 210174 658596 210202
rect 658844 210066 658872 210310
rect 659764 210202 659792 219710
rect 661132 219700 661184 219706
rect 661132 219642 661184 219648
rect 660040 210310 660344 210338
rect 660040 210202 660068 210310
rect 659732 210174 660068 210202
rect 660316 210066 660344 210310
rect 661144 210202 661172 219642
rect 662800 218142 662828 230386
rect 662788 218136 662840 218142
rect 662788 218078 662840 218084
rect 662892 210338 662920 230454
rect 663432 219632 663484 219638
rect 663432 219574 663484 219580
rect 662972 218136 663024 218142
rect 662972 218078 663024 218084
rect 661420 210310 661724 210338
rect 661420 210202 661448 210310
rect 661112 210174 661448 210202
rect 661696 210066 661724 210310
rect 662800 210310 662920 210338
rect 662800 210202 662828 210310
rect 662984 210202 663012 218078
rect 663444 210202 663472 219574
rect 664352 219564 664404 219570
rect 664352 219506 664404 219512
rect 663892 219428 663944 219434
rect 663892 219370 663944 219376
rect 663904 210202 663932 219370
rect 664364 210202 664392 219506
rect 664812 219496 664864 219502
rect 664812 219438 664864 219444
rect 664824 210202 664852 219438
rect 665732 215892 665784 215898
rect 665732 215834 665784 215840
rect 665272 215756 665324 215762
rect 665272 215698 665324 215704
rect 665284 210202 665312 215698
rect 665744 210202 665772 215834
rect 666192 215824 666244 215830
rect 666192 215766 666244 215772
rect 666204 210202 666232 215766
rect 662492 210174 662828 210202
rect 662952 210174 663012 210202
rect 663412 210174 663472 210202
rect 663872 210174 663932 210202
rect 664332 210174 664392 210202
rect 664792 210174 664852 210202
rect 665252 210174 665312 210202
rect 665712 210174 665772 210202
rect 666172 210174 666232 210202
rect 642100 210038 642436 210052
rect 643480 210038 643816 210052
rect 644952 210038 645288 210052
rect 646332 210038 646668 210052
rect 647712 210038 648048 210066
rect 649092 210038 649428 210066
rect 650472 210038 650808 210066
rect 651944 210038 652280 210066
rect 653324 210038 653660 210066
rect 654704 210038 655040 210066
rect 656084 210038 656420 210066
rect 657464 210038 657800 210066
rect 658844 210038 659272 210066
rect 660316 210038 660652 210066
rect 661696 210038 662032 210066
rect 600044 209908 600096 209914
rect 600044 209850 600096 209856
rect 599950 208584 600006 208593
rect 599950 208519 600006 208528
rect 599858 207496 599914 207505
rect 599858 207431 599914 207440
rect 600056 206553 600084 209850
rect 601148 207120 601200 207126
rect 601148 207062 601200 207068
rect 600964 207052 601016 207058
rect 600964 206994 601016 207000
rect 600042 206544 600098 206553
rect 600042 206479 600098 206488
rect 599122 205456 599178 205465
rect 599122 205391 599178 205400
rect 600976 204513 601004 206994
rect 600962 204504 601018 204513
rect 600962 204439 601018 204448
rect 582288 204332 582340 204338
rect 582288 204274 582340 204280
rect 599952 204332 600004 204338
rect 599952 204274 600004 204280
rect 581826 204096 581882 204105
rect 581826 204031 581882 204040
rect 581090 202600 581146 202609
rect 581090 202535 581146 202544
rect 581104 201550 581132 202535
rect 581840 201618 581868 204031
rect 599964 202473 599992 204274
rect 601160 203425 601188 207062
rect 601146 203416 601202 203425
rect 601146 203351 601202 203360
rect 599950 202464 600006 202473
rect 599950 202399 600006 202408
rect 581828 201612 581880 201618
rect 581828 201554 581880 201560
rect 599032 201612 599084 201618
rect 599032 201554 599084 201560
rect 581092 201544 581144 201550
rect 581092 201486 581144 201492
rect 599044 201385 599072 201554
rect 599952 201544 600004 201550
rect 599952 201486 600004 201492
rect 599030 201376 599086 201385
rect 599030 201311 599086 201320
rect 581090 201104 581146 201113
rect 581090 201039 581146 201048
rect 581104 200122 581132 201039
rect 599964 200433 599992 201486
rect 599950 200424 600006 200433
rect 599950 200359 600006 200368
rect 581092 200116 581144 200122
rect 581092 200058 581144 200064
rect 599952 200116 600004 200122
rect 599952 200058 600004 200064
rect 582286 199608 582342 199617
rect 582286 199543 582342 199552
rect 582300 198762 582328 199543
rect 599964 199345 599992 200058
rect 599950 199336 600006 199345
rect 599950 199271 600006 199280
rect 582288 198756 582340 198762
rect 582288 198698 582340 198704
rect 599124 198756 599176 198762
rect 599124 198698 599176 198704
rect 599136 198393 599164 198698
rect 599122 198384 599178 198393
rect 599122 198319 599178 198328
rect 581274 197976 581330 197985
rect 581274 197911 581330 197920
rect 580816 197396 580868 197402
rect 580816 197338 580868 197344
rect 580828 196489 580856 197338
rect 581288 197334 581316 197911
rect 599308 197396 599360 197402
rect 599308 197338 599360 197344
rect 581276 197328 581328 197334
rect 599320 197305 599348 197338
rect 599952 197328 600004 197334
rect 581276 197270 581328 197276
rect 599306 197296 599362 197305
rect 599952 197270 600004 197276
rect 599306 197231 599362 197240
rect 580814 196480 580870 196489
rect 580814 196415 580870 196424
rect 599964 196353 599992 197270
rect 599950 196344 600006 196353
rect 599950 196279 600006 196288
rect 599950 195256 600006 195265
rect 599950 195191 600006 195200
rect 582286 194984 582342 194993
rect 582286 194919 582342 194928
rect 582196 194676 582248 194682
rect 582196 194618 582248 194624
rect 582208 193497 582236 194618
rect 582300 194614 582328 194919
rect 599124 194676 599176 194682
rect 599124 194618 599176 194624
rect 582288 194608 582340 194614
rect 582288 194550 582340 194556
rect 599136 194313 599164 194618
rect 599964 194614 599992 195191
rect 599952 194608 600004 194614
rect 599952 194550 600004 194556
rect 599122 194304 599178 194313
rect 599122 194239 599178 194248
rect 582194 193488 582250 193497
rect 582194 193423 582250 193432
rect 599858 193216 599914 193225
rect 599858 193151 599914 193160
rect 582286 191992 582342 192001
rect 582286 191927 582342 191936
rect 582300 191894 582328 191927
rect 599872 191894 599900 193151
rect 599950 192264 600006 192273
rect 599950 192199 600006 192208
rect 582288 191888 582340 191894
rect 582288 191830 582340 191836
rect 599860 191888 599912 191894
rect 599860 191830 599912 191836
rect 599964 191826 599992 192199
rect 581276 191820 581328 191826
rect 581276 191762 581328 191768
rect 599952 191820 600004 191826
rect 599952 191762 600004 191768
rect 581288 190505 581316 191762
rect 599858 191176 599914 191185
rect 599858 191111 599914 191120
rect 581274 190496 581330 190505
rect 579712 190460 579764 190466
rect 599872 190466 599900 191111
rect 581274 190431 581330 190440
rect 599860 190460 599912 190466
rect 579712 190402 579764 190408
rect 599860 190402 599912 190408
rect 579724 188873 579752 190402
rect 600962 190224 601018 190233
rect 600962 190159 601018 190168
rect 579710 188864 579766 188873
rect 579710 188799 579766 188808
rect 582196 187672 582248 187678
rect 582196 187614 582248 187620
rect 582208 185881 582236 187614
rect 600976 187610 601004 190159
rect 601606 189136 601662 189145
rect 601606 189071 601662 189080
rect 601514 188184 601570 188193
rect 601514 188119 601570 188128
rect 582288 187604 582340 187610
rect 582288 187546 582340 187552
rect 600964 187604 601016 187610
rect 600964 187546 601016 187552
rect 582300 187377 582328 187546
rect 582286 187368 582342 187377
rect 582286 187303 582342 187312
rect 599950 187096 600006 187105
rect 599950 187031 600006 187040
rect 582194 185872 582250 185881
rect 582194 185807 582250 185816
rect 599858 185056 599914 185065
rect 599858 184991 599914 185000
rect 580264 184884 580316 184890
rect 580264 184826 580316 184832
rect 580276 182889 580304 184826
rect 580908 184816 580960 184822
rect 580908 184758 580960 184764
rect 580920 184385 580948 184758
rect 580906 184376 580962 184385
rect 580906 184311 580962 184320
rect 599766 184104 599822 184113
rect 599766 184039 599822 184048
rect 580262 182880 580318 182889
rect 580262 182815 580318 182824
rect 581828 182164 581880 182170
rect 581828 182106 581880 182112
rect 580540 182096 580592 182102
rect 580540 182038 580592 182044
rect 580552 181393 580580 182038
rect 580538 181384 580594 181393
rect 580538 181319 580594 181328
rect 581840 179761 581868 182106
rect 581826 179752 581882 179761
rect 581826 179687 581882 179696
rect 580724 179376 580776 179382
rect 580724 179318 580776 179324
rect 580736 176769 580764 179318
rect 599780 179314 599808 184039
rect 599872 182170 599900 184991
rect 599964 184890 599992 187031
rect 600042 186144 600098 186153
rect 600042 186079 600098 186088
rect 599952 184884 600004 184890
rect 599952 184826 600004 184832
rect 599950 183016 600006 183025
rect 599950 182951 600006 182960
rect 599860 182164 599912 182170
rect 599860 182106 599912 182112
rect 599858 182064 599914 182073
rect 599858 181999 599914 182008
rect 581092 179308 581144 179314
rect 581092 179250 581144 179256
rect 599768 179308 599820 179314
rect 599768 179250 599820 179256
rect 581104 178265 581132 179250
rect 599674 178936 599730 178945
rect 599674 178871 599730 178880
rect 581090 178256 581146 178265
rect 581090 178191 581146 178200
rect 598938 176896 598994 176905
rect 598938 176831 598994 176840
rect 580722 176760 580778 176769
rect 598952 176730 598980 176831
rect 580722 176695 580778 176704
rect 581092 176724 581144 176730
rect 581092 176666 581144 176672
rect 598940 176724 598992 176730
rect 598940 176666 598992 176672
rect 580816 173936 580868 173942
rect 580816 173878 580868 173884
rect 579712 173868 579764 173874
rect 579712 173810 579764 173816
rect 579724 172281 579752 173810
rect 579710 172272 579766 172281
rect 579710 172207 579766 172216
rect 579896 171148 579948 171154
rect 579896 171090 579948 171096
rect 579712 168564 579764 168570
rect 579712 168506 579764 168512
rect 579724 158545 579752 168506
rect 579908 161537 579936 171090
rect 580080 171012 580132 171018
rect 580080 170954 580132 170960
rect 580092 169153 580120 170954
rect 580078 169144 580134 169153
rect 580078 169079 580134 169088
rect 580264 168428 580316 168434
rect 580264 168370 580316 168376
rect 580172 168360 580224 168366
rect 580172 168302 580224 168308
rect 580184 166161 580212 168302
rect 580170 166152 580226 166161
rect 580170 166087 580226 166096
rect 580080 165708 580132 165714
rect 580080 165650 580132 165656
rect 579894 161528 579950 161537
rect 579894 161463 579950 161472
rect 579710 158536 579766 158545
rect 579710 158471 579766 158480
rect 580092 152425 580120 165650
rect 580276 155553 580304 168370
rect 580828 164665 580856 173878
rect 580908 171080 580960 171086
rect 580908 171022 580960 171028
rect 580920 170649 580948 171022
rect 580906 170640 580962 170649
rect 580906 170575 580962 170584
rect 581104 167657 581132 176666
rect 581460 176656 581512 176662
rect 581460 176598 581512 176604
rect 581472 175273 581500 176598
rect 581458 175264 581514 175273
rect 581458 175199 581514 175208
rect 582288 173800 582340 173806
rect 582286 173768 582288 173777
rect 582340 173768 582342 173777
rect 582286 173703 582342 173712
rect 582196 171216 582248 171222
rect 582196 171158 582248 171164
rect 581920 168496 581972 168502
rect 581920 168438 581972 168444
rect 581090 167648 581146 167657
rect 581090 167583 581146 167592
rect 581552 165640 581604 165646
rect 581552 165582 581604 165588
rect 580814 164656 580870 164665
rect 580814 164591 580870 164600
rect 581092 162920 581144 162926
rect 581092 162862 581144 162868
rect 580908 157548 580960 157554
rect 580908 157490 580960 157496
rect 580724 157412 580776 157418
rect 580724 157354 580776 157360
rect 580262 155544 580318 155553
rect 580262 155479 580318 155488
rect 580632 154624 580684 154630
rect 580632 154566 580684 154572
rect 580078 152416 580134 152425
rect 580078 152351 580134 152360
rect 579712 143676 579764 143682
rect 579712 143618 579764 143624
rect 579724 122097 579752 143618
rect 579804 143608 579856 143614
rect 579804 143550 579856 143556
rect 579710 122088 579766 122097
rect 579710 122023 579766 122032
rect 579816 119105 579844 143550
rect 580644 138825 580672 154566
rect 580736 143313 580764 157354
rect 580816 151836 580868 151842
rect 580816 151778 580868 151784
rect 580722 143304 580778 143313
rect 580722 143239 580778 143248
rect 580630 138816 580686 138825
rect 580630 138751 580686 138760
rect 579896 138032 579948 138038
rect 579896 137974 579948 137980
rect 579802 119096 579858 119105
rect 579802 119031 579858 119040
rect 579908 112985 579936 137974
rect 580080 135380 580132 135386
rect 580080 135322 580132 135328
rect 579988 132524 580040 132530
rect 579988 132466 580040 132472
rect 579894 112976 579950 112985
rect 579894 112911 579950 112920
rect 580000 105369 580028 132466
rect 580092 108497 580120 135322
rect 580172 135312 580224 135318
rect 580172 135254 580224 135260
rect 580078 108488 580134 108497
rect 580078 108423 580134 108432
rect 580184 106865 580212 135254
rect 580828 134201 580856 151778
rect 580920 137329 580948 157490
rect 581000 157480 581052 157486
rect 581000 157422 581052 157428
rect 581012 141817 581040 157422
rect 581104 147937 581132 162862
rect 581184 160132 581236 160138
rect 581184 160074 581236 160080
rect 581090 147928 581146 147937
rect 581090 147863 581146 147872
rect 581196 144945 581224 160074
rect 581564 150929 581592 165582
rect 581828 165572 581880 165578
rect 581828 165514 581880 165520
rect 581840 163169 581868 165514
rect 581826 163160 581882 163169
rect 581826 163095 581882 163104
rect 581644 162988 581696 162994
rect 581644 162930 581696 162936
rect 581550 150920 581606 150929
rect 581550 150855 581606 150864
rect 581656 149433 581684 162930
rect 581736 160200 581788 160206
rect 581736 160142 581788 160148
rect 581642 149424 581698 149433
rect 581642 149359 581698 149368
rect 581460 149184 581512 149190
rect 581460 149126 581512 149132
rect 581276 146328 581328 146334
rect 581276 146270 581328 146276
rect 581182 144936 581238 144945
rect 581182 144871 581238 144880
rect 580998 141808 581054 141817
rect 580998 141743 581054 141752
rect 581184 140820 581236 140826
rect 581184 140762 581236 140768
rect 581092 138168 581144 138174
rect 581092 138110 581144 138116
rect 581000 138100 581052 138106
rect 581000 138042 581052 138048
rect 580906 137320 580962 137329
rect 580906 137255 580962 137264
rect 580814 134192 580870 134201
rect 580814 134127 580870 134136
rect 580908 132660 580960 132666
rect 580908 132602 580960 132608
rect 580264 132592 580316 132598
rect 580264 132534 580316 132540
rect 580170 106856 580226 106865
rect 580170 106791 580226 106800
rect 579986 105360 580042 105369
rect 579986 105295 580042 105304
rect 580276 103873 580304 132534
rect 580540 129940 580592 129946
rect 580540 129882 580592 129888
rect 580356 129872 580408 129878
rect 580356 129814 580408 129820
rect 580262 103864 580318 103873
rect 580262 103799 580318 103808
rect 580368 97753 580396 129814
rect 580448 129804 580500 129810
rect 580448 129746 580500 129752
rect 580460 100881 580488 129746
rect 580446 100872 580502 100881
rect 580446 100807 580502 100816
rect 580552 99385 580580 129882
rect 580724 127016 580776 127022
rect 580724 126958 580776 126964
rect 580632 124228 580684 124234
rect 580632 124170 580684 124176
rect 580538 99376 580594 99385
rect 580538 99311 580594 99320
rect 580354 97744 580410 97753
rect 580354 97679 580410 97688
rect 580644 91769 580672 124170
rect 580736 96257 580764 126958
rect 580816 124296 580868 124302
rect 580816 124238 580868 124244
rect 580722 96248 580778 96257
rect 580722 96183 580778 96192
rect 580828 93265 580856 124238
rect 580920 102377 580948 132602
rect 581012 111489 581040 138042
rect 580998 111480 581054 111489
rect 580998 111415 581054 111424
rect 581104 109993 581132 138110
rect 581196 114481 581224 140762
rect 581288 123593 581316 146270
rect 581368 140888 581420 140894
rect 581368 140830 581420 140836
rect 581274 123584 581330 123593
rect 581274 123519 581330 123528
rect 581276 116000 581328 116006
rect 581380 115977 581408 140830
rect 581472 125089 581500 149126
rect 581644 149116 581696 149122
rect 581644 149058 581696 149064
rect 581552 140956 581604 140962
rect 581552 140898 581604 140904
rect 581458 125080 581514 125089
rect 581458 125015 581514 125024
rect 581564 117609 581592 140898
rect 581656 126721 581684 149058
rect 581748 146441 581776 160142
rect 581932 157049 581960 168438
rect 582012 160268 582064 160274
rect 582012 160210 582064 160216
rect 581918 157040 581974 157049
rect 581918 156975 581974 156984
rect 581920 151904 581972 151910
rect 581920 151846 581972 151852
rect 581828 149252 581880 149258
rect 581828 149194 581880 149200
rect 581734 146432 581790 146441
rect 581734 146367 581790 146376
rect 581736 143744 581788 143750
rect 581736 143686 581788 143692
rect 581642 126712 581698 126721
rect 581642 126647 581698 126656
rect 581748 120601 581776 143686
rect 581840 129713 581868 149194
rect 581932 131209 581960 151846
rect 582024 140321 582052 160210
rect 582208 160041 582236 171158
rect 599688 171086 599716 178871
rect 599766 177984 599822 177993
rect 599766 177919 599822 177928
rect 599676 171080 599728 171086
rect 599676 171022 599728 171028
rect 599780 171018 599808 177919
rect 599872 176662 599900 181999
rect 599964 179382 599992 182951
rect 600056 182102 600084 186079
rect 601528 184822 601556 188119
rect 601620 187678 601648 189071
rect 601608 187672 601660 187678
rect 601608 187614 601660 187620
rect 601516 184816 601568 184822
rect 601516 184758 601568 184764
rect 600044 182096 600096 182102
rect 600044 182038 600096 182044
rect 600134 180976 600190 180985
rect 600134 180911 600190 180920
rect 600042 180024 600098 180033
rect 600042 179959 600098 179968
rect 599952 179376 600004 179382
rect 599952 179318 600004 179324
rect 599860 176656 599912 176662
rect 599860 176598 599912 176604
rect 599950 174856 600006 174865
rect 599950 174791 600006 174800
rect 599964 173942 599992 174791
rect 599952 173936 600004 173942
rect 599952 173878 600004 173884
rect 600056 173874 600084 179959
rect 600044 173868 600096 173874
rect 600044 173810 600096 173816
rect 600148 173806 600176 180911
rect 600226 175944 600282 175953
rect 600226 175879 600282 175888
rect 600136 173800 600188 173806
rect 600136 173742 600188 173748
rect 599858 172816 599914 172825
rect 599858 172751 599914 172760
rect 599872 171154 599900 172751
rect 599950 171864 600006 171873
rect 599950 171799 600006 171808
rect 599964 171222 599992 171799
rect 599952 171216 600004 171222
rect 599952 171158 600004 171164
rect 599860 171148 599912 171154
rect 599860 171090 599912 171096
rect 599768 171012 599820 171018
rect 599768 170954 599820 170960
rect 598938 170776 598994 170785
rect 598938 170711 598994 170720
rect 598952 168570 598980 170711
rect 599950 169824 600006 169833
rect 599950 169759 600006 169768
rect 599490 168736 599546 168745
rect 599490 168671 599546 168680
rect 598940 168564 598992 168570
rect 598940 168506 598992 168512
rect 599504 168434 599532 168671
rect 599964 168502 599992 169759
rect 599952 168496 600004 168502
rect 599952 168438 600004 168444
rect 599492 168428 599544 168434
rect 599492 168370 599544 168376
rect 600240 168366 600268 175879
rect 601422 173904 601478 173913
rect 601422 173839 601478 173848
rect 600228 168360 600280 168366
rect 600228 168302 600280 168308
rect 599858 167784 599914 167793
rect 599858 167719 599914 167728
rect 599872 165782 599900 167719
rect 600042 166696 600098 166705
rect 600042 166631 600098 166640
rect 582288 165776 582340 165782
rect 582288 165718 582340 165724
rect 599860 165776 599912 165782
rect 599860 165718 599912 165724
rect 599950 165744 600006 165753
rect 582194 160032 582250 160041
rect 582194 159967 582250 159976
rect 582104 154692 582156 154698
rect 582104 154634 582156 154640
rect 582010 140312 582066 140321
rect 582010 140247 582066 140256
rect 582116 135833 582144 154634
rect 582300 154057 582328 165718
rect 600056 165714 600084 166631
rect 599950 165679 600006 165688
rect 600044 165708 600096 165714
rect 599964 165646 599992 165679
rect 600044 165650 600096 165656
rect 599952 165640 600004 165646
rect 599952 165582 600004 165588
rect 601436 165578 601464 173839
rect 601424 165572 601476 165578
rect 601424 165514 601476 165520
rect 599858 164656 599914 164665
rect 599858 164591 599914 164600
rect 599872 162994 599900 164591
rect 599950 163704 600006 163713
rect 599950 163639 600006 163648
rect 599860 162988 599912 162994
rect 599860 162930 599912 162936
rect 599964 162926 599992 163639
rect 599952 162920 600004 162926
rect 599952 162862 600004 162868
rect 600042 162616 600098 162625
rect 600042 162551 600098 162560
rect 599858 161664 599914 161673
rect 599858 161599 599914 161608
rect 599872 160138 599900 161599
rect 599950 160576 600006 160585
rect 599950 160511 600006 160520
rect 599964 160274 599992 160511
rect 599952 160268 600004 160274
rect 599952 160210 600004 160216
rect 600056 160206 600084 162551
rect 600044 160200 600096 160206
rect 600044 160142 600096 160148
rect 599860 160132 599912 160138
rect 599860 160074 599912 160080
rect 600042 159624 600098 159633
rect 600042 159559 600098 159568
rect 599858 158536 599914 158545
rect 599858 158471 599914 158480
rect 599872 157418 599900 158471
rect 599950 157584 600006 157593
rect 599950 157519 599952 157528
rect 600004 157519 600006 157528
rect 599952 157490 600004 157496
rect 600056 157486 600084 159559
rect 600044 157480 600096 157486
rect 600044 157422 600096 157428
rect 599860 157412 599912 157418
rect 599860 157354 599912 157360
rect 599858 156496 599914 156505
rect 599858 156431 599914 156440
rect 599872 154630 599900 156431
rect 599950 155544 600006 155553
rect 599950 155479 600006 155488
rect 599964 154698 599992 155479
rect 599952 154692 600004 154698
rect 599952 154634 600004 154640
rect 599860 154624 599912 154630
rect 599860 154566 599912 154572
rect 600042 154456 600098 154465
rect 600042 154391 600098 154400
rect 582286 154048 582342 154057
rect 582286 153983 582342 153992
rect 599858 153504 599914 153513
rect 599858 153439 599914 153448
rect 599872 151978 599900 153439
rect 599950 152416 600006 152425
rect 599950 152351 600006 152360
rect 582196 151972 582248 151978
rect 582196 151914 582248 151920
rect 599860 151972 599912 151978
rect 599860 151914 599912 151920
rect 582102 135824 582158 135833
rect 582102 135759 582158 135768
rect 582208 132705 582236 151914
rect 599964 151910 599992 152351
rect 599952 151904 600004 151910
rect 599952 151846 600004 151852
rect 600056 151842 600084 154391
rect 600044 151836 600096 151842
rect 600044 151778 600096 151784
rect 598938 151464 598994 151473
rect 598938 151399 598994 151408
rect 598952 149258 598980 151399
rect 599858 150376 599914 150385
rect 599858 150311 599914 150320
rect 598940 149252 598992 149258
rect 598940 149194 598992 149200
rect 599872 149190 599900 150311
rect 599950 149424 600006 149433
rect 599950 149359 600006 149368
rect 599860 149184 599912 149190
rect 599860 149126 599912 149132
rect 599964 149122 599992 149359
rect 599952 149116 600004 149122
rect 599952 149058 600004 149064
rect 599858 148336 599914 148345
rect 599858 148271 599914 148280
rect 599872 146402 599900 148271
rect 599950 147384 600006 147393
rect 599950 147319 600006 147328
rect 582288 146396 582340 146402
rect 582288 146338 582340 146344
rect 599860 146396 599912 146402
rect 599860 146338 599912 146344
rect 582194 132696 582250 132705
rect 582194 132631 582250 132640
rect 581918 131200 581974 131209
rect 581918 131135 581974 131144
rect 581826 129704 581882 129713
rect 581826 129639 581882 129648
rect 582300 128217 582328 146338
rect 599964 146334 599992 147319
rect 599952 146328 600004 146334
rect 599582 146296 599638 146305
rect 599952 146270 600004 146276
rect 599582 146231 599638 146240
rect 599596 143682 599624 146231
rect 599950 145344 600006 145353
rect 599950 145279 600006 145288
rect 599674 144256 599730 144265
rect 599674 144191 599730 144200
rect 599584 143676 599636 143682
rect 599584 143618 599636 143624
rect 599688 143614 599716 144191
rect 599964 143750 599992 145279
rect 599952 143744 600004 143750
rect 599952 143686 600004 143692
rect 599676 143608 599728 143614
rect 599676 143550 599728 143556
rect 599858 143304 599914 143313
rect 599858 143239 599914 143248
rect 599306 141264 599362 141273
rect 599306 141199 599362 141208
rect 599320 140826 599348 141199
rect 599872 140962 599900 143239
rect 599950 142216 600006 142225
rect 599950 142151 600006 142160
rect 599860 140956 599912 140962
rect 599860 140898 599912 140904
rect 599964 140894 599992 142151
rect 599952 140888 600004 140894
rect 599952 140830 600004 140836
rect 599308 140820 599360 140826
rect 599308 140762 599360 140768
rect 600042 140176 600098 140185
rect 600042 140111 600098 140120
rect 599858 139224 599914 139233
rect 599858 139159 599914 139168
rect 599872 138106 599900 139159
rect 599952 138168 600004 138174
rect 599950 138136 599952 138145
rect 600004 138136 600006 138145
rect 599860 138100 599912 138106
rect 599950 138071 600006 138080
rect 599860 138042 599912 138048
rect 600056 138038 600084 140111
rect 600044 138032 600096 138038
rect 600044 137974 600096 137980
rect 599858 137184 599914 137193
rect 599858 137119 599914 137128
rect 599872 135386 599900 137119
rect 599950 136096 600006 136105
rect 599950 136031 600006 136040
rect 599860 135380 599912 135386
rect 599860 135322 599912 135328
rect 599964 135318 599992 136031
rect 599952 135312 600004 135318
rect 599952 135254 600004 135260
rect 599858 135144 599914 135153
rect 599858 135079 599914 135088
rect 599306 133104 599362 133113
rect 599306 133039 599362 133048
rect 599320 132666 599348 133039
rect 599308 132660 599360 132666
rect 599308 132602 599360 132608
rect 599872 132530 599900 135079
rect 599950 134056 600006 134065
rect 599950 133991 600006 134000
rect 599964 132598 599992 133991
rect 599952 132592 600004 132598
rect 599952 132534 600004 132540
rect 599860 132524 599912 132530
rect 599860 132466 599912 132472
rect 598938 132016 598994 132025
rect 598938 131951 598994 131960
rect 598952 129810 598980 131951
rect 599858 131064 599914 131073
rect 599858 130999 599914 131008
rect 599872 129946 599900 130999
rect 599950 129976 600006 129985
rect 599860 129940 599912 129946
rect 599950 129911 600006 129920
rect 599860 129882 599912 129888
rect 599964 129878 599992 129911
rect 599952 129872 600004 129878
rect 599952 129814 600004 129820
rect 598940 129804 598992 129810
rect 598940 129746 598992 129752
rect 599858 129024 599914 129033
rect 599858 128959 599914 128968
rect 582286 128208 582342 128217
rect 582286 128143 582342 128152
rect 582196 127084 582248 127090
rect 582196 127026 582248 127032
rect 582012 124364 582064 124370
rect 582012 124306 582064 124312
rect 581920 121508 581972 121514
rect 581920 121450 581972 121456
rect 581734 120592 581790 120601
rect 581734 120527 581790 120536
rect 581644 118788 581696 118794
rect 581644 118730 581696 118736
rect 581550 117600 581606 117609
rect 581550 117535 581606 117544
rect 581276 115942 581328 115948
rect 581366 115968 581422 115977
rect 581182 114472 581238 114481
rect 581182 114407 581238 114416
rect 581184 110492 581236 110498
rect 581184 110434 581236 110440
rect 581090 109984 581146 109993
rect 581090 109919 581146 109928
rect 581000 107704 581052 107710
rect 581000 107646 581052 107652
rect 580906 102368 580962 102377
rect 580906 102303 580962 102312
rect 580908 99408 580960 99414
rect 580908 99350 580960 99356
rect 580814 93256 580870 93265
rect 580814 93191 580870 93200
rect 580630 91760 580686 91769
rect 580630 91695 580686 91704
rect 578148 85604 578200 85610
rect 578148 85546 578200 85552
rect 576768 55208 576820 55214
rect 576768 55150 576820 55156
rect 571340 53644 571392 53650
rect 571340 53586 571392 53592
rect 84824 52686 85160 52714
rect 52276 47048 52328 47054
rect 52276 46990 52328 46996
rect 85132 45558 85160 52686
rect 150314 52454 150342 52700
rect 215832 52686 216168 52714
rect 281336 52686 281488 52714
rect 150268 52426 150342 52454
rect 150268 48414 150296 52426
rect 212448 51400 212500 51406
rect 212448 51342 212500 51348
rect 149980 48408 150032 48414
rect 149980 48350 150032 48356
rect 150256 48408 150308 48414
rect 150256 48350 150308 48356
rect 149992 47054 150020 48350
rect 149980 47048 150032 47054
rect 149980 46990 150032 46996
rect 141804 46702 142370 46730
rect 85120 45552 85172 45558
rect 85120 45494 85172 45500
rect 52184 42900 52236 42906
rect 52184 42842 52236 42848
rect 141804 41546 141832 46702
rect 209688 43308 209740 43314
rect 209688 43250 209740 43256
rect 194414 42256 194470 42265
rect 194414 42191 194470 42200
rect 194428 42106 194456 42191
rect 194074 42078 194456 42106
rect 187606 41848 187662 41857
rect 187358 41806 187606 41834
rect 187606 41783 187662 41792
rect 209700 41546 209728 43250
rect 141792 41540 141844 41546
rect 141792 41482 141844 41488
rect 207020 41540 207072 41546
rect 207020 41482 207072 41488
rect 209688 41540 209740 41546
rect 209688 41482 209740 41488
rect 141804 40202 141832 41482
rect 141758 40174 141832 40202
rect 141758 39984 141786 40174
rect 207032 17490 207060 41482
rect 212460 41313 212488 51342
rect 215208 48476 215260 48482
rect 215208 48418 215260 48424
rect 215220 47122 215248 48418
rect 216140 48346 216168 52686
rect 230388 51468 230440 51474
rect 230388 51410 230440 51416
rect 218060 48408 218112 48414
rect 218060 48350 218112 48356
rect 216128 48340 216180 48346
rect 216128 48282 216180 48288
rect 213828 47116 213880 47122
rect 213828 47058 213880 47064
rect 215208 47116 215260 47122
rect 215208 47058 215260 47064
rect 209778 41304 209834 41313
rect 209778 41239 209834 41248
rect 212446 41304 212502 41313
rect 212446 41239 212502 41248
rect 209792 17490 209820 41239
rect 213840 24818 213868 47058
rect 215300 42900 215352 42906
rect 215300 42842 215352 42848
rect 213184 24812 213236 24818
rect 213184 24754 213236 24760
rect 213828 24812 213880 24818
rect 213828 24754 213880 24760
rect 213196 17490 213224 24754
rect 207032 17462 207184 17490
rect 209792 17462 210036 17490
rect 212888 17462 213224 17490
rect 215312 17490 215340 42842
rect 218072 41313 218100 48350
rect 226248 43444 226300 43450
rect 226248 43386 226300 43392
rect 223488 43376 223540 43382
rect 223488 43318 223540 43324
rect 218058 41304 218114 41313
rect 218058 41239 218114 41248
rect 218072 33134 218100 41239
rect 218072 33106 218192 33134
rect 218164 17490 218192 33106
rect 223500 22574 223528 43318
rect 226260 23050 226288 43386
rect 224592 23044 224644 23050
rect 224592 22986 224644 22992
rect 226248 23044 226300 23050
rect 226248 22986 226300 22992
rect 221740 22568 221792 22574
rect 221740 22510 221792 22516
rect 223488 22568 223540 22574
rect 223488 22510 223540 22516
rect 221752 17490 221780 22510
rect 224604 17490 224632 22986
rect 215312 17462 215740 17490
rect 218164 17462 218592 17490
rect 221444 17462 221780 17490
rect 224296 17462 224632 17490
rect 230400 6225 230428 51410
rect 281460 48414 281488 52686
rect 346504 52686 346900 52714
rect 412344 52686 412680 52714
rect 477848 52686 478184 52714
rect 346504 48482 346532 52686
rect 346872 52426 346900 52686
rect 346860 52420 346912 52426
rect 346860 52362 346912 52368
rect 412652 48482 412680 52686
rect 478156 48550 478184 52686
rect 543016 52686 543352 52714
rect 478144 48544 478196 48550
rect 478144 48486 478196 48492
rect 526168 48544 526220 48550
rect 526168 48486 526220 48492
rect 346492 48476 346544 48482
rect 346492 48418 346544 48424
rect 412640 48476 412692 48482
rect 412640 48418 412692 48424
rect 494060 48476 494112 48482
rect 494060 48418 494112 48424
rect 281448 48408 281500 48414
rect 281448 48350 281500 48356
rect 494072 46918 494100 48418
rect 506388 48408 506440 48414
rect 506388 48350 506440 48356
rect 494060 46912 494112 46918
rect 494060 46854 494112 46860
rect 502248 46912 502300 46918
rect 502248 46854 502300 46860
rect 460664 45824 460716 45830
rect 460664 45766 460716 45772
rect 367100 45756 367152 45762
rect 367100 45698 367152 45704
rect 312820 45688 312872 45694
rect 312820 45630 312872 45636
rect 230848 45620 230900 45626
rect 230848 45562 230900 45568
rect 230572 43852 230624 43858
rect 230572 43794 230624 43800
rect 230480 43512 230532 43518
rect 230480 43454 230532 43460
rect 230492 10713 230520 43454
rect 230478 10704 230534 10713
rect 230478 10639 230534 10648
rect 230584 7721 230612 43794
rect 230756 43648 230808 43654
rect 230756 43590 230808 43596
rect 230664 43580 230716 43586
rect 230664 43522 230716 43528
rect 230676 9217 230704 43522
rect 230768 13705 230796 43590
rect 230860 16697 230888 45562
rect 312832 44198 312860 45630
rect 367112 44198 367140 45698
rect 312820 44192 312872 44198
rect 312820 44134 312872 44140
rect 367100 44192 367152 44198
rect 367100 44134 367152 44140
rect 310428 44124 310480 44130
rect 310428 44066 310480 44072
rect 365168 44124 365220 44130
rect 365168 44066 365220 44072
rect 444564 44124 444616 44130
rect 444564 44066 444616 44072
rect 231032 43784 231084 43790
rect 231032 43726 231084 43732
rect 230940 43716 230992 43722
rect 230940 43658 230992 43664
rect 230846 16688 230902 16697
rect 230846 16623 230902 16632
rect 230754 13696 230810 13705
rect 230754 13631 230810 13640
rect 230952 12209 230980 43658
rect 231044 15201 231072 43726
rect 310440 42106 310468 44066
rect 365180 42106 365208 44066
rect 419724 43988 419776 43994
rect 419724 43930 419776 43936
rect 405556 43920 405608 43926
rect 405556 43862 405608 43868
rect 310132 42078 310468 42106
rect 364918 42078 365208 42106
rect 405568 42092 405596 43862
rect 419736 42772 419764 43930
rect 415490 41984 415546 41993
rect 415426 41942 415490 41970
rect 415490 41919 415546 41928
rect 307298 41848 307354 41857
rect 307004 41806 307298 41834
rect 362038 41848 362094 41857
rect 361790 41806 362038 41834
rect 307298 41783 307354 41792
rect 416622 41818 416728 41834
rect 416622 41812 416740 41818
rect 416622 41806 416688 41812
rect 362038 41783 362094 41792
rect 416688 41754 416740 41760
rect 420736 41812 420788 41818
rect 420736 41754 420788 41760
rect 420748 38622 420776 41754
rect 444576 38690 444604 44066
rect 460676 42106 460704 45766
rect 475660 45552 475712 45558
rect 475660 45494 475712 45500
rect 474464 44056 474516 44062
rect 474464 43998 474516 44004
rect 474476 42500 474504 43998
rect 460368 42078 460704 42106
rect 470322 41848 470378 41857
rect 470166 41806 470322 41834
rect 471408 41818 471744 41834
rect 471408 41812 471756 41818
rect 471408 41806 471704 41812
rect 470322 41783 470378 41792
rect 471704 41754 471756 41760
rect 475568 41812 475620 41818
rect 475568 41754 475620 41760
rect 444564 38684 444616 38690
rect 444564 38626 444616 38632
rect 475580 38622 475608 41754
rect 420736 38616 420788 38622
rect 420736 38558 420788 38564
rect 475568 38616 475620 38622
rect 475568 38558 475620 38564
rect 475672 38554 475700 45494
rect 502260 41886 502288 46854
rect 506400 41954 506428 48350
rect 518532 48340 518584 48346
rect 518532 48282 518584 48288
rect 507860 42288 507912 42294
rect 507860 42230 507912 42236
rect 506388 41948 506440 41954
rect 506388 41890 506440 41896
rect 502248 41880 502300 41886
rect 502248 41822 502300 41828
rect 507872 38622 507900 42230
rect 518544 42129 518572 48282
rect 524052 45552 524104 45558
rect 524052 45494 524104 45500
rect 518530 42120 518586 42129
rect 518530 42055 518586 42064
rect 521658 42120 521714 42129
rect 521714 42078 521870 42106
rect 521658 42055 521714 42064
rect 524064 41993 524092 45494
rect 526180 42092 526208 48486
rect 543016 47258 543044 52686
rect 559472 51060 559524 51066
rect 559472 51002 559524 51008
rect 535460 47252 535512 47258
rect 535460 47194 535512 47200
rect 543004 47252 543056 47258
rect 543004 47194 543056 47200
rect 530676 42288 530728 42294
rect 531044 42288 531096 42294
rect 530728 42236 531044 42242
rect 530676 42230 531096 42236
rect 530688 42214 531084 42230
rect 535472 41993 535500 47194
rect 559484 45558 559512 51002
rect 565820 49700 565872 49706
rect 565820 49642 565872 49648
rect 559472 45552 559524 45558
rect 559472 45494 559524 45500
rect 565832 44282 565860 49642
rect 565740 44254 565860 44282
rect 565740 42294 565768 44254
rect 571352 44198 571380 53586
rect 576780 44198 576808 55150
rect 565820 44192 565872 44198
rect 565820 44134 565872 44140
rect 571340 44192 571392 44198
rect 571340 44134 571392 44140
rect 576768 44192 576820 44198
rect 576768 44134 576820 44140
rect 565728 42288 565780 42294
rect 565728 42230 565780 42236
rect 524050 41984 524106 41993
rect 520384 41954 520674 41970
rect 520372 41948 520674 41954
rect 520424 41942 520674 41948
rect 529662 41984 529718 41993
rect 529322 41942 529662 41970
rect 524050 41919 524106 41928
rect 529662 41919 529718 41928
rect 535458 41984 535514 41993
rect 535458 41919 535514 41928
rect 520372 41890 520424 41896
rect 518532 41880 518584 41886
rect 514864 41818 515154 41834
rect 518584 41828 518834 41834
rect 518532 41822 518834 41828
rect 514024 41812 514076 41818
rect 514024 41754 514076 41760
rect 514852 41812 515154 41818
rect 514904 41806 515154 41812
rect 518544 41806 518834 41822
rect 514852 41754 514904 41760
rect 507860 38616 507912 38622
rect 507860 38558 507912 38564
rect 514036 38554 514064 41754
rect 565832 41585 565860 44134
rect 578160 43994 578188 85546
rect 579620 82680 579672 82686
rect 579618 82648 579620 82657
rect 579672 82648 579674 82657
rect 579618 82583 579674 82592
rect 580816 81524 580868 81530
rect 580816 81466 580868 81472
rect 578240 75812 578292 75818
rect 578240 75754 578292 75760
rect 578252 51066 578280 75754
rect 578332 69080 578384 69086
rect 578332 69022 578384 69028
rect 578240 51060 578292 51066
rect 578240 51002 578292 51008
rect 578344 49774 578372 69022
rect 580724 66020 580776 66026
rect 580724 65962 580776 65968
rect 580736 65929 580764 65962
rect 580722 65920 580778 65929
rect 580722 65855 580778 65864
rect 580828 64433 580856 81466
rect 580814 64424 580870 64433
rect 580814 64359 580870 64368
rect 579620 59900 579672 59906
rect 579620 59842 579672 59848
rect 579632 59809 579660 59842
rect 579618 59800 579674 59809
rect 579618 59735 579674 59744
rect 579804 59084 579856 59090
rect 579804 59026 579856 59032
rect 579620 58676 579672 58682
rect 579620 58618 579672 58624
rect 579632 58313 579660 58618
rect 579618 58304 579674 58313
rect 579618 58239 579674 58248
rect 579816 55282 579844 59026
rect 579804 55276 579856 55282
rect 579804 55218 579856 55224
rect 580920 53825 580948 99350
rect 581012 81410 581040 107646
rect 581092 104916 581144 104922
rect 581092 104858 581144 104864
rect 581104 81530 581132 104858
rect 581092 81524 581144 81530
rect 581092 81466 581144 81472
rect 581012 81382 581132 81410
rect 581000 72208 581052 72214
rect 581000 72150 581052 72156
rect 581012 69086 581040 72150
rect 581000 69080 581052 69086
rect 581000 69022 581052 69028
rect 581104 67425 581132 81382
rect 581196 70417 581224 110434
rect 581288 78033 581316 115942
rect 581366 115903 581422 115912
rect 581368 113280 581420 113286
rect 581368 113222 581420 113228
rect 581274 78024 581330 78033
rect 581274 77959 581330 77968
rect 581380 75041 581408 113222
rect 581552 113212 581604 113218
rect 581552 113154 581604 113160
rect 581460 110560 581512 110566
rect 581460 110502 581512 110508
rect 581366 75032 581422 75041
rect 581366 74967 581422 74976
rect 581472 72049 581500 110502
rect 581564 76537 581592 113154
rect 581656 81161 581684 118730
rect 581828 118720 581880 118726
rect 581828 118662 581880 118668
rect 581736 116068 581788 116074
rect 581736 116010 581788 116016
rect 581642 81152 581698 81161
rect 581642 81087 581698 81096
rect 581748 79529 581776 116010
rect 581840 84153 581868 118662
rect 581932 85649 581960 121450
rect 582024 90273 582052 124306
rect 582104 121576 582156 121582
rect 582104 121518 582156 121524
rect 582010 90264 582066 90273
rect 582010 90199 582066 90208
rect 582116 87145 582144 121518
rect 582208 94761 582236 127026
rect 599872 127022 599900 128959
rect 599950 127936 600006 127945
rect 599950 127871 600006 127880
rect 599964 127090 599992 127871
rect 599952 127084 600004 127090
rect 599952 127026 600004 127032
rect 599860 127016 599912 127022
rect 599860 126958 599912 126964
rect 600042 126984 600098 126993
rect 600042 126919 600098 126928
rect 599858 125896 599914 125905
rect 599858 125831 599914 125840
rect 599872 124234 599900 125831
rect 599950 124944 600006 124953
rect 599950 124879 600006 124888
rect 599964 124370 599992 124879
rect 599952 124364 600004 124370
rect 599952 124306 600004 124312
rect 600056 124302 600084 126919
rect 600044 124296 600096 124302
rect 600044 124238 600096 124244
rect 599860 124228 599912 124234
rect 599860 124170 599912 124176
rect 598938 123856 598994 123865
rect 598938 123791 598994 123800
rect 598952 121650 598980 123791
rect 599858 122904 599914 122913
rect 599858 122839 599914 122848
rect 582288 121644 582340 121650
rect 582288 121586 582340 121592
rect 598940 121644 598992 121650
rect 598940 121586 598992 121592
rect 582194 94752 582250 94761
rect 582194 94687 582250 94696
rect 582300 88641 582328 121586
rect 599872 121582 599900 122839
rect 599950 121816 600006 121825
rect 599950 121751 600006 121760
rect 599860 121576 599912 121582
rect 599860 121518 599912 121524
rect 599964 121514 599992 121751
rect 599952 121508 600004 121514
rect 599952 121450 600004 121456
rect 600042 120864 600098 120873
rect 600042 120799 600098 120808
rect 599858 119776 599914 119785
rect 599858 119711 599914 119720
rect 599872 118862 599900 119711
rect 583668 118856 583720 118862
rect 583668 118798 583720 118804
rect 599860 118856 599912 118862
rect 599860 118798 599912 118804
rect 599950 118824 600006 118833
rect 582286 88632 582342 88641
rect 582286 88567 582342 88576
rect 582102 87136 582158 87145
rect 582102 87071 582158 87080
rect 581918 85640 581974 85649
rect 581918 85575 581974 85584
rect 582288 84448 582340 84454
rect 582288 84390 582340 84396
rect 582012 84380 582064 84386
rect 582012 84322 582064 84328
rect 581920 84176 581972 84182
rect 581826 84144 581882 84153
rect 581920 84118 581972 84124
rect 581826 84079 581882 84088
rect 581734 79520 581790 79529
rect 581734 79455 581790 79464
rect 581550 76528 581606 76537
rect 581550 76463 581606 76472
rect 581458 72040 581514 72049
rect 581458 71975 581514 71984
rect 581182 70408 581238 70417
rect 581182 70343 581238 70352
rect 581090 67416 581146 67425
rect 581090 67351 581146 67360
rect 581932 56817 581960 84118
rect 582024 62937 582052 84322
rect 582196 84312 582248 84318
rect 582196 84254 582248 84260
rect 582104 84244 582156 84250
rect 582104 84186 582156 84192
rect 582010 62928 582066 62937
rect 582010 62863 582066 62872
rect 581918 56808 581974 56817
rect 581918 56743 581974 56752
rect 582116 55321 582144 84186
rect 582208 61305 582236 84254
rect 582300 68921 582328 84390
rect 583680 82686 583708 118798
rect 599950 118759 599952 118768
rect 600004 118759 600006 118768
rect 599952 118730 600004 118736
rect 600056 118726 600084 120799
rect 600044 118720 600096 118726
rect 600044 118662 600096 118668
rect 599858 117736 599914 117745
rect 599858 117671 599914 117680
rect 599872 116074 599900 117671
rect 599950 116784 600006 116793
rect 599950 116719 600006 116728
rect 599860 116068 599912 116074
rect 599860 116010 599912 116016
rect 599964 116006 599992 116719
rect 599952 116000 600004 116006
rect 599952 115942 600004 115948
rect 599858 115696 599914 115705
rect 599858 115631 599914 115640
rect 599872 113218 599900 115631
rect 599950 114744 600006 114753
rect 599950 114679 600006 114688
rect 599964 113286 599992 114679
rect 599952 113280 600004 113286
rect 599952 113222 600004 113228
rect 599860 113212 599912 113218
rect 599860 113154 599912 113160
rect 599950 112704 600006 112713
rect 599950 112639 600006 112648
rect 599766 111616 599822 111625
rect 599766 111551 599822 111560
rect 599780 110498 599808 111551
rect 599964 110566 599992 112639
rect 600226 110664 600282 110673
rect 600226 110599 600282 110608
rect 599952 110560 600004 110566
rect 599952 110502 600004 110508
rect 599768 110492 599820 110498
rect 599768 110434 599820 110440
rect 599950 109576 600006 109585
rect 599950 109511 600006 109520
rect 599964 107710 599992 109511
rect 599952 107704 600004 107710
rect 599952 107646 600004 107652
rect 599950 107536 600006 107545
rect 599950 107471 600006 107480
rect 599964 104922 599992 107471
rect 599952 104916 600004 104922
rect 599952 104858 600004 104864
rect 599950 100464 600006 100473
rect 599950 100399 600006 100408
rect 599964 99414 599992 100399
rect 599952 99408 600004 99414
rect 599952 99350 600004 99356
rect 589188 95260 589240 95266
rect 589188 95202 589240 95208
rect 589200 85610 589228 95202
rect 597468 95124 597520 95130
rect 597468 95066 597520 95072
rect 590660 89684 590712 89690
rect 590660 89626 590712 89632
rect 589188 85604 589240 85610
rect 589188 85546 589240 85552
rect 586428 84652 586480 84658
rect 586428 84594 586480 84600
rect 583852 84584 583904 84590
rect 583852 84526 583904 84532
rect 583760 84516 583812 84522
rect 583760 84458 583812 84464
rect 583668 82680 583720 82686
rect 583668 82622 583720 82628
rect 582286 68912 582342 68921
rect 582286 68847 582342 68856
rect 582194 61296 582250 61305
rect 582194 61231 582250 61240
rect 583772 59906 583800 84458
rect 583760 59900 583812 59906
rect 583760 59842 583812 59848
rect 583864 58682 583892 84526
rect 586440 66026 586468 84594
rect 590672 75818 590700 89626
rect 590660 75812 590712 75818
rect 590660 75754 590712 75760
rect 594708 66292 594760 66298
rect 594708 66234 594760 66240
rect 587900 66224 587952 66230
rect 587900 66166 587952 66172
rect 586428 66020 586480 66026
rect 586428 65962 586480 65968
rect 583852 58676 583904 58682
rect 583852 58618 583904 58624
rect 582102 55312 582158 55321
rect 582102 55247 582158 55256
rect 580906 53816 580962 53825
rect 580906 53751 580962 53760
rect 587912 53718 587940 66166
rect 594340 63776 594392 63782
rect 594340 63718 594392 63724
rect 594352 59090 594380 63718
rect 594340 59084 594392 59090
rect 594340 59026 594392 59032
rect 587900 53712 587952 53718
rect 587900 53654 587952 53660
rect 578332 49768 578384 49774
rect 578332 49710 578384 49716
rect 590660 49768 590712 49774
rect 590660 49710 590712 49716
rect 590672 44198 590700 49710
rect 590752 48340 590804 48346
rect 590752 48282 590804 48288
rect 590660 44192 590712 44198
rect 590660 44134 590712 44140
rect 578148 43988 578200 43994
rect 578148 43930 578200 43936
rect 590764 41721 590792 48282
rect 594720 41857 594748 66234
rect 597480 66230 597508 95066
rect 600240 84454 600268 110599
rect 600318 108624 600374 108633
rect 600318 108559 600374 108568
rect 600332 84658 600360 108559
rect 600410 106584 600466 106593
rect 600410 106519 600466 106528
rect 600320 84652 600372 84658
rect 600320 84594 600372 84600
rect 600228 84448 600280 84454
rect 600228 84390 600280 84396
rect 600424 84386 600452 106519
rect 600594 105496 600650 105505
rect 600594 105431 600650 105440
rect 600502 103456 600558 103465
rect 600502 103391 600558 103400
rect 600516 84590 600544 103391
rect 600504 84584 600556 84590
rect 600504 84526 600556 84532
rect 600412 84380 600464 84386
rect 600412 84322 600464 84328
rect 600608 84318 600636 105431
rect 600686 104544 600742 104553
rect 600686 104479 600742 104488
rect 600700 84522 600728 104479
rect 600870 102504 600926 102513
rect 600870 102439 600926 102448
rect 600778 101416 600834 101425
rect 600778 101351 600834 101360
rect 600688 84516 600740 84522
rect 600688 84458 600740 84464
rect 600596 84312 600648 84318
rect 600596 84254 600648 84260
rect 600792 84250 600820 101351
rect 600780 84244 600832 84250
rect 600780 84186 600832 84192
rect 600884 84182 600912 102439
rect 606404 100014 606740 100042
rect 603540 95668 603592 95674
rect 603540 95610 603592 95616
rect 603552 89690 603580 95610
rect 606404 95606 606432 100014
rect 607370 99770 607398 100028
rect 607324 99742 607398 99770
rect 607692 100014 608028 100042
rect 608244 100014 608672 100042
rect 608980 100014 609316 100042
rect 609960 100014 610388 100042
rect 604460 95600 604512 95606
rect 604460 95542 604512 95548
rect 606392 95600 606444 95606
rect 606392 95542 606444 95548
rect 603540 89684 603592 89690
rect 603540 89626 603592 89632
rect 600872 84176 600924 84182
rect 600872 84118 600924 84124
rect 598940 82816 598992 82822
rect 598940 82758 598992 82764
rect 598952 74610 598980 82758
rect 600320 75404 600372 75410
rect 600320 75346 600372 75352
rect 598860 74582 598980 74610
rect 598860 72214 598888 74582
rect 598848 72208 598900 72214
rect 598848 72150 598900 72156
rect 600332 66298 600360 75346
rect 602620 71800 602672 71806
rect 602620 71742 602672 71748
rect 600320 66292 600372 66298
rect 600320 66234 600372 66240
rect 597468 66224 597520 66230
rect 597468 66166 597520 66172
rect 602632 63578 602660 71742
rect 597560 63572 597612 63578
rect 597560 63514 597612 63520
rect 602620 63572 602672 63578
rect 602620 63514 602672 63520
rect 597572 49774 597600 63514
rect 604472 55554 604500 95542
rect 607220 83836 607272 83842
rect 607220 83778 607272 83784
rect 605748 82884 605800 82890
rect 605748 82826 605800 82832
rect 605760 63782 605788 82826
rect 607232 75410 607260 83778
rect 607220 75404 607272 75410
rect 607220 75346 607272 75352
rect 605748 63776 605800 63782
rect 605748 63718 605800 63724
rect 599124 55548 599176 55554
rect 599124 55490 599176 55496
rect 604460 55548 604512 55554
rect 604460 55490 604512 55496
rect 597560 49768 597612 49774
rect 597560 49710 597612 49716
rect 599136 48346 599164 55490
rect 599124 48340 599176 48346
rect 599124 48282 599176 48288
rect 607324 45762 607352 99742
rect 607496 95600 607548 95606
rect 607496 95542 607548 95548
rect 607312 45756 607364 45762
rect 607312 45698 607364 45704
rect 607508 43926 607536 95542
rect 607692 95130 607720 100014
rect 607680 95124 607732 95130
rect 607680 95066 607732 95072
rect 608244 91094 608272 100014
rect 608980 95606 609008 100014
rect 608968 95600 609020 95606
rect 608968 95542 609020 95548
rect 610256 95600 610308 95606
rect 610256 95542 610308 95548
rect 610164 95532 610216 95538
rect 610164 95474 610216 95480
rect 607600 91066 608272 91094
rect 607600 45694 607628 91066
rect 610176 82958 610204 95474
rect 610164 82952 610216 82958
rect 610164 82894 610216 82900
rect 610268 45830 610296 95542
rect 610360 82890 610388 100014
rect 610452 100014 610604 100042
rect 610912 100014 611248 100042
rect 611556 100014 611892 100042
rect 612200 100014 612536 100042
rect 612936 100014 613180 100042
rect 613580 100014 613916 100042
rect 614560 100014 614896 100042
rect 610452 95674 610480 100014
rect 610440 95668 610492 95674
rect 610440 95610 610492 95616
rect 610912 95266 610940 100014
rect 611556 95606 611584 100014
rect 611544 95600 611596 95606
rect 611544 95542 611596 95548
rect 612200 95538 612228 100014
rect 612832 95600 612884 95606
rect 612832 95542 612884 95548
rect 612188 95532 612240 95538
rect 612188 95474 612240 95480
rect 610900 95260 610952 95266
rect 610900 95202 610952 95208
rect 610348 82884 610400 82890
rect 610348 82826 610400 82832
rect 612844 71806 612872 95542
rect 612936 83842 612964 100014
rect 613580 95606 613608 100014
rect 613568 95600 613620 95606
rect 613568 95542 613620 95548
rect 614868 94994 614896 100014
rect 614960 100014 615204 100042
rect 615848 100014 616184 100042
rect 616492 100014 616828 100042
rect 617136 100014 617472 100042
rect 617780 100014 618116 100042
rect 618424 100014 618760 100042
rect 619068 100014 619404 100042
rect 619712 100014 620048 100042
rect 614856 94988 614908 94994
rect 614856 94930 614908 94936
rect 614960 91730 614988 100014
rect 616156 95402 616184 100014
rect 616800 95810 616828 100014
rect 616788 95804 616840 95810
rect 616788 95746 616840 95752
rect 617444 95538 617472 100014
rect 617432 95532 617484 95538
rect 617432 95474 617484 95480
rect 616144 95396 616196 95402
rect 616144 95338 616196 95344
rect 615408 94988 615460 94994
rect 615408 94930 615460 94936
rect 613016 91724 613068 91730
rect 613016 91666 613068 91672
rect 614948 91724 615000 91730
rect 614948 91666 615000 91672
rect 612924 83836 612976 83842
rect 612924 83778 612976 83784
rect 612832 71800 612884 71806
rect 612832 71742 612884 71748
rect 610256 45824 610308 45830
rect 610256 45766 610308 45772
rect 607588 45688 607640 45694
rect 607588 45630 607640 45636
rect 613028 45626 613056 91666
rect 613016 45620 613068 45626
rect 613016 45562 613068 45568
rect 607496 43920 607548 43926
rect 607496 43862 607548 43868
rect 615420 42974 615448 94930
rect 618088 94586 618116 100014
rect 618260 95600 618312 95606
rect 618260 95542 618312 95548
rect 618076 94580 618128 94586
rect 618076 94522 618128 94528
rect 618272 43858 618300 95542
rect 618732 94790 618760 100014
rect 619376 95674 619404 100014
rect 619364 95668 619416 95674
rect 619364 95610 619416 95616
rect 620020 95470 620048 100014
rect 620112 100014 620448 100042
rect 621092 100014 621336 100042
rect 620112 95606 620140 100014
rect 621204 95736 621256 95742
rect 621204 95678 621256 95684
rect 620100 95600 620152 95606
rect 620100 95542 620152 95548
rect 620008 95464 620060 95470
rect 620008 95406 620060 95412
rect 618720 94784 618772 94790
rect 618720 94726 618772 94732
rect 618260 43852 618312 43858
rect 618260 43794 618312 43800
rect 621216 43722 621244 95678
rect 621204 43716 621256 43722
rect 621204 43658 621256 43664
rect 621308 43586 621336 100014
rect 621400 100014 621736 100042
rect 622044 100014 622380 100042
rect 622504 100014 623024 100042
rect 623332 100014 623668 100042
rect 623976 100014 624312 100042
rect 624620 100014 624956 100042
rect 625600 100014 625936 100042
rect 626244 100014 626488 100042
rect 626980 100014 627316 100042
rect 627624 100014 627960 100042
rect 628268 100014 628328 100042
rect 621296 43580 621348 43586
rect 621296 43522 621348 43528
rect 621400 43518 621428 100014
rect 622044 95742 622072 100014
rect 622032 95736 622084 95742
rect 622032 95678 622084 95684
rect 621480 95600 621532 95606
rect 622504 95588 622532 100014
rect 623228 95804 623280 95810
rect 623228 95746 623280 95752
rect 621480 95542 621532 95548
rect 621584 95560 622532 95588
rect 621492 43790 621520 95542
rect 621480 43784 621532 43790
rect 621480 43726 621532 43732
rect 621584 43654 621612 95560
rect 623136 95532 623188 95538
rect 623136 95474 623188 95480
rect 622308 95464 622360 95470
rect 622308 95406 622360 95412
rect 621940 94580 621992 94586
rect 621940 94522 621992 94528
rect 621952 84153 621980 94522
rect 622320 87009 622348 95406
rect 622492 95396 622544 95402
rect 622492 95338 622544 95344
rect 622504 87961 622532 95338
rect 622490 87952 622546 87961
rect 622490 87887 622546 87896
rect 622306 87000 622362 87009
rect 622306 86935 622362 86944
rect 621938 84144 621994 84153
rect 621938 84079 621994 84088
rect 623148 83201 623176 95474
rect 623240 88913 623268 95746
rect 623332 95606 623360 100014
rect 623412 95668 623464 95674
rect 623412 95610 623464 95616
rect 623320 95600 623372 95606
rect 623320 95542 623372 95548
rect 623320 94784 623372 94790
rect 623320 94726 623372 94732
rect 623226 88904 623282 88913
rect 623226 88839 623282 88848
rect 623332 85105 623360 94726
rect 623424 86057 623452 95610
rect 623780 95600 623832 95606
rect 623780 95542 623832 95548
rect 623792 90681 623820 95542
rect 623778 90672 623834 90681
rect 623778 90607 623834 90616
rect 623976 89729 624004 100014
rect 624620 95606 624648 100014
rect 624608 95600 624660 95606
rect 624608 95542 624660 95548
rect 625908 91633 625936 100014
rect 626460 92585 626488 100014
rect 627288 93537 627316 100014
rect 627932 94489 627960 100014
rect 628300 95985 628328 100014
rect 628760 100014 628912 100042
rect 629556 100014 629708 100042
rect 630200 100014 630628 100042
rect 630844 100014 631180 100042
rect 631488 100014 631824 100042
rect 632132 100014 632468 100042
rect 632776 100014 633112 100042
rect 633512 100014 633848 100042
rect 634156 100014 634492 100042
rect 634800 100014 635136 100042
rect 635444 100014 635780 100042
rect 636088 100014 636332 100042
rect 636732 100014 637068 100042
rect 637376 100014 637528 100042
rect 638020 100014 638356 100042
rect 638664 100014 638908 100042
rect 639308 100014 639644 100042
rect 639952 100014 640104 100042
rect 640688 100014 640932 100042
rect 641332 100014 641668 100042
rect 641976 100014 642312 100042
rect 642620 100014 642680 100042
rect 643264 100014 643508 100042
rect 643908 100014 644244 100042
rect 644552 100014 644796 100042
rect 628286 95976 628342 95985
rect 628286 95911 628342 95920
rect 628760 95826 628788 100014
rect 628728 95798 628788 95826
rect 629680 95826 629708 100014
rect 630600 95826 630628 100014
rect 631152 96082 631180 100014
rect 631140 96076 631192 96082
rect 631140 96018 631192 96024
rect 631796 95946 631824 100014
rect 632440 96082 632468 100014
rect 633084 96626 633112 100014
rect 633072 96620 633124 96626
rect 633072 96562 633124 96568
rect 633820 96558 633848 100014
rect 633808 96552 633860 96558
rect 633808 96494 633860 96500
rect 634464 96490 634492 100014
rect 634452 96484 634504 96490
rect 634452 96426 634504 96432
rect 635108 96082 635136 100014
rect 635280 96620 635332 96626
rect 635280 96562 635332 96568
rect 632106 96076 632158 96082
rect 632106 96018 632158 96024
rect 632428 96076 632480 96082
rect 632428 96018 632480 96024
rect 634406 96076 634458 96082
rect 634406 96018 634458 96024
rect 635096 96076 635148 96082
rect 635096 96018 635148 96024
rect 631784 95940 631836 95946
rect 631784 95882 631836 95888
rect 629680 95798 629832 95826
rect 630600 95798 631028 95826
rect 632118 95812 632146 96018
rect 632980 95940 633032 95946
rect 632980 95882 633032 95888
rect 632992 95826 633020 95882
rect 632992 95798 633328 95826
rect 634418 95812 634446 96018
rect 635292 95826 635320 96562
rect 635752 96422 635780 100014
rect 636304 96626 636332 100014
rect 636292 96620 636344 96626
rect 636292 96562 636344 96568
rect 637040 96558 637068 100014
rect 636384 96552 636436 96558
rect 636384 96494 636436 96500
rect 637028 96552 637080 96558
rect 637028 96494 637080 96500
rect 635740 96416 635792 96422
rect 635740 96358 635792 96364
rect 636396 95826 636424 96494
rect 635292 95798 635628 95826
rect 636396 95798 636732 95826
rect 637500 95742 637528 100014
rect 637580 96484 637632 96490
rect 637580 96426 637632 96432
rect 637592 95826 637620 96426
rect 637592 95798 637928 95826
rect 637488 95736 637540 95742
rect 637488 95678 637540 95684
rect 638328 95606 638356 100014
rect 638880 95878 638908 100014
rect 639006 96076 639058 96082
rect 639006 96018 639058 96024
rect 638868 95872 638920 95878
rect 638868 95814 638920 95820
rect 639018 95812 639046 96018
rect 639616 95810 639644 100014
rect 639880 96416 639932 96422
rect 639880 96358 639932 96364
rect 639892 95826 639920 96358
rect 640076 95946 640104 100014
rect 640064 95940 640116 95946
rect 640064 95882 640116 95888
rect 639604 95804 639656 95810
rect 639892 95798 640228 95826
rect 639604 95746 639656 95752
rect 640904 95742 640932 100014
rect 640984 96620 641036 96626
rect 640984 96562 641036 96568
rect 640996 95826 641024 96562
rect 640996 95798 641332 95826
rect 640524 95736 640576 95742
rect 640522 95704 640524 95713
rect 640892 95736 640944 95742
rect 640576 95704 640578 95713
rect 640892 95678 640944 95684
rect 641640 95674 641668 100014
rect 640522 95639 640578 95648
rect 641628 95668 641680 95674
rect 641628 95610 641680 95616
rect 642284 95606 642312 100014
rect 642364 96552 642416 96558
rect 642364 96494 642416 96500
rect 642376 95826 642404 96494
rect 642376 95798 642528 95826
rect 638316 95600 638368 95606
rect 638316 95542 638368 95548
rect 642272 95600 642324 95606
rect 642272 95542 642324 95548
rect 627918 94480 627974 94489
rect 627918 94415 627974 94424
rect 627274 93528 627330 93537
rect 627274 93463 627330 93472
rect 626446 92576 626502 92585
rect 626446 92511 626502 92520
rect 625894 91624 625950 91633
rect 625894 91559 625950 91568
rect 623962 89720 624018 89729
rect 623962 89655 624018 89664
rect 623410 86048 623466 86057
rect 623410 85983 623466 85992
rect 623318 85096 623374 85105
rect 623318 85031 623374 85040
rect 623134 83192 623190 83201
rect 623134 83127 623190 83136
rect 622306 82240 622362 82249
rect 622306 82175 622362 82184
rect 621572 43648 621624 43654
rect 621572 43590 621624 43596
rect 621388 43512 621440 43518
rect 621388 43454 621440 43460
rect 622320 43382 622348 82175
rect 622490 81424 622546 81433
rect 622490 81359 622546 81368
rect 622504 43450 622532 81359
rect 631520 80974 631856 81002
rect 639308 80974 639368 81002
rect 631520 72010 631548 80974
rect 629300 72004 629352 72010
rect 629300 71946 629352 71952
rect 631508 72004 631560 72010
rect 631508 71946 631560 71952
rect 622492 43444 622544 43450
rect 622492 43386 622544 43392
rect 622308 43376 622360 43382
rect 622308 43318 622360 43324
rect 629312 43314 629340 71946
rect 639340 51406 639368 80974
rect 639328 51400 639380 51406
rect 639328 51342 639380 51348
rect 641258 43616 641314 43625
rect 641258 43551 641314 43560
rect 629300 43308 629352 43314
rect 629300 43250 629352 43256
rect 615408 42968 615460 42974
rect 641168 42968 641220 42974
rect 615408 42910 615460 42916
rect 641166 42936 641168 42945
rect 641220 42936 641222 42945
rect 641166 42871 641222 42880
rect 641272 42265 641300 43551
rect 641258 42256 641314 42265
rect 641258 42191 641314 42200
rect 594706 41848 594762 41857
rect 594706 41783 594762 41792
rect 590750 41712 590806 41721
rect 590750 41647 590806 41656
rect 565818 41576 565874 41585
rect 565818 41511 565874 41520
rect 642652 41313 642680 100014
rect 642824 95668 642876 95674
rect 642824 95610 642876 95616
rect 642732 95532 642784 95538
rect 642732 95474 642784 95480
rect 642744 92721 642772 95474
rect 642730 92712 642786 92721
rect 642730 92647 642786 92656
rect 642836 51474 642864 95610
rect 642916 95600 642968 95606
rect 642916 95542 642968 95548
rect 642928 52426 642956 95542
rect 643480 94246 643508 100014
rect 643560 95260 643612 95266
rect 643560 95202 643612 95208
rect 643468 94240 643520 94246
rect 643468 94182 643520 94188
rect 643572 85270 643600 95202
rect 644216 94110 644244 100014
rect 644204 94104 644256 94110
rect 644204 94046 644256 94052
rect 644768 93906 644796 100014
rect 644860 100014 645196 100042
rect 645840 100014 646176 100042
rect 646484 100014 646820 100042
rect 647220 100014 647556 100042
rect 647864 100014 648108 100042
rect 644860 95266 644888 100014
rect 646044 95940 646096 95946
rect 646044 95882 646096 95888
rect 645952 95804 646004 95810
rect 645952 95746 646004 95752
rect 645860 95736 645912 95742
rect 645860 95678 645912 95684
rect 644848 95260 644900 95266
rect 644848 95202 644900 95208
rect 644756 93900 644808 93906
rect 644756 93842 644808 93848
rect 643560 85264 643612 85270
rect 643560 85206 643612 85212
rect 645872 82249 645900 95678
rect 645964 94874 645992 95746
rect 646056 95010 646084 95882
rect 646148 95198 646176 100014
rect 646228 95872 646280 95878
rect 646228 95814 646280 95820
rect 646136 95192 646188 95198
rect 646136 95134 646188 95140
rect 646056 94982 646176 95010
rect 645964 94846 646084 94874
rect 645952 94784 646004 94790
rect 645952 94726 646004 94732
rect 645964 89729 645992 94726
rect 645950 89720 646006 89729
rect 645950 89655 646006 89664
rect 646056 87145 646084 94846
rect 646042 87136 646098 87145
rect 646042 87071 646098 87080
rect 646148 84697 646176 94982
rect 646240 94790 646268 95814
rect 646792 95334 646820 100014
rect 647528 96082 647556 100014
rect 647516 96076 647568 96082
rect 647516 96018 647568 96024
rect 646780 95328 646832 95334
rect 646780 95270 646832 95276
rect 646688 95124 646740 95130
rect 646688 95066 646740 95072
rect 646228 94784 646280 94790
rect 646228 94726 646280 94732
rect 646700 85202 646728 95066
rect 648080 94518 648108 100014
rect 648172 100014 648508 100042
rect 649152 100014 649396 100042
rect 648172 95130 648200 100014
rect 648160 95124 648212 95130
rect 648160 95066 648212 95072
rect 648896 95124 648948 95130
rect 648896 95066 648948 95072
rect 648712 94852 648764 94858
rect 648712 94794 648764 94800
rect 648068 94512 648120 94518
rect 648068 94454 648120 94460
rect 648724 85338 648752 94794
rect 648804 94716 648856 94722
rect 648804 94658 648856 94664
rect 648816 85406 648844 94658
rect 648908 85542 648936 95066
rect 649368 94042 649396 100014
rect 649460 100014 649796 100042
rect 650104 100014 650440 100042
rect 650748 100014 651084 100042
rect 651728 100014 652064 100042
rect 652372 100014 652708 100042
rect 653016 100014 653352 100042
rect 649460 94722 649488 100014
rect 650104 94858 650132 100014
rect 650748 95130 650776 100014
rect 652036 96490 652064 100014
rect 652024 96484 652076 96490
rect 652024 96426 652076 96432
rect 651472 95260 651524 95266
rect 651472 95202 651524 95208
rect 650736 95124 650788 95130
rect 650736 95066 650788 95072
rect 650092 94852 650144 94858
rect 650092 94794 650144 94800
rect 649448 94716 649500 94722
rect 649448 94658 649500 94664
rect 649356 94036 649408 94042
rect 649356 93978 649408 93984
rect 648896 85536 648948 85542
rect 648896 85478 648948 85484
rect 651484 85474 651512 95202
rect 652680 95130 652708 100014
rect 653220 96076 653272 96082
rect 653220 96018 653272 96024
rect 652668 95124 652720 95130
rect 652668 95066 652720 95072
rect 653232 92585 653260 96018
rect 653324 94722 653352 100014
rect 653416 100014 653752 100042
rect 654396 100014 654732 100042
rect 655040 100014 655376 100042
rect 655684 100014 656020 100042
rect 656328 100014 656664 100042
rect 656972 100014 657308 100042
rect 653416 95266 653444 100014
rect 654704 96558 654732 100014
rect 654692 96552 654744 96558
rect 654692 96494 654744 96500
rect 653404 95260 653456 95266
rect 653404 95202 653456 95208
rect 653312 94716 653364 94722
rect 653312 94658 653364 94664
rect 654048 94104 654100 94110
rect 654048 94046 654100 94052
rect 653496 93900 653548 93906
rect 653496 93842 653548 93848
rect 653218 92576 653274 92585
rect 653218 92511 653274 92520
rect 653508 90681 653536 93842
rect 654060 91497 654088 94046
rect 655348 93401 655376 100014
rect 655992 96626 656020 100014
rect 655980 96620 656032 96626
rect 655980 96562 656032 96568
rect 656636 95402 656664 100014
rect 656992 95600 657044 95606
rect 656992 95542 657044 95548
rect 656624 95396 656676 95402
rect 656624 95338 656676 95344
rect 656900 94580 656952 94586
rect 656900 94522 656952 94528
rect 656912 94042 656940 94522
rect 656900 94036 656952 94042
rect 656900 93978 656952 93984
rect 655334 93392 655390 93401
rect 655334 93327 655390 93336
rect 654046 91488 654102 91497
rect 654046 91423 654102 91432
rect 653494 90672 653550 90681
rect 653494 90607 653550 90616
rect 657004 90409 657032 95542
rect 657084 95260 657136 95266
rect 657084 95202 657136 95208
rect 656990 90400 657046 90409
rect 656990 90335 657046 90344
rect 657096 88874 657124 95202
rect 657280 94654 657308 100014
rect 657372 100014 657616 100042
rect 657924 100014 658260 100042
rect 658904 100014 659148 100042
rect 657372 94761 657400 100014
rect 657728 99816 657780 99822
rect 657728 99758 657780 99764
rect 657740 95132 657768 99758
rect 657924 95266 657952 100014
rect 659120 96558 659148 100014
rect 659212 100014 659548 100042
rect 660284 100014 660620 100042
rect 658280 96552 658332 96558
rect 658280 96494 658332 96500
rect 659108 96552 659160 96558
rect 659108 96494 659160 96500
rect 657912 95260 657964 95266
rect 657912 95202 657964 95208
rect 658292 95132 658320 96494
rect 659212 95606 659240 100014
rect 659568 96620 659620 96626
rect 659568 96562 659620 96568
rect 659200 95600 659252 95606
rect 659200 95542 659252 95548
rect 659580 95132 659608 96562
rect 660592 95538 660620 100014
rect 660914 99822 660942 100028
rect 661572 100014 661908 100042
rect 662216 100014 662276 100042
rect 662860 100014 663288 100042
rect 663504 100014 663656 100042
rect 660902 99816 660954 99822
rect 660902 99758 660954 99764
rect 661880 96626 661908 100014
rect 661868 96620 661920 96626
rect 661868 96562 661920 96568
rect 661960 96484 662012 96490
rect 661960 96426 662012 96432
rect 660580 95532 660632 95538
rect 660580 95474 660632 95480
rect 661408 95532 661460 95538
rect 661408 95474 661460 95480
rect 661420 95132 661448 95474
rect 661972 95132 662000 96426
rect 662248 95577 662276 100014
rect 663064 96620 663116 96626
rect 663064 96562 663116 96568
rect 662512 96552 662564 96558
rect 662512 96494 662564 96500
rect 662234 95568 662290 95577
rect 662234 95503 662290 95512
rect 662524 95132 662552 96494
rect 663076 95132 663104 96562
rect 663156 95396 663208 95402
rect 663156 95338 663208 95344
rect 657358 94752 657414 94761
rect 657358 94687 657414 94696
rect 657268 94648 657320 94654
rect 657268 94590 657320 94596
rect 658568 94586 658858 94602
rect 658556 94580 658858 94586
rect 658608 94574 658858 94580
rect 658556 94522 658608 94528
rect 659844 94512 659896 94518
rect 660396 94512 660448 94518
rect 659896 94460 660146 94466
rect 659844 94454 660146 94460
rect 660448 94460 660698 94466
rect 660396 94454 660698 94460
rect 659856 94438 660146 94454
rect 660408 94438 660698 94454
rect 663168 91066 663196 95338
rect 663260 93809 663288 100014
rect 663340 95328 663392 95334
rect 663340 95270 663392 95276
rect 663246 93800 663302 93809
rect 663246 93735 663302 93744
rect 663352 93129 663380 95270
rect 663432 95192 663484 95198
rect 663432 95134 663484 95140
rect 663338 93120 663394 93129
rect 663338 93055 663394 93064
rect 663444 92313 663472 95134
rect 663524 94648 663576 94654
rect 663524 94590 663576 94596
rect 663430 92304 663486 92313
rect 663430 92239 663486 92248
rect 663246 91080 663302 91089
rect 663168 91038 663246 91066
rect 663246 91015 663302 91024
rect 663536 89593 663564 94590
rect 663522 89584 663578 89593
rect 663522 89519 663578 89528
rect 658016 88874 658306 88890
rect 659488 88874 659594 88890
rect 663628 88874 663656 100014
rect 663800 95124 663852 95130
rect 663800 95066 663852 95072
rect 663708 94716 663760 94722
rect 663708 94658 663760 94664
rect 663720 90409 663748 94658
rect 663706 90400 663762 90409
rect 663706 90335 663762 90344
rect 657084 88868 657136 88874
rect 657084 88810 657136 88816
rect 658004 88868 658306 88874
rect 658056 88862 658306 88868
rect 659476 88868 659594 88874
rect 658004 88810 658056 88816
rect 659528 88862 659594 88868
rect 663616 88868 663668 88874
rect 659476 88810 659528 88816
rect 663616 88810 663668 88816
rect 662142 88768 662198 88777
rect 661986 88726 662142 88754
rect 663812 88754 663840 95066
rect 662538 88726 663840 88754
rect 662142 88703 662198 88712
rect 657188 85542 657216 88196
rect 657176 85536 657228 85542
rect 657176 85478 657228 85484
rect 651472 85468 651524 85474
rect 651472 85410 651524 85416
rect 648804 85400 648856 85406
rect 648804 85342 648856 85348
rect 657740 85338 657768 88196
rect 658844 85474 658872 88196
rect 658832 85468 658884 85474
rect 658832 85410 658884 85416
rect 648712 85332 648764 85338
rect 648712 85274 648764 85280
rect 657728 85332 657780 85338
rect 657728 85274 657780 85280
rect 660132 85270 660160 88196
rect 660684 85406 660712 88196
rect 660672 85400 660724 85406
rect 660672 85342 660724 85348
rect 660120 85264 660172 85270
rect 660120 85206 660172 85212
rect 661420 85202 661448 88196
rect 646688 85196 646740 85202
rect 646688 85138 646740 85144
rect 661408 85196 661460 85202
rect 661408 85138 661460 85144
rect 646134 84688 646190 84697
rect 646134 84623 646190 84632
rect 645858 82240 645914 82249
rect 645858 82175 645914 82184
rect 642916 52420 642968 52426
rect 642916 52362 642968 52368
rect 642824 51468 642876 51474
rect 642824 51410 642876 51416
rect 666572 46918 666600 989402
rect 666652 987828 666704 987834
rect 666652 987770 666704 987776
rect 666664 149054 666692 987770
rect 666928 987760 666980 987766
rect 666928 987702 666980 987708
rect 666744 987624 666796 987630
rect 666744 987566 666796 987572
rect 666756 183938 666784 987566
rect 666836 984904 666888 984910
rect 666836 984846 666888 984852
rect 666744 183932 666796 183938
rect 666744 183874 666796 183880
rect 666742 183832 666798 183841
rect 666742 183767 666798 183776
rect 666756 180441 666784 183767
rect 666742 180432 666798 180441
rect 666742 180367 666798 180376
rect 666742 178800 666798 178809
rect 666742 178735 666798 178744
rect 666756 175409 666784 178735
rect 666848 176662 666876 984846
rect 666940 179382 666968 987702
rect 669228 987692 669280 987698
rect 669228 987634 669280 987640
rect 668768 985380 668820 985386
rect 668768 985322 668820 985328
rect 668676 982932 668728 982938
rect 668676 982874 668728 982880
rect 667112 841832 667164 841838
rect 667112 841774 667164 841780
rect 667020 761796 667072 761802
rect 667020 761738 667072 761744
rect 667032 624034 667060 761738
rect 667124 715766 667152 841774
rect 668584 756424 668636 756430
rect 668584 756366 668636 756372
rect 667112 715760 667164 715766
rect 667112 715702 667164 715708
rect 668596 712910 668624 756366
rect 668584 712904 668636 712910
rect 668584 712846 668636 712852
rect 667204 629332 667256 629338
rect 667204 629274 667256 629280
rect 667020 624028 667072 624034
rect 667020 623970 667072 623976
rect 667112 536444 667164 536450
rect 667112 536386 667164 536392
rect 667020 510672 667072 510678
rect 667020 510614 667072 510620
rect 667032 356386 667060 510614
rect 667124 403306 667152 536386
rect 667216 532914 667244 629274
rect 667204 532908 667256 532914
rect 667204 532850 667256 532856
rect 667112 403300 667164 403306
rect 667112 403242 667164 403248
rect 667112 364404 667164 364410
rect 667112 364346 667164 364352
rect 667020 356380 667072 356386
rect 667020 356322 667072 356328
rect 667020 336864 667072 336870
rect 667020 336806 667072 336812
rect 666928 179376 666980 179382
rect 666928 179318 666980 179324
rect 667032 176866 667060 336806
rect 667124 220998 667152 364346
rect 668596 278186 668624 712846
rect 668688 621625 668716 982874
rect 668780 667321 668808 985322
rect 669134 983376 669190 983385
rect 669134 983311 669190 983320
rect 669044 983000 669096 983006
rect 669044 982942 669096 982948
rect 668952 815652 669004 815658
rect 668952 815594 669004 815600
rect 668860 749012 668912 749018
rect 668860 748954 668912 748960
rect 668766 667312 668822 667321
rect 668766 667247 668822 667256
rect 668872 624170 668900 748954
rect 668964 671022 668992 815594
rect 669056 713250 669084 982942
rect 669044 713244 669096 713250
rect 669044 713186 669096 713192
rect 669148 712502 669176 983311
rect 669136 712496 669188 712502
rect 669136 712438 669188 712444
rect 669136 683460 669188 683466
rect 669136 683402 669188 683408
rect 668952 671016 669004 671022
rect 668952 670958 669004 670964
rect 668860 624164 668912 624170
rect 668860 624106 668912 624112
rect 668674 621616 668730 621625
rect 668674 621551 668730 621560
rect 669044 590708 669096 590714
rect 669044 590650 669096 590656
rect 669056 491706 669084 590650
rect 669148 580106 669176 683402
rect 669136 580100 669188 580106
rect 669136 580042 669188 580048
rect 669136 550248 669188 550254
rect 669136 550190 669188 550196
rect 669044 491700 669096 491706
rect 669044 491642 669096 491648
rect 669148 403442 669176 550190
rect 669136 403436 669188 403442
rect 669136 403378 669188 403384
rect 669136 323944 669188 323950
rect 669136 323886 669188 323892
rect 668584 278180 668636 278186
rect 668584 278122 668636 278128
rect 667112 220992 667164 220998
rect 667112 220934 667164 220940
rect 667112 183932 667164 183938
rect 667112 183874 667164 183880
rect 667020 176860 667072 176866
rect 667020 176802 667072 176808
rect 666836 176656 666888 176662
rect 666836 176598 666888 176604
rect 667124 176594 667152 183874
rect 669148 177002 669176 323886
rect 669136 176996 669188 177002
rect 669136 176938 669188 176944
rect 667112 176588 667164 176594
rect 667112 176530 667164 176536
rect 666742 175400 666798 175409
rect 666742 175335 666798 175344
rect 666742 173632 666798 173641
rect 666742 173567 666798 173576
rect 666756 170241 666784 173567
rect 666742 170232 666798 170241
rect 666742 170167 666798 170176
rect 666742 168600 666798 168609
rect 666742 168535 666798 168544
rect 666756 165209 666784 168535
rect 666742 165200 666798 165209
rect 666742 165135 666798 165144
rect 666742 163568 666798 163577
rect 666742 163503 666798 163512
rect 666756 160177 666784 163503
rect 666742 160168 666798 160177
rect 666742 160103 666798 160112
rect 666742 158400 666798 158409
rect 666742 158335 666798 158344
rect 666756 155009 666784 158335
rect 666742 155000 666798 155009
rect 666742 154935 666798 154944
rect 666742 153368 666798 153377
rect 666742 153303 666798 153312
rect 666756 149977 666784 153303
rect 666742 149968 666798 149977
rect 666742 149903 666798 149912
rect 666664 149026 666784 149054
rect 666650 148200 666706 148209
rect 666650 148135 666706 148144
rect 666664 144945 666692 148135
rect 666650 144936 666706 144945
rect 666650 144871 666706 144880
rect 666650 143168 666706 143177
rect 666650 143103 666706 143112
rect 666664 139777 666692 143103
rect 666650 139768 666706 139777
rect 666650 139703 666706 139712
rect 666650 132968 666706 132977
rect 666650 132903 666706 132912
rect 666664 129577 666692 132903
rect 666756 129810 666784 149026
rect 669240 129878 669268 987634
rect 669504 986876 669556 986882
rect 669504 986818 669556 986824
rect 669412 986808 669464 986814
rect 669412 986750 669464 986756
rect 669320 986740 669372 986746
rect 669320 986682 669372 986688
rect 669332 353394 669360 986682
rect 669424 353530 669452 986750
rect 669516 356114 669544 986818
rect 675668 985584 675720 985590
rect 672722 985552 672778 985561
rect 669596 985516 669648 985522
rect 675668 985526 675720 985532
rect 672722 985487 672778 985496
rect 669596 985458 669648 985464
rect 669608 488578 669636 985458
rect 670424 985448 670476 985454
rect 670424 985390 670476 985396
rect 672538 985416 672594 985425
rect 669686 983240 669742 983249
rect 669686 983175 669742 983184
rect 669596 488572 669648 488578
rect 669596 488514 669648 488520
rect 669700 488102 669728 983175
rect 670238 983104 670294 983113
rect 670238 983039 670294 983048
rect 670054 982968 670110 982977
rect 670054 982903 670110 982912
rect 669872 922276 669924 922282
rect 669872 922218 669924 922224
rect 669884 759626 669912 922218
rect 669872 759620 669924 759626
rect 669872 759562 669924 759568
rect 669778 759248 669834 759257
rect 669778 759183 669834 759192
rect 669688 488096 669740 488102
rect 669688 488038 669740 488044
rect 669596 389836 669648 389842
rect 669596 389778 669648 389784
rect 669504 356108 669556 356114
rect 669504 356050 669556 356056
rect 669412 353524 669464 353530
rect 669412 353466 669464 353472
rect 669320 353388 669372 353394
rect 669320 353330 669372 353336
rect 669412 350600 669464 350606
rect 669412 350542 669464 350548
rect 669320 311704 669372 311710
rect 669320 311646 669372 311652
rect 669332 132666 669360 311646
rect 669424 177138 669452 350542
rect 669504 298444 669556 298450
rect 669504 298386 669556 298392
rect 669412 177132 669464 177138
rect 669412 177074 669464 177080
rect 669516 132802 669544 298386
rect 669608 221066 669636 389778
rect 669688 378208 669740 378214
rect 669688 378150 669740 378156
rect 669700 221202 669728 378150
rect 669792 278050 669820 759183
rect 669964 756356 670016 756362
rect 669964 756298 670016 756304
rect 669872 756288 669924 756294
rect 669872 756230 669924 756236
rect 669884 278390 669912 756230
rect 669872 278384 669924 278390
rect 669872 278326 669924 278332
rect 669976 278118 670004 756298
rect 670068 532846 670096 982903
rect 670148 935740 670200 935746
rect 670148 935682 670200 935688
rect 670160 756294 670188 935682
rect 670148 756288 670200 756294
rect 670148 756230 670200 756236
rect 670252 714950 670280 983039
rect 670332 935808 670384 935814
rect 670332 935750 670384 935756
rect 670344 756362 670372 935750
rect 670332 756356 670384 756362
rect 670332 756298 670384 756304
rect 670240 714944 670292 714950
rect 670240 714886 670292 714892
rect 670148 714876 670200 714882
rect 670148 714818 670200 714824
rect 670056 532840 670108 532846
rect 670056 532782 670108 532788
rect 670056 483336 670108 483342
rect 670056 483278 670108 483284
rect 670068 356522 670096 483278
rect 670056 356516 670108 356522
rect 670056 356458 670108 356464
rect 670056 284776 670108 284782
rect 670056 284718 670108 284724
rect 669964 278112 670016 278118
rect 669964 278054 670016 278060
rect 669780 278044 669832 278050
rect 669780 277986 669832 277992
rect 669688 221196 669740 221202
rect 669688 221138 669740 221144
rect 669596 221060 669648 221066
rect 669596 221002 669648 221008
rect 670068 132938 670096 284718
rect 670160 278322 670188 714818
rect 670252 670342 670280 714886
rect 670332 713652 670384 713658
rect 670332 713594 670384 713600
rect 670240 670336 670292 670342
rect 670240 670278 670292 670284
rect 670240 623824 670292 623830
rect 670240 623766 670292 623772
rect 670252 580242 670280 623766
rect 670240 580236 670292 580242
rect 670240 580178 670292 580184
rect 670148 278316 670200 278322
rect 670148 278258 670200 278264
rect 670344 278254 670372 713594
rect 670436 623830 670464 985390
rect 672538 985351 672594 985360
rect 670976 985176 671028 985182
rect 670976 985118 671028 985124
rect 670884 984972 670936 984978
rect 670884 984914 670936 984920
rect 670792 984632 670844 984638
rect 670792 984574 670844 984580
rect 670700 984360 670752 984366
rect 670700 984302 670752 984308
rect 670516 759076 670568 759082
rect 670516 759018 670568 759024
rect 670528 715290 670556 759018
rect 670608 756492 670660 756498
rect 670608 756434 670660 756440
rect 670516 715284 670568 715290
rect 670516 715226 670568 715232
rect 670528 714882 670556 715226
rect 670516 714876 670568 714882
rect 670516 714818 670568 714824
rect 670620 713658 670648 756434
rect 670608 713652 670660 713658
rect 670608 713594 670660 713600
rect 670608 713244 670660 713250
rect 670608 713186 670660 713192
rect 670516 712496 670568 712502
rect 670516 712438 670568 712444
rect 670528 699786 670556 712438
rect 670516 699780 670568 699786
rect 670516 699722 670568 699728
rect 670620 699666 670648 713186
rect 670528 699638 670648 699666
rect 670528 668710 670556 699638
rect 670608 699576 670660 699582
rect 670608 699518 670660 699524
rect 670516 668704 670568 668710
rect 670516 668646 670568 668652
rect 670620 667758 670648 699518
rect 670608 667752 670660 667758
rect 670608 667694 670660 667700
rect 670608 624300 670660 624306
rect 670608 624242 670660 624248
rect 670424 623824 670476 623830
rect 670424 623766 670476 623772
rect 670516 621104 670568 621110
rect 670516 621046 670568 621052
rect 670424 621036 670476 621042
rect 670424 620978 670476 620984
rect 670436 278526 670464 620978
rect 670528 577182 670556 621046
rect 670516 577176 670568 577182
rect 670516 577118 670568 577124
rect 670424 278520 670476 278526
rect 670424 278462 670476 278468
rect 670528 278458 670556 577118
rect 670620 278594 670648 624242
rect 670608 278588 670660 278594
rect 670608 278530 670660 278536
rect 670516 278452 670568 278458
rect 670516 278394 670568 278400
rect 670332 278248 670384 278254
rect 670332 278190 670384 278196
rect 670712 189009 670740 984302
rect 670804 194041 670832 984574
rect 670896 199073 670924 984914
rect 670988 204241 671016 985118
rect 671988 984836 672040 984842
rect 671988 984778 672040 984784
rect 671068 984768 671120 984774
rect 671068 984710 671120 984716
rect 671080 209273 671108 984710
rect 671804 705492 671856 705498
rect 671804 705434 671856 705440
rect 671160 314628 671212 314634
rect 671160 314570 671212 314576
rect 671172 312118 671200 314570
rect 671160 312112 671212 312118
rect 671160 312054 671212 312060
rect 671160 311840 671212 311846
rect 671160 311782 671212 311788
rect 671172 309670 671200 311782
rect 671160 309664 671212 309670
rect 671160 309606 671212 309612
rect 671160 218068 671212 218074
rect 671160 218010 671212 218016
rect 671066 209264 671122 209273
rect 671066 209199 671122 209208
rect 671080 205873 671108 209199
rect 671066 205864 671122 205873
rect 671066 205799 671122 205808
rect 670974 204232 671030 204241
rect 670974 204167 671030 204176
rect 670988 200841 671016 204167
rect 670974 200832 671030 200841
rect 670974 200767 671030 200776
rect 670882 199064 670938 199073
rect 670882 198999 670938 199008
rect 670896 195673 670924 198999
rect 670882 195664 670938 195673
rect 670882 195599 670938 195608
rect 670790 194032 670846 194041
rect 670790 193967 670846 193976
rect 670804 190641 670832 193967
rect 670790 190632 670846 190641
rect 670790 190567 670846 190576
rect 670698 189000 670754 189009
rect 670698 188935 670754 188944
rect 670712 185609 670740 188935
rect 670698 185600 670754 185609
rect 670698 185535 670754 185544
rect 670698 138136 670754 138145
rect 670698 138071 670754 138080
rect 670712 134745 670740 138071
rect 670698 134736 670754 134745
rect 670698 134671 670754 134680
rect 670056 132932 670108 132938
rect 670056 132874 670108 132880
rect 669504 132796 669556 132802
rect 669504 132738 669556 132744
rect 669320 132660 669372 132666
rect 669320 132602 669372 132608
rect 670792 131708 670844 131714
rect 670792 131650 670844 131656
rect 670804 129878 670832 131650
rect 670884 130076 670936 130082
rect 670884 130018 670936 130024
rect 669228 129872 669280 129878
rect 669228 129814 669280 129820
rect 670792 129872 670844 129878
rect 670792 129814 670844 129820
rect 666744 129804 666796 129810
rect 666744 129746 666796 129752
rect 666650 129568 666706 129577
rect 666650 129503 666706 129512
rect 666650 127936 666706 127945
rect 666650 127871 666706 127880
rect 666664 124545 666692 127871
rect 666650 124536 666706 124545
rect 666650 124471 666706 124480
rect 666650 122904 666706 122913
rect 666650 122839 666706 122848
rect 666664 119513 666692 122839
rect 666650 119504 666706 119513
rect 666650 119439 666706 119448
rect 670804 104145 670832 129814
rect 670896 129810 670924 130018
rect 670884 129804 670936 129810
rect 670884 129746 670936 129752
rect 670790 104136 670846 104145
rect 670790 104071 670846 104080
rect 670896 100881 670924 129746
rect 671172 107545 671200 218010
rect 671436 179376 671488 179382
rect 671436 179318 671488 179324
rect 671448 176934 671476 179318
rect 671436 176928 671488 176934
rect 671436 176870 671488 176876
rect 671816 173641 671844 705434
rect 671896 310480 671948 310486
rect 671896 310422 671948 310428
rect 671908 266150 671936 310422
rect 671896 266144 671948 266150
rect 671896 266086 671948 266092
rect 671896 176656 671948 176662
rect 671896 176598 671948 176604
rect 671908 175302 671936 176598
rect 671896 175296 671948 175302
rect 671896 175238 671948 175244
rect 671896 174480 671948 174486
rect 671896 174422 671948 174428
rect 671802 173632 671858 173641
rect 671802 173567 671858 173576
rect 671908 129742 671936 174422
rect 671896 129736 671948 129742
rect 671896 129678 671948 129684
rect 672000 129470 672028 984778
rect 672080 927444 672132 927450
rect 672080 927386 672132 927392
rect 672092 183841 672120 927386
rect 672172 749964 672224 749970
rect 672172 749906 672224 749912
rect 672078 183832 672134 183841
rect 672078 183767 672134 183776
rect 672184 178809 672212 749906
rect 672356 659728 672408 659734
rect 672356 659670 672408 659676
rect 672264 312112 672316 312118
rect 672264 312054 672316 312060
rect 672276 267510 672304 312054
rect 672264 267504 672316 267510
rect 672264 267446 672316 267452
rect 672170 178800 672226 178809
rect 672170 178735 672226 178744
rect 672172 176588 672224 176594
rect 672172 176530 672224 176536
rect 672184 174486 672212 176530
rect 672264 175296 672316 175302
rect 672264 175238 672316 175244
rect 672172 174480 672224 174486
rect 672172 174422 672224 174428
rect 672172 167884 672224 167890
rect 672172 167826 672224 167832
rect 672080 167476 672132 167482
rect 672080 167418 672132 167424
rect 671988 129464 672040 129470
rect 671988 129406 672040 129412
rect 671436 123140 671488 123146
rect 671436 123082 671488 123088
rect 671448 112713 671476 123082
rect 671434 112704 671490 112713
rect 671434 112639 671490 112648
rect 671158 107536 671214 107545
rect 671158 107471 671214 107480
rect 672000 102513 672028 129406
rect 672092 114345 672120 167418
rect 672184 116113 672212 167826
rect 672276 130694 672304 175238
rect 672368 168609 672396 659670
rect 672448 614780 672500 614786
rect 672448 614722 672500 614728
rect 672354 168600 672410 168609
rect 672354 168535 672410 168544
rect 672356 168292 672408 168298
rect 672356 168234 672408 168240
rect 672264 130688 672316 130694
rect 672264 130630 672316 130636
rect 672264 122324 672316 122330
rect 672264 122266 672316 122272
rect 672170 116104 672226 116113
rect 672170 116039 672226 116048
rect 672078 114336 672134 114345
rect 672078 114271 672134 114280
rect 672276 109313 672304 122266
rect 672368 117745 672396 168234
rect 672460 163577 672488 614722
rect 672552 579290 672580 985351
rect 672540 579284 672592 579290
rect 672540 579226 672592 579232
rect 672736 577658 672764 985487
rect 675680 970154 675708 985526
rect 674840 970148 674892 970154
rect 674840 970090 674892 970096
rect 675668 970148 675720 970154
rect 675668 970090 675720 970096
rect 674748 966204 674800 966210
rect 674748 966146 674800 966152
rect 673552 965796 673604 965802
rect 673552 965738 673604 965744
rect 673460 962056 673512 962062
rect 673460 961998 673512 962004
rect 673472 950774 673500 961998
rect 673460 950768 673512 950774
rect 673460 950710 673512 950716
rect 673564 933366 673592 965738
rect 673736 965048 673788 965054
rect 673736 964990 673788 964996
rect 673644 962532 673696 962538
rect 673644 962474 673696 962480
rect 673656 950858 673684 962474
rect 673748 950978 673776 964990
rect 673920 963212 673972 963218
rect 673920 963154 673972 963160
rect 673828 961376 673880 961382
rect 673828 961318 673880 961324
rect 673736 950972 673788 950978
rect 673736 950914 673788 950920
rect 673656 950830 673776 950858
rect 673644 950768 673696 950774
rect 673644 950710 673696 950716
rect 673552 933360 673604 933366
rect 673552 933302 673604 933308
rect 673656 932754 673684 950710
rect 673748 932822 673776 950830
rect 673736 932816 673788 932822
rect 673736 932758 673788 932764
rect 673644 932748 673696 932754
rect 673644 932690 673696 932696
rect 673840 932142 673868 961318
rect 673932 935338 673960 963154
rect 674656 958860 674708 958866
rect 674656 958802 674708 958808
rect 674288 958384 674340 958390
rect 674288 958326 674340 958332
rect 674012 954032 674064 954038
rect 674012 953974 674064 953980
rect 674024 951114 674052 953974
rect 674012 951108 674064 951114
rect 674012 951050 674064 951056
rect 674012 950972 674064 950978
rect 674012 950914 674064 950920
rect 674024 935474 674052 950914
rect 674012 935468 674064 935474
rect 674012 935410 674064 935416
rect 673920 935332 673972 935338
rect 673920 935274 673972 935280
rect 674300 932686 674328 958326
rect 674380 957772 674432 957778
rect 674380 957714 674432 957720
rect 674288 932680 674340 932686
rect 674288 932622 674340 932628
rect 673828 932136 673880 932142
rect 673828 932078 673880 932084
rect 674392 931734 674420 957714
rect 674564 957024 674616 957030
rect 674564 956966 674616 956972
rect 674472 955732 674524 955738
rect 674472 955674 674524 955680
rect 674484 932890 674512 955674
rect 674472 932884 674524 932890
rect 674472 932826 674524 932832
rect 674380 931728 674432 931734
rect 674380 931670 674432 931676
rect 674576 931326 674604 956966
rect 674668 935542 674696 958802
rect 674760 954038 674788 966146
rect 674748 954032 674800 954038
rect 674748 953974 674800 953980
rect 674748 953896 674800 953902
rect 674748 953838 674800 953844
rect 674760 935610 674788 953838
rect 674852 952202 674880 970090
rect 675404 966210 675432 966723
rect 675392 966204 675444 966210
rect 675392 966146 675444 966152
rect 675404 965802 675432 966076
rect 675392 965796 675444 965802
rect 675392 965738 675444 965744
rect 675496 965054 675524 965435
rect 675484 965048 675536 965054
rect 675484 964990 675536 964996
rect 675404 963218 675432 963595
rect 675392 963212 675444 963218
rect 675392 963154 675444 963160
rect 675496 962538 675524 963016
rect 675484 962532 675536 962538
rect 675484 962474 675536 962480
rect 675404 962062 675432 962404
rect 675392 962056 675444 962062
rect 675392 961998 675444 962004
rect 675404 961382 675432 961755
rect 675392 961376 675444 961382
rect 675392 961318 675444 961324
rect 675024 960560 675076 960566
rect 675024 960502 675076 960508
rect 675036 955534 675064 960502
rect 675404 958866 675432 959276
rect 675392 958860 675444 958866
rect 675392 958802 675444 958808
rect 675404 958390 675432 958732
rect 675392 958384 675444 958390
rect 675392 958326 675444 958332
rect 675496 957778 675524 958052
rect 675484 957772 675536 957778
rect 675484 957714 675536 957720
rect 675404 957030 675432 957440
rect 675392 957024 675444 957030
rect 675392 956966 675444 956972
rect 675496 955738 675524 956216
rect 675484 955732 675536 955738
rect 675484 955674 675536 955680
rect 675024 955528 675076 955534
rect 675024 955470 675076 955476
rect 675484 955528 675536 955534
rect 675484 955470 675536 955476
rect 675496 955060 675524 955470
rect 675404 953902 675432 954380
rect 675392 953896 675444 953902
rect 675392 953838 675444 953844
rect 674840 952196 674892 952202
rect 674840 952138 674892 952144
rect 675404 952066 675432 952544
rect 674840 952060 674892 952066
rect 674840 952002 674892 952008
rect 675392 952060 675444 952066
rect 675392 952002 675444 952008
rect 674748 935604 674800 935610
rect 674748 935546 674800 935552
rect 674656 935536 674708 935542
rect 674656 935478 674708 935484
rect 674852 934998 674880 952002
rect 675668 951788 675720 951794
rect 675668 951730 675720 951736
rect 675680 938777 675708 951730
rect 675760 951108 675812 951114
rect 675760 951050 675812 951056
rect 675666 938768 675722 938777
rect 675666 938703 675722 938712
rect 674840 934992 674892 934998
rect 674840 934934 674892 934940
rect 675772 934697 675800 951050
rect 703452 942948 703504 942954
rect 703452 942890 703504 942896
rect 709340 942948 709392 942954
rect 709340 942890 709392 942896
rect 703464 940522 703492 942890
rect 709352 940930 709380 942890
rect 703556 940914 703708 940930
rect 703544 940908 703708 940914
rect 703596 940902 703708 940908
rect 708880 940908 708932 940914
rect 703544 940850 703596 940856
rect 709228 940902 709380 940930
rect 708880 940850 708932 940856
rect 708052 940840 708104 940846
rect 704628 940778 704964 940794
rect 708104 940788 708308 940794
rect 708052 940782 708308 940788
rect 704628 940772 704976 940778
rect 704628 940766 704924 940772
rect 704924 940714 704976 940720
rect 707960 940772 708012 940778
rect 708064 940766 708308 940782
rect 707960 940714 708012 940720
rect 704832 940704 704884 940710
rect 704168 940630 704504 940658
rect 707040 940704 707092 940710
rect 704832 940646 704884 940652
rect 703464 940494 703708 940522
rect 704476 940302 704504 940630
rect 704844 940522 704872 940646
rect 705088 940630 705424 940658
rect 705548 940630 705884 940658
rect 706008 940630 706344 940658
rect 704628 940494 704872 940522
rect 705396 940438 705424 940630
rect 705752 940568 705804 940574
rect 705548 940516 705752 940522
rect 705548 940510 705804 940516
rect 705548 940494 705792 940510
rect 705856 940506 705884 940630
rect 706316 940574 706344 940630
rect 706212 940568 706264 940574
rect 706008 940516 706212 940522
rect 706008 940510 706264 940516
rect 706304 940568 706356 940574
rect 706304 940510 706356 940516
rect 705844 940500 705896 940506
rect 706008 940494 706252 940510
rect 706454 940508 706482 940644
rect 706684 940642 706928 940658
rect 707092 940652 707388 940658
rect 707040 940646 707388 940652
rect 706672 940636 706928 940642
rect 706724 940630 706928 940636
rect 707052 940630 707388 940646
rect 707604 940630 707848 940658
rect 706672 940578 706724 940584
rect 706580 940568 706632 940574
rect 706632 940516 706928 940522
rect 706580 940510 706928 940516
rect 706592 940494 706928 940510
rect 707052 940506 707388 940522
rect 707604 940506 707632 940630
rect 707972 940522 708000 940714
rect 708524 940630 708768 940658
rect 707040 940500 707388 940506
rect 705844 940442 705896 940448
rect 707092 940494 707388 940500
rect 707592 940500 707644 940506
rect 707040 940442 707092 940448
rect 707972 940494 708308 940522
rect 707592 940442 707644 940448
rect 705384 940432 705436 940438
rect 705088 940370 705332 940386
rect 705384 940374 705436 940380
rect 707500 940432 707552 940438
rect 707552 940380 707848 940386
rect 707500 940374 707848 940380
rect 705088 940364 705344 940370
rect 705088 940358 705292 940364
rect 707512 940358 707848 940374
rect 708524 940370 708552 940630
rect 708892 940522 708920 940850
rect 708892 940494 709228 940522
rect 708512 940364 708564 940370
rect 705292 940306 705344 940312
rect 708512 940306 708564 940312
rect 704464 940296 704516 940302
rect 704168 940234 704412 940250
rect 704464 940238 704516 940244
rect 708420 940296 708472 940302
rect 708472 940244 708768 940250
rect 708420 940238 708768 940244
rect 704168 940228 704424 940234
rect 704168 940222 704372 940228
rect 708432 940222 708768 940238
rect 704372 940170 704424 940176
rect 676310 939720 676366 939729
rect 676310 939655 676366 939664
rect 676126 939312 676182 939321
rect 676126 939247 676182 939256
rect 676140 938602 676168 939247
rect 676218 938904 676274 938913
rect 676218 938839 676220 938848
rect 676272 938839 676274 938848
rect 676220 938810 676272 938816
rect 676324 938738 676352 939655
rect 676312 938732 676364 938738
rect 676312 938674 676364 938680
rect 676128 938596 676180 938602
rect 676128 938538 676180 938544
rect 678978 937680 679034 937689
rect 678978 937615 679034 937624
rect 676218 936456 676274 936465
rect 676218 936391 676274 936400
rect 676034 935912 676090 935921
rect 676034 935847 676090 935856
rect 676048 935814 676076 935847
rect 676036 935808 676088 935814
rect 676036 935750 676088 935756
rect 676232 935746 676260 936391
rect 676220 935740 676272 935746
rect 676220 935682 676272 935688
rect 678992 935678 679020 937615
rect 678980 935672 679032 935678
rect 678980 935614 679032 935620
rect 676036 935604 676088 935610
rect 676036 935546 676088 935552
rect 675942 935504 675998 935513
rect 675942 935439 675944 935448
rect 675996 935439 675998 935448
rect 675944 935410 675996 935416
rect 675944 935332 675996 935338
rect 675944 935274 675996 935280
rect 675758 934688 675814 934697
rect 675758 934623 675814 934632
rect 675956 934289 675984 935274
rect 676048 935105 676076 935546
rect 676128 935536 676180 935542
rect 676128 935478 676180 935484
rect 676034 935096 676090 935105
rect 676034 935031 676090 935040
rect 676036 934992 676088 934998
rect 676036 934934 676088 934940
rect 675942 934280 675998 934289
rect 675942 934215 675998 934224
rect 676048 933473 676076 934934
rect 676140 934017 676168 935478
rect 676126 934008 676182 934017
rect 676126 933943 676182 933952
rect 676034 933464 676090 933473
rect 676034 933399 676090 933408
rect 676036 933360 676088 933366
rect 676036 933302 676088 933308
rect 676048 933065 676076 933302
rect 676034 933056 676090 933065
rect 676034 932991 676090 933000
rect 676036 932884 676088 932890
rect 676036 932826 676088 932832
rect 675944 932748 675996 932754
rect 675944 932690 675996 932696
rect 675956 932249 675984 932690
rect 675942 932240 675998 932249
rect 675942 932175 675998 932184
rect 675944 932136 675996 932142
rect 675944 932078 675996 932084
rect 674564 931320 674616 931326
rect 674564 931262 674616 931268
rect 675956 931025 675984 932078
rect 676048 931841 676076 932826
rect 676128 932816 676180 932822
rect 676126 932784 676128 932793
rect 676180 932784 676182 932793
rect 676126 932719 676182 932728
rect 676128 932680 676180 932686
rect 676128 932622 676180 932628
rect 676034 931832 676090 931841
rect 676034 931767 676090 931776
rect 676036 931728 676088 931734
rect 676036 931670 676088 931676
rect 676048 931433 676076 931670
rect 676034 931424 676090 931433
rect 676034 931359 676090 931368
rect 676036 931320 676088 931326
rect 676036 931262 676088 931268
rect 675942 931016 675998 931025
rect 675942 930951 675998 930960
rect 676048 930209 676076 931262
rect 676140 930753 676168 932622
rect 676126 930744 676182 930753
rect 676126 930679 676182 930688
rect 676034 930200 676090 930209
rect 676034 930135 676090 930144
rect 678978 929520 679034 929529
rect 678978 929455 679034 929464
rect 678992 929121 679020 929455
rect 678978 929112 679034 929121
rect 678978 929047 679034 929056
rect 684498 929112 684554 929121
rect 684498 929047 684554 929056
rect 678992 927450 679020 929047
rect 684512 928713 684540 929047
rect 684498 928704 684554 928713
rect 684498 928639 684554 928648
rect 678980 927444 679032 927450
rect 678980 927386 679032 927392
rect 675772 877305 675800 877540
rect 675758 877296 675814 877305
rect 675758 877231 675814 877240
rect 675680 876625 675708 876860
rect 675666 876616 675722 876625
rect 675666 876551 675722 876560
rect 675404 875945 675432 876248
rect 675390 875936 675446 875945
rect 675390 875871 675446 875880
rect 675496 874041 675524 874412
rect 675482 874032 675538 874041
rect 675482 873967 675538 873976
rect 675404 873526 675432 873868
rect 673552 873520 673604 873526
rect 673552 873462 673604 873468
rect 675392 873520 675444 873526
rect 675392 873462 675444 873468
rect 673460 782944 673512 782950
rect 673460 782886 673512 782892
rect 673472 770302 673500 782886
rect 673460 770296 673512 770302
rect 673460 770238 673512 770244
rect 673458 760336 673514 760345
rect 673458 760271 673514 760280
rect 673472 759257 673500 760271
rect 673458 759248 673514 759257
rect 673458 759183 673514 759192
rect 673368 759144 673420 759150
rect 673368 759086 673420 759092
rect 673380 723178 673408 759086
rect 673564 754934 673592 873462
rect 675404 872710 675432 873188
rect 674748 872704 674800 872710
rect 674748 872646 674800 872652
rect 675392 872704 675444 872710
rect 675392 872646 675444 872652
rect 673644 869848 673696 869854
rect 673644 869790 673696 869796
rect 673656 756158 673684 869790
rect 674196 869032 674248 869038
rect 674196 868974 674248 868980
rect 673736 868556 673788 868562
rect 673736 868498 673788 868504
rect 673644 756152 673696 756158
rect 673644 756094 673696 756100
rect 673552 754928 673604 754934
rect 673552 754870 673604 754876
rect 673748 753302 673776 868498
rect 673828 866516 673880 866522
rect 673828 866458 673880 866464
rect 673840 753506 673868 866458
rect 674012 864680 674064 864686
rect 674012 864622 674064 864628
rect 673920 862844 673972 862850
rect 673920 862786 673972 862792
rect 673932 756226 673960 862786
rect 674024 759014 674052 864622
rect 674208 792033 674236 868974
rect 674288 867808 674340 867814
rect 674288 867750 674340 867756
rect 674300 797745 674328 867750
rect 674760 854282 674788 872646
rect 675772 872273 675800 872576
rect 675758 872264 675814 872273
rect 675758 872199 675814 872208
rect 674932 870800 674984 870806
rect 674932 870742 674984 870748
rect 674944 866318 674972 870742
rect 675404 869854 675432 870060
rect 675392 869848 675444 869854
rect 675392 869790 675444 869796
rect 675404 869038 675432 869516
rect 675392 869032 675444 869038
rect 675392 868974 675444 868980
rect 675404 868562 675432 868875
rect 675392 868556 675444 868562
rect 675392 868498 675444 868504
rect 675404 867814 675432 868224
rect 675392 867808 675444 867814
rect 675392 867750 675444 867756
rect 675404 866522 675432 867035
rect 675392 866516 675444 866522
rect 675392 866458 675444 866464
rect 674932 866312 674984 866318
rect 674932 866254 674984 866260
rect 675392 866312 675444 866318
rect 675392 866254 675444 866260
rect 675404 865844 675432 866254
rect 675404 864686 675432 865195
rect 675392 864680 675444 864686
rect 675392 864622 675444 864628
rect 675496 862850 675524 863328
rect 675484 862844 675536 862850
rect 675484 862786 675536 862792
rect 674748 854276 674800 854282
rect 674748 854218 674800 854224
rect 675576 854276 675628 854282
rect 675576 854218 675628 854224
rect 674286 797736 674342 797745
rect 674286 797671 674342 797680
rect 675588 796278 675616 854218
rect 674564 796272 674616 796278
rect 674564 796214 674616 796220
rect 675576 796272 675628 796278
rect 675576 796214 675628 796220
rect 674194 792024 674250 792033
rect 674194 791959 674250 791968
rect 674380 784984 674432 784990
rect 674380 784926 674432 784932
rect 674288 780632 674340 780638
rect 674288 780574 674340 780580
rect 674196 779340 674248 779346
rect 674196 779282 674248 779288
rect 674208 770386 674236 779282
rect 674300 770574 674328 780574
rect 674392 777481 674420 784926
rect 674472 779816 674524 779822
rect 674472 779758 674524 779764
rect 674378 777472 674434 777481
rect 674378 777407 674434 777416
rect 674380 777368 674432 777374
rect 674380 777310 674432 777316
rect 674288 770568 674340 770574
rect 674288 770510 674340 770516
rect 674392 770522 674420 777310
rect 674484 773430 674512 779758
rect 674576 776914 674604 796214
rect 675404 787817 675432 788324
rect 675390 787808 675446 787817
rect 675390 787743 675446 787752
rect 675404 787409 675432 787679
rect 675390 787400 675446 787409
rect 675390 787335 675446 787344
rect 675404 786865 675432 787032
rect 675390 786856 675446 786865
rect 675390 786791 675446 786800
rect 675404 784990 675432 785196
rect 675392 784984 675444 784990
rect 675392 784926 675444 784932
rect 675404 784145 675432 784652
rect 675390 784136 675446 784145
rect 675390 784071 675446 784080
rect 675496 783873 675524 783972
rect 675482 783864 675538 783873
rect 675482 783799 675538 783808
rect 675496 782950 675524 783360
rect 675484 782944 675536 782950
rect 675484 782886 675536 782892
rect 674656 782468 674708 782474
rect 674656 782410 674708 782416
rect 674668 777102 674696 782410
rect 675496 780638 675524 780844
rect 675484 780632 675536 780638
rect 675484 780574 675536 780580
rect 675496 779822 675524 780300
rect 675484 779816 675536 779822
rect 675484 779758 675536 779764
rect 675404 779346 675432 779688
rect 675392 779340 675444 779346
rect 675392 779282 675444 779288
rect 675496 778666 675524 779008
rect 674748 778660 674800 778666
rect 674748 778602 674800 778608
rect 675484 778660 675536 778666
rect 675484 778602 675536 778608
rect 674656 777096 674708 777102
rect 674656 777038 674708 777044
rect 674576 776886 674696 776914
rect 674564 775532 674616 775538
rect 674564 775474 674616 775480
rect 674472 773424 674524 773430
rect 674472 773366 674524 773372
rect 674576 770658 674604 775474
rect 674668 773906 674696 776886
rect 674656 773900 674708 773906
rect 674656 773842 674708 773848
rect 674656 773628 674708 773634
rect 674656 773570 674708 773576
rect 674668 770794 674696 773570
rect 674760 773158 674788 778602
rect 675404 777374 675432 777852
rect 675392 777368 675444 777374
rect 675392 777310 675444 777316
rect 675392 777096 675444 777102
rect 675392 777038 675444 777044
rect 675404 776628 675432 777038
rect 675404 775538 675432 776016
rect 675392 775532 675444 775538
rect 675392 775474 675444 775480
rect 675208 773900 675260 773906
rect 675208 773842 675260 773848
rect 675220 773362 675248 773842
rect 675496 773634 675524 774180
rect 675484 773628 675536 773634
rect 675484 773570 675536 773576
rect 675668 773424 675720 773430
rect 675668 773366 675720 773372
rect 675208 773356 675260 773362
rect 675208 773298 675260 773304
rect 675576 773356 675628 773362
rect 675576 773298 675628 773304
rect 674748 773152 674800 773158
rect 674748 773094 674800 773100
rect 675484 773152 675536 773158
rect 675484 773094 675536 773100
rect 674668 770766 674788 770794
rect 674576 770630 674696 770658
rect 674564 770568 674616 770574
rect 674392 770494 674512 770522
rect 674564 770510 674616 770516
rect 674208 770358 674420 770386
rect 674288 770296 674340 770302
rect 674194 770264 674250 770273
rect 674288 770238 674340 770244
rect 674194 770199 674250 770208
rect 674012 759008 674064 759014
rect 674012 758950 674064 758956
rect 673920 756220 673972 756226
rect 673920 756162 673972 756168
rect 673828 753500 673880 753506
rect 673828 753442 673880 753448
rect 673736 753296 673788 753302
rect 673736 753238 673788 753244
rect 673920 738472 673972 738478
rect 673920 738414 673972 738420
rect 673736 734800 673788 734806
rect 673736 734742 673788 734748
rect 673644 734392 673696 734398
rect 673644 734334 673696 734340
rect 673552 733644 673604 733650
rect 673552 733586 673604 733592
rect 673368 723172 673420 723178
rect 673368 723114 673420 723120
rect 673092 714060 673144 714066
rect 673092 714002 673144 714008
rect 673000 688628 673052 688634
rect 673000 688570 673052 688576
rect 673012 616758 673040 688570
rect 673104 679046 673132 714002
rect 673564 710734 673592 733586
rect 673552 710728 673604 710734
rect 673552 710670 673604 710676
rect 673656 699825 673684 734334
rect 673748 730674 673776 734742
rect 673828 732352 673880 732358
rect 673828 732294 673880 732300
rect 673840 730810 673868 732294
rect 673932 731762 673960 738414
rect 674012 735480 674064 735486
rect 674012 735422 674064 735428
rect 674024 731950 674052 735422
rect 674012 731944 674064 731950
rect 674012 731886 674064 731892
rect 673932 731734 674052 731762
rect 673840 730782 673960 730810
rect 673748 730646 673868 730674
rect 673736 730516 673788 730522
rect 673736 730458 673788 730464
rect 673748 711090 673776 730458
rect 673840 714134 673868 730646
rect 673932 722906 673960 730782
rect 673920 722900 673972 722906
rect 673920 722842 673972 722848
rect 674024 721206 674052 731734
rect 674208 721342 674236 770199
rect 674196 721336 674248 721342
rect 674196 721278 674248 721284
rect 674012 721200 674064 721206
rect 674012 721142 674064 721148
rect 674196 721200 674248 721206
rect 674196 721142 674248 721148
rect 673828 714128 673880 714134
rect 673828 714070 673880 714076
rect 674208 711958 674236 721142
rect 674196 711952 674248 711958
rect 674196 711894 674248 711900
rect 673748 711062 673960 711090
rect 673736 710660 673788 710666
rect 673736 710602 673788 710608
rect 673642 699816 673698 699825
rect 673642 699751 673698 699760
rect 673644 690464 673696 690470
rect 673644 690406 673696 690412
rect 673184 689172 673236 689178
rect 673184 689114 673236 689120
rect 673092 679040 673144 679046
rect 673092 678982 673144 678988
rect 673092 668092 673144 668098
rect 673092 668034 673144 668040
rect 673104 637906 673132 668034
rect 673092 637900 673144 637906
rect 673092 637842 673144 637848
rect 673196 617982 673224 689114
rect 673276 687336 673328 687342
rect 673276 687278 673328 687284
rect 673288 618254 673316 687278
rect 673552 647760 673604 647766
rect 673552 647702 673604 647708
rect 673368 623960 673420 623966
rect 673368 623902 673420 623908
rect 673276 618248 673328 618254
rect 673276 618190 673328 618196
rect 673184 617976 673236 617982
rect 673184 617918 673236 617924
rect 673000 616752 673052 616758
rect 673000 616694 673052 616700
rect 673380 587926 673408 623902
rect 673368 587920 673420 587926
rect 673368 587862 673420 587868
rect 673276 579284 673328 579290
rect 673276 579226 673328 579232
rect 673092 578468 673144 578474
rect 673092 578410 673144 578416
rect 672724 577652 672776 577658
rect 672724 577594 672776 577600
rect 672540 568608 672592 568614
rect 672540 568550 672592 568556
rect 672446 163568 672502 163577
rect 672446 163503 672502 163512
rect 672552 158409 672580 568550
rect 673104 546310 673132 578410
rect 673184 577652 673236 577658
rect 673184 577594 673236 577600
rect 673092 546304 673144 546310
rect 673092 546246 673144 546252
rect 673196 533322 673224 577594
rect 673288 534954 673316 579226
rect 673368 576972 673420 576978
rect 673368 576914 673420 576920
rect 673276 534948 673328 534954
rect 673276 534890 673328 534896
rect 673184 533316 673236 533322
rect 673184 533258 673236 533264
rect 673380 532642 673408 576914
rect 673564 572422 673592 647702
rect 673656 620906 673684 690406
rect 673748 665106 673776 710602
rect 673828 683664 673880 683670
rect 673828 683606 673880 683612
rect 673736 665100 673788 665106
rect 673736 665042 673788 665048
rect 673736 645448 673788 645454
rect 673736 645390 673788 645396
rect 673748 637226 673776 645390
rect 673736 637220 673788 637226
rect 673736 637162 673788 637168
rect 673840 620974 673868 683606
rect 673932 667894 673960 711062
rect 674012 710728 674064 710734
rect 674012 710670 674064 710676
rect 674024 699689 674052 710670
rect 674300 707878 674328 770238
rect 674392 708286 674420 770358
rect 674484 709306 674512 770494
rect 674576 712026 674604 770510
rect 674668 738478 674696 770630
rect 674656 738472 674708 738478
rect 674656 738414 674708 738420
rect 674656 738336 674708 738342
rect 674656 738278 674708 738284
rect 674668 732086 674696 738278
rect 674656 732080 674708 732086
rect 674656 732022 674708 732028
rect 674656 731944 674708 731950
rect 674656 731886 674708 731892
rect 674564 712020 674616 712026
rect 674564 711962 674616 711968
rect 674668 710734 674696 731886
rect 674656 710728 674708 710734
rect 674656 710670 674708 710676
rect 674760 710598 674788 770766
rect 675496 744161 675524 773094
rect 675588 753817 675616 773298
rect 675574 753808 675630 753817
rect 675574 753743 675630 753752
rect 675482 744152 675538 744161
rect 675482 744087 675538 744096
rect 675680 744025 675708 773366
rect 679070 772712 679126 772721
rect 679070 772647 679126 772656
rect 678978 761288 679034 761297
rect 678978 761223 679034 761232
rect 676218 760880 676274 760889
rect 676218 760815 676274 760824
rect 676126 760472 676182 760481
rect 676126 760407 676182 760416
rect 676140 759354 676168 760407
rect 676232 759626 676260 760815
rect 676310 759656 676366 759665
rect 676220 759620 676272 759626
rect 676310 759591 676366 759600
rect 676220 759562 676272 759568
rect 676128 759348 676180 759354
rect 676128 759290 676180 759296
rect 676036 759144 676088 759150
rect 676034 759112 676036 759121
rect 676088 759112 676090 759121
rect 676324 759082 676352 759591
rect 678992 759490 679020 761223
rect 679084 759665 679112 772647
rect 708512 762544 708564 762550
rect 704168 762482 704504 762498
rect 708564 762492 708768 762498
rect 708512 762486 708768 762492
rect 704168 762476 704516 762482
rect 704168 762470 704464 762476
rect 704464 762418 704516 762424
rect 708420 762476 708472 762482
rect 708524 762470 708768 762486
rect 708420 762418 708472 762424
rect 704372 762408 704424 762414
rect 703556 762334 703708 762362
rect 707500 762408 707552 762414
rect 704372 762350 704424 762356
rect 703556 761870 703584 762334
rect 704384 762090 704412 762350
rect 704628 762334 704964 762362
rect 705088 762334 705424 762362
rect 705548 762334 705884 762362
rect 706008 762334 706344 762362
rect 704168 762062 704412 762090
rect 704936 762006 704964 762334
rect 705292 762272 705344 762278
rect 705292 762214 705344 762220
rect 705304 762090 705332 762214
rect 705088 762062 705332 762090
rect 705396 762074 705424 762334
rect 705752 762272 705804 762278
rect 705752 762214 705804 762220
rect 705764 762090 705792 762214
rect 705856 762210 705884 762334
rect 706212 762272 706264 762278
rect 706212 762214 706264 762220
rect 705844 762204 705896 762210
rect 705844 762146 705896 762152
rect 706224 762090 706252 762214
rect 706316 762142 706344 762334
rect 706592 762334 706928 762362
rect 707052 762346 707388 762362
rect 707552 762356 707848 762362
rect 707500 762350 707848 762356
rect 707040 762340 707388 762346
rect 706592 762278 706620 762334
rect 707092 762334 707388 762340
rect 707512 762334 707848 762350
rect 708064 762334 708308 762362
rect 707040 762282 707092 762288
rect 706580 762272 706632 762278
rect 706580 762214 706632 762220
rect 705384 762068 705436 762074
rect 705548 762062 705792 762090
rect 706008 762062 706252 762090
rect 706304 762136 706356 762142
rect 706304 762078 706356 762084
rect 706454 762076 706482 762212
rect 707040 762204 707092 762210
rect 707040 762146 707092 762152
rect 706580 762136 706632 762142
rect 707052 762090 707080 762146
rect 706632 762084 706928 762090
rect 706580 762078 706928 762084
rect 706592 762062 706928 762078
rect 707052 762062 707388 762090
rect 707512 762074 707848 762090
rect 708064 762074 708092 762334
rect 708432 762090 708460 762418
rect 708984 762334 709228 762362
rect 707500 762068 707848 762074
rect 705384 762010 705436 762016
rect 707552 762062 707848 762068
rect 708052 762068 708104 762074
rect 707500 762010 707552 762016
rect 708432 762062 708768 762090
rect 708052 762010 708104 762016
rect 704924 762000 704976 762006
rect 704628 761938 704872 761954
rect 704924 761942 704976 761948
rect 707960 762000 708012 762006
rect 708012 761948 708308 761954
rect 707960 761942 708308 761948
rect 704628 761932 704884 761938
rect 704628 761926 704832 761932
rect 707972 761926 708308 761942
rect 708984 761938 709012 762334
rect 708972 761932 709024 761938
rect 704832 761874 704884 761880
rect 708972 761874 709024 761880
rect 703544 761864 703596 761870
rect 708880 761864 708932 761870
rect 703544 761806 703596 761812
rect 703708 761802 704044 761818
rect 708932 761812 709228 761818
rect 708880 761806 709228 761812
rect 703708 761796 704056 761802
rect 703708 761790 704004 761796
rect 708892 761790 709228 761806
rect 704004 761738 704056 761744
rect 679070 759656 679126 759665
rect 679070 759591 679126 759600
rect 678980 759484 679032 759490
rect 678980 759426 679032 759432
rect 676034 759047 676090 759056
rect 676312 759076 676364 759082
rect 676312 759018 676364 759024
rect 676036 759008 676088 759014
rect 676036 758950 676088 758956
rect 676048 756673 676076 758950
rect 678978 758432 679034 758441
rect 678978 758367 679034 758376
rect 676126 758024 676182 758033
rect 676126 757959 676182 757968
rect 676034 756664 676090 756673
rect 676034 756599 676090 756608
rect 676140 756498 676168 757959
rect 676310 757616 676366 757625
rect 676310 757551 676366 757560
rect 676218 757208 676274 757217
rect 676218 757143 676274 757152
rect 676128 756492 676180 756498
rect 676128 756434 676180 756440
rect 676232 756430 676260 757143
rect 676220 756424 676272 756430
rect 676220 756366 676272 756372
rect 676324 756362 676352 757551
rect 676312 756356 676364 756362
rect 676312 756298 676364 756304
rect 678992 756294 679020 758367
rect 678980 756288 679032 756294
rect 678980 756230 679032 756236
rect 676036 756220 676088 756226
rect 676036 756162 676088 756168
rect 676048 755041 676076 756162
rect 676128 756152 676180 756158
rect 676128 756094 676180 756100
rect 676140 755585 676168 756094
rect 676126 755576 676182 755585
rect 676126 755511 676182 755520
rect 676034 755032 676090 755041
rect 676034 754967 676090 754976
rect 676036 754928 676088 754934
rect 676036 754870 676088 754876
rect 676048 754225 676076 754870
rect 676034 754216 676090 754225
rect 676034 754151 676090 754160
rect 676036 753500 676088 753506
rect 676036 753442 676088 753448
rect 676048 753409 676076 753442
rect 676034 753400 676090 753409
rect 676034 753335 676090 753344
rect 676036 753296 676088 753302
rect 676036 753238 676088 753244
rect 676048 753001 676076 753238
rect 676034 752992 676090 753001
rect 676034 752927 676090 752936
rect 679254 751088 679310 751097
rect 679254 751023 679310 751032
rect 679268 750689 679296 751023
rect 678978 750680 679034 750689
rect 678978 750615 679034 750624
rect 679254 750680 679310 750689
rect 679254 750615 679310 750624
rect 678992 750281 679020 750615
rect 678978 750272 679034 750281
rect 678978 750207 679034 750216
rect 679268 749970 679296 750615
rect 679256 749964 679308 749970
rect 679256 749906 679308 749912
rect 675666 744016 675722 744025
rect 675666 743951 675722 743960
rect 675772 742937 675800 743308
rect 675758 742928 675814 742937
rect 675758 742863 675814 742872
rect 675772 742529 675800 742696
rect 675758 742520 675814 742529
rect 675758 742455 675814 742464
rect 675496 741713 675524 742016
rect 675482 741704 675538 741713
rect 675482 741639 675538 741648
rect 675404 739809 675432 740180
rect 675390 739800 675446 739809
rect 675390 739735 675446 739744
rect 675404 739129 675432 739636
rect 675390 739120 675446 739129
rect 675390 739055 675446 739064
rect 675680 738585 675708 739024
rect 675666 738576 675722 738585
rect 675666 738511 675722 738520
rect 675772 738041 675800 738344
rect 675758 738032 675814 738041
rect 675758 737967 675814 737976
rect 675404 735486 675432 735896
rect 675392 735480 675444 735486
rect 675392 735422 675444 735428
rect 675404 734806 675432 735319
rect 675392 734800 675444 734806
rect 675392 734742 675444 734748
rect 675404 734398 675432 734672
rect 675392 734392 675444 734398
rect 675392 734334 675444 734340
rect 675404 733650 675432 734031
rect 675392 733644 675444 733650
rect 675392 733586 675444 733592
rect 675404 732358 675432 732836
rect 675392 732352 675444 732358
rect 675392 732294 675444 732300
rect 675392 732080 675444 732086
rect 675392 732022 675444 732028
rect 675404 731612 675432 732022
rect 675404 730522 675432 731000
rect 675392 730516 675444 730522
rect 675392 730458 675444 730464
rect 675496 728958 675524 729164
rect 674840 728952 674892 728958
rect 674840 728894 674892 728900
rect 675484 728952 675536 728958
rect 675484 728894 675536 728900
rect 674852 710666 674880 728894
rect 678980 723172 679032 723178
rect 678980 723114 679032 723120
rect 675484 722900 675536 722906
rect 675484 722842 675536 722848
rect 674932 721336 674984 721342
rect 674932 721278 674984 721284
rect 674944 712094 674972 721278
rect 674932 712088 674984 712094
rect 674932 712030 674984 712036
rect 674840 710660 674892 710666
rect 674840 710602 674892 710608
rect 674748 710592 674800 710598
rect 674748 710534 674800 710540
rect 674472 709300 674524 709306
rect 674472 709242 674524 709248
rect 674380 708280 674432 708286
rect 674380 708222 674432 708228
rect 674288 707872 674340 707878
rect 674288 707814 674340 707820
rect 675496 699718 675524 722842
rect 676036 716576 676088 716582
rect 676034 716544 676036 716553
rect 676088 716544 676090 716553
rect 676034 716479 676090 716488
rect 676036 716168 676088 716174
rect 676034 716136 676036 716145
rect 676088 716136 676090 716145
rect 676034 716071 676090 716080
rect 676036 715760 676088 715766
rect 676034 715728 676036 715737
rect 676088 715728 676090 715737
rect 676034 715663 676090 715672
rect 676034 715320 676090 715329
rect 676034 715255 676036 715264
rect 676088 715255 676090 715264
rect 676036 715226 676088 715232
rect 676036 714944 676088 714950
rect 676034 714912 676036 714921
rect 676088 714912 676090 714921
rect 676034 714847 676090 714856
rect 678992 714513 679020 723114
rect 703452 720452 703504 720458
rect 703452 720394 703504 720400
rect 709248 720452 709300 720458
rect 709248 720394 709300 720400
rect 703464 717482 703492 720394
rect 709260 719522 709288 720394
rect 709260 719494 709380 719522
rect 704464 717528 704516 717534
rect 703464 717454 703708 717482
rect 704177 717476 704464 717482
rect 704177 717470 704516 717476
rect 708420 717528 708472 717534
rect 708420 717470 708472 717476
rect 704177 717454 704504 717470
rect 704464 717392 704516 717398
rect 705384 717392 705436 717398
rect 704464 717334 704516 717340
rect 704476 717074 704504 717334
rect 704637 717318 704964 717346
rect 705097 717340 705384 717346
rect 707500 717392 707552 717398
rect 705097 717334 705436 717340
rect 705097 717318 705424 717334
rect 705557 717318 705884 717346
rect 706017 717318 706344 717346
rect 704168 717046 704504 717074
rect 704936 716990 704964 717318
rect 705752 717256 705804 717262
rect 705752 717198 705804 717204
rect 705764 717074 705792 717198
rect 705856 717194 705884 717318
rect 706212 717256 706264 717262
rect 706212 717198 706264 717204
rect 705844 717188 705896 717194
rect 705844 717130 705896 717136
rect 706224 717074 706252 717198
rect 706316 717126 706344 717318
rect 706454 717196 706482 717332
rect 706592 717318 706928 717346
rect 707052 717330 707388 717346
rect 707500 717334 707552 717340
rect 707040 717324 707388 717330
rect 706592 717262 706620 717318
rect 707092 717318 707388 717324
rect 707040 717266 707092 717272
rect 706580 717256 706632 717262
rect 706580 717198 706632 717204
rect 707040 717188 707092 717194
rect 707040 717130 707092 717136
rect 705088 717058 705424 717074
rect 705088 717052 705436 717058
rect 705088 717046 705384 717052
rect 705548 717046 705792 717074
rect 706008 717046 706252 717074
rect 706304 717120 706356 717126
rect 706304 717062 706356 717068
rect 706580 717120 706632 717126
rect 707052 717074 707080 717130
rect 707512 717074 707540 717334
rect 707604 717318 707848 717346
rect 708064 717318 708308 717346
rect 707604 717194 707632 717318
rect 707592 717188 707644 717194
rect 707592 717130 707644 717136
rect 706632 717068 706928 717074
rect 706580 717062 706928 717068
rect 706592 717046 706928 717062
rect 707052 717046 707388 717074
rect 707512 717046 707848 717074
rect 708064 717058 708092 717318
rect 708432 717074 708460 717470
rect 708524 717466 708768 717482
rect 708512 717460 708768 717466
rect 708564 717454 708768 717460
rect 708512 717402 708564 717408
rect 708892 717318 709228 717346
rect 708052 717052 708104 717058
rect 705384 716994 705436 717000
rect 708432 717046 708768 717074
rect 708052 716994 708104 717000
rect 704924 716984 704976 716990
rect 704628 716922 704872 716938
rect 704924 716926 704976 716932
rect 707960 716984 708012 716990
rect 708012 716932 708308 716938
rect 707960 716926 708308 716932
rect 704628 716916 704884 716922
rect 704628 716910 704832 716916
rect 707972 716910 708308 716926
rect 704832 716858 704884 716864
rect 708892 716854 708920 717318
rect 709352 717074 709380 719494
rect 709228 717046 709380 717074
rect 703544 716848 703596 716854
rect 708880 716848 708932 716854
rect 703596 716796 703708 716802
rect 703544 716790 703708 716796
rect 708880 716790 708932 716796
rect 703556 716774 703708 716790
rect 678978 714504 679034 714513
rect 678978 714439 679034 714448
rect 675668 714128 675720 714134
rect 675668 714070 675720 714076
rect 676034 714096 676090 714105
rect 675576 710728 675628 710734
rect 675576 710670 675628 710676
rect 674748 699712 674800 699718
rect 674010 699680 674066 699689
rect 674748 699654 674800 699660
rect 675484 699712 675536 699718
rect 675484 699654 675536 699660
rect 674010 699615 674066 699624
rect 674656 699644 674708 699650
rect 674656 699586 674708 699592
rect 674564 691416 674616 691422
rect 674564 691358 674616 691364
rect 674576 687070 674604 691358
rect 674564 687064 674616 687070
rect 674564 687006 674616 687012
rect 674288 685500 674340 685506
rect 674288 685442 674340 685448
rect 673920 667888 673972 667894
rect 673920 667830 673972 667836
rect 673920 644156 673972 644162
rect 673920 644098 673972 644104
rect 673828 620968 673880 620974
rect 673828 620910 673880 620916
rect 673644 620900 673696 620906
rect 673644 620842 673696 620848
rect 673736 599140 673788 599146
rect 673736 599082 673788 599088
rect 673644 598460 673696 598466
rect 673644 598402 673696 598408
rect 673656 583778 673684 598402
rect 673644 583772 673696 583778
rect 673644 583714 673696 583720
rect 673552 572416 673604 572422
rect 673552 572358 673604 572364
rect 673552 559564 673604 559570
rect 673552 559506 673604 559512
rect 673460 554600 673512 554606
rect 673460 554542 673512 554548
rect 672816 532636 672868 532642
rect 672816 532578 672868 532584
rect 673368 532636 673420 532642
rect 673368 532578 673420 532584
rect 672632 524476 672684 524482
rect 672632 524418 672684 524424
rect 672538 158400 672594 158409
rect 672538 158335 672594 158344
rect 672644 153377 672672 524418
rect 672724 481092 672776 481098
rect 672724 481034 672776 481040
rect 672630 153368 672686 153377
rect 672630 153303 672686 153312
rect 672736 148209 672764 481034
rect 672828 278497 672856 532578
rect 673472 482934 673500 554542
rect 673564 487490 673592 559506
rect 673644 553240 673696 553246
rect 673644 553182 673696 553188
rect 673552 487484 673604 487490
rect 673552 487426 673604 487432
rect 673656 483002 673684 553182
rect 673748 527882 673776 599082
rect 673828 597168 673880 597174
rect 673828 597110 673880 597116
rect 673840 583914 673868 597110
rect 673828 583908 673880 583914
rect 673828 583850 673880 583856
rect 673828 583772 673880 583778
rect 673828 583714 673880 583720
rect 673736 527876 673788 527882
rect 673736 527818 673788 527824
rect 673840 527134 673868 583714
rect 673932 572830 673960 644098
rect 674196 643408 674248 643414
rect 674196 643350 674248 643356
rect 674012 642116 674064 642122
rect 674012 642058 674064 642064
rect 674024 637362 674052 642058
rect 674208 638058 674236 643350
rect 674300 638178 674328 685442
rect 674564 669044 674616 669050
rect 674564 668986 674616 668992
rect 674380 649596 674432 649602
rect 674380 649538 674432 649544
rect 674392 638178 674420 649538
rect 674472 647352 674524 647358
rect 674472 647294 674524 647300
rect 674484 641714 674512 647294
rect 674472 641708 674524 641714
rect 674472 641650 674524 641656
rect 674472 640280 674524 640286
rect 674472 640222 674524 640228
rect 674288 638172 674340 638178
rect 674288 638114 674340 638120
rect 674380 638172 674432 638178
rect 674380 638114 674432 638120
rect 674208 638030 674420 638058
rect 674196 637968 674248 637974
rect 674196 637910 674248 637916
rect 674208 637786 674236 637910
rect 674208 637758 674328 637786
rect 674012 637356 674064 637362
rect 674012 637298 674064 637304
rect 674196 637356 674248 637362
rect 674196 637298 674248 637304
rect 674012 637220 674064 637226
rect 674012 637162 674064 637168
rect 674024 576094 674052 637162
rect 674012 576088 674064 576094
rect 674012 576030 674064 576036
rect 674208 573646 674236 637298
rect 674300 623762 674328 637758
rect 674288 623756 674340 623762
rect 674288 623698 674340 623704
rect 674392 608977 674420 638030
rect 674378 608968 674434 608977
rect 674378 608903 674434 608912
rect 674380 608796 674432 608802
rect 674380 608738 674432 608744
rect 674288 600432 674340 600438
rect 674288 600374 674340 600380
rect 674196 573640 674248 573646
rect 674196 573582 674248 573588
rect 673920 572824 673972 572830
rect 673920 572766 673972 572772
rect 674196 555280 674248 555286
rect 674196 555222 674248 555228
rect 673920 553784 673972 553790
rect 673920 553726 673972 553732
rect 673828 527128 673880 527134
rect 673828 527070 673880 527076
rect 673932 483886 673960 553726
rect 674012 551948 674064 551954
rect 674012 551890 674064 551896
rect 674024 485518 674052 551890
rect 674208 487150 674236 555222
rect 674300 531146 674328 600374
rect 674392 596714 674420 608738
rect 674484 596834 674512 640222
rect 674576 624306 674604 668986
rect 674668 667826 674696 699586
rect 674760 671294 674788 699654
rect 675588 699650 675616 710670
rect 675576 699644 675628 699650
rect 675576 699586 675628 699592
rect 675680 699553 675708 714070
rect 676034 714031 676036 714040
rect 676088 714031 676090 714040
rect 676036 714002 676088 714008
rect 676034 713688 676090 713697
rect 676034 713623 676036 713632
rect 676088 713623 676090 713632
rect 676036 713594 676088 713600
rect 676034 713280 676090 713289
rect 676034 713215 676036 713224
rect 676088 713215 676090 713224
rect 676036 713186 676088 713192
rect 676036 712904 676088 712910
rect 676034 712872 676036 712881
rect 676088 712872 676090 712881
rect 676034 712807 676090 712816
rect 676036 712496 676088 712502
rect 676034 712464 676036 712473
rect 676088 712464 676090 712473
rect 676034 712399 676090 712408
rect 676036 712088 676088 712094
rect 676036 712030 676088 712036
rect 675944 712020 675996 712026
rect 675944 711962 675996 711968
rect 675852 711952 675904 711958
rect 675852 711894 675904 711900
rect 675864 711657 675892 711894
rect 675850 711648 675906 711657
rect 675850 711583 675906 711592
rect 675850 710560 675906 710569
rect 675850 710495 675906 710504
rect 675864 707169 675892 710495
rect 675956 710433 675984 711962
rect 676048 710841 676076 712030
rect 676034 710832 676090 710841
rect 676034 710767 676090 710776
rect 676036 710592 676088 710598
rect 676036 710534 676088 710540
rect 676586 710594 676642 710603
rect 675942 710424 675998 710433
rect 675942 710359 675998 710368
rect 676048 710025 676076 710534
rect 676586 710529 676642 710538
rect 676034 710016 676090 710025
rect 676034 709951 676090 709960
rect 676036 709300 676088 709306
rect 676036 709242 676088 709248
rect 676048 708393 676076 709242
rect 676034 708384 676090 708393
rect 676034 708319 676090 708328
rect 676036 708280 676088 708286
rect 676036 708222 676088 708228
rect 676048 707985 676076 708222
rect 676034 707976 676090 707985
rect 676034 707911 676090 707920
rect 676036 707872 676088 707878
rect 676036 707814 676088 707820
rect 676048 707577 676076 707814
rect 676034 707568 676090 707577
rect 676034 707503 676090 707512
rect 676600 707470 676628 710529
rect 676036 707464 676088 707470
rect 676036 707406 676088 707412
rect 676588 707464 676640 707470
rect 676588 707406 676640 707412
rect 675850 707160 675906 707169
rect 675850 707095 675906 707104
rect 676048 706761 676076 707406
rect 676034 706752 676090 706761
rect 676034 706687 676090 706696
rect 675942 706344 675998 706353
rect 675942 706279 675998 706288
rect 675956 705537 675984 706279
rect 676034 705936 676090 705945
rect 676034 705871 676090 705880
rect 675942 705528 675998 705537
rect 675942 705463 675944 705472
rect 675996 705463 675998 705472
rect 675944 705434 675996 705440
rect 675956 705403 675984 705434
rect 676048 705129 676076 705871
rect 676034 705120 676090 705129
rect 676034 705055 676090 705064
rect 675666 699544 675722 699553
rect 675666 699479 675722 699488
rect 675496 698193 675524 698323
rect 675482 698184 675538 698193
rect 675482 698119 675538 698128
rect 675404 697377 675432 697680
rect 675390 697368 675446 697377
rect 675390 697303 675446 697312
rect 675404 696697 675432 697035
rect 675390 696688 675446 696697
rect 675390 696623 675446 696632
rect 675404 694793 675432 695195
rect 675390 694784 675446 694793
rect 675390 694719 675446 694728
rect 675496 694385 675524 694620
rect 675482 694376 675538 694385
rect 675482 694311 675538 694320
rect 675404 693569 675432 694008
rect 675390 693560 675446 693569
rect 675390 693495 675446 693504
rect 675772 693025 675800 693328
rect 675758 693016 675814 693025
rect 675758 692951 675814 692960
rect 675404 690470 675432 690880
rect 675392 690464 675444 690470
rect 675392 690406 675444 690412
rect 675772 690169 675800 690336
rect 675758 690160 675814 690169
rect 675758 690095 675814 690104
rect 675496 689178 675524 689656
rect 675484 689172 675536 689178
rect 675484 689114 675536 689120
rect 675404 688634 675432 689044
rect 675392 688628 675444 688634
rect 675392 688570 675444 688576
rect 675404 687342 675432 687820
rect 675392 687336 675444 687342
rect 675392 687278 675444 687284
rect 675484 687064 675536 687070
rect 675484 687006 675536 687012
rect 675496 686664 675524 687006
rect 675404 685506 675432 685984
rect 675392 685500 675444 685506
rect 675392 685442 675444 685448
rect 675496 683670 675524 684148
rect 675484 683664 675536 683670
rect 675484 683606 675536 683612
rect 678980 679040 679032 679046
rect 678980 678982 679032 678988
rect 674748 671288 674800 671294
rect 674748 671230 674800 671236
rect 675208 671288 675260 671294
rect 675208 671230 675260 671236
rect 674748 667956 674800 667962
rect 674748 667898 674800 667904
rect 674656 667820 674708 667826
rect 674656 667762 674708 667768
rect 674760 647358 674788 667898
rect 675220 665174 675248 671230
rect 676218 671120 676274 671129
rect 676218 671055 676274 671064
rect 676036 671016 676088 671022
rect 676034 670984 676036 670993
rect 676088 670984 676090 670993
rect 676034 670919 676090 670928
rect 676232 670818 676260 671055
rect 676220 670812 676272 670818
rect 676220 670754 676272 670760
rect 676036 670608 676088 670614
rect 676034 670576 676036 670585
rect 676088 670576 676090 670585
rect 676034 670511 676090 670520
rect 676220 670336 676272 670342
rect 676218 670304 676220 670313
rect 676272 670304 676274 670313
rect 676218 670239 676274 670248
rect 676034 669760 676090 669769
rect 676034 669695 676090 669704
rect 676048 669050 676076 669695
rect 678992 669497 679020 678982
rect 703452 672376 703504 672382
rect 703452 672318 703504 672324
rect 703464 671922 703492 672318
rect 703556 672314 703708 672330
rect 708984 672314 709228 672330
rect 703544 672308 703708 672314
rect 703596 672302 703708 672308
rect 708880 672308 708932 672314
rect 703544 672250 703596 672256
rect 708880 672250 708932 672256
rect 708972 672308 709228 672314
rect 709024 672302 709228 672308
rect 708972 672250 709024 672256
rect 708052 672240 708104 672246
rect 704628 672178 704964 672194
rect 708104 672188 708308 672194
rect 708052 672182 708308 672188
rect 704628 672172 704976 672178
rect 704628 672166 704924 672172
rect 704924 672114 704976 672120
rect 707960 672172 708012 672178
rect 708064 672166 708308 672182
rect 707960 672114 708012 672120
rect 704832 672104 704884 672110
rect 704168 672030 704504 672058
rect 707040 672104 707092 672110
rect 704832 672046 704884 672052
rect 703464 671894 703708 671922
rect 704476 671702 704504 672030
rect 704844 671922 704872 672046
rect 705088 672030 705424 672058
rect 705548 672030 705884 672058
rect 706008 672030 706344 672058
rect 704628 671894 704872 671922
rect 705396 671838 705424 672030
rect 705752 671968 705804 671974
rect 705548 671916 705752 671922
rect 705548 671910 705804 671916
rect 705548 671894 705792 671910
rect 705856 671906 705884 672030
rect 706316 671974 706344 672030
rect 706212 671968 706264 671974
rect 706008 671916 706212 671922
rect 706008 671910 706264 671916
rect 706304 671968 706356 671974
rect 706304 671910 706356 671916
rect 705844 671900 705896 671906
rect 706008 671894 706252 671910
rect 706454 671908 706482 672044
rect 706684 672042 706928 672058
rect 707092 672052 707388 672058
rect 707040 672046 707388 672052
rect 706672 672036 706928 672042
rect 706724 672030 706928 672036
rect 707052 672030 707388 672046
rect 707604 672030 707848 672058
rect 706672 671978 706724 671984
rect 706580 671968 706632 671974
rect 706632 671916 706928 671922
rect 706580 671910 706928 671916
rect 706592 671894 706928 671910
rect 707052 671906 707388 671922
rect 707604 671906 707632 672030
rect 707972 671922 708000 672114
rect 708524 672030 708768 672058
rect 707040 671900 707388 671906
rect 705844 671842 705896 671848
rect 707092 671894 707388 671900
rect 707592 671900 707644 671906
rect 707040 671842 707092 671848
rect 707972 671894 708308 671922
rect 707592 671842 707644 671848
rect 705384 671832 705436 671838
rect 705088 671770 705332 671786
rect 705384 671774 705436 671780
rect 707500 671832 707552 671838
rect 707552 671780 707848 671786
rect 707500 671774 707848 671780
rect 705088 671764 705344 671770
rect 705088 671758 705292 671764
rect 707512 671758 707848 671774
rect 708524 671770 708552 672030
rect 708892 671922 708920 672250
rect 708892 671894 709228 671922
rect 708512 671764 708564 671770
rect 705292 671706 705344 671712
rect 708512 671706 708564 671712
rect 704464 671696 704516 671702
rect 704168 671634 704412 671650
rect 704464 671638 704516 671644
rect 708420 671696 708472 671702
rect 708472 671644 708768 671650
rect 708420 671638 708768 671644
rect 704168 671628 704424 671634
rect 704168 671622 704372 671628
rect 708432 671622 708768 671638
rect 704372 671570 704424 671576
rect 678978 669488 679034 669497
rect 678978 669423 679034 669432
rect 676036 669044 676088 669050
rect 676036 668986 676088 668992
rect 676034 668944 676090 668953
rect 676034 668879 676090 668888
rect 675942 668128 675998 668137
rect 675942 668063 675944 668072
rect 675996 668063 675998 668072
rect 675944 668034 675996 668040
rect 676048 667962 676076 668879
rect 676220 668704 676272 668710
rect 676218 668672 676220 668681
rect 676272 668672 676274 668681
rect 676218 668607 676274 668616
rect 676036 667956 676088 667962
rect 676036 667898 676088 667904
rect 676128 667888 676180 667894
rect 676128 667830 676180 667836
rect 676036 667820 676088 667826
rect 676036 667762 676088 667768
rect 675944 667752 675996 667758
rect 675942 667720 675944 667729
rect 675996 667720 675998 667729
rect 675942 667655 675998 667664
rect 676048 665281 676076 667762
rect 676140 666641 676168 667830
rect 676126 666632 676182 666641
rect 676126 666567 676182 666576
rect 676034 665272 676090 665281
rect 676034 665207 676090 665216
rect 675208 665168 675260 665174
rect 675208 665110 675260 665116
rect 676036 665168 676088 665174
rect 676036 665110 676088 665116
rect 676048 663241 676076 665110
rect 676128 665100 676180 665106
rect 676128 665042 676180 665048
rect 676140 665009 676168 665042
rect 676126 665000 676182 665009
rect 676126 664935 676182 664944
rect 676034 663232 676090 663241
rect 676034 663167 676090 663176
rect 678978 660920 679034 660929
rect 678978 660855 679034 660864
rect 678992 660521 679020 660855
rect 678978 660512 679034 660521
rect 678978 660447 679034 660456
rect 684498 660512 684554 660521
rect 684498 660447 684554 660456
rect 678992 659734 679020 660447
rect 684512 660113 684540 660447
rect 684498 660104 684554 660113
rect 684498 660039 684554 660048
rect 678980 659728 679032 659734
rect 678980 659670 679032 659676
rect 675404 652905 675432 653140
rect 675390 652896 675446 652905
rect 675390 652831 675446 652840
rect 675496 652225 675524 652460
rect 675482 652216 675538 652225
rect 675482 652151 675538 652160
rect 675404 651681 675432 651848
rect 675390 651672 675446 651681
rect 675390 651607 675446 651616
rect 675404 649602 675432 650012
rect 675392 649596 675444 649602
rect 675392 649538 675444 649544
rect 675404 648961 675432 649468
rect 675390 648952 675446 648961
rect 675390 648887 675446 648896
rect 675772 648689 675800 648788
rect 675758 648680 675814 648689
rect 675758 648615 675814 648624
rect 675496 647766 675524 648176
rect 675484 647760 675536 647766
rect 675484 647702 675536 647708
rect 674748 647352 674800 647358
rect 674748 647294 674800 647300
rect 674748 647216 674800 647222
rect 674748 647158 674800 647164
rect 674656 644632 674708 644638
rect 674656 644574 674708 644580
rect 674668 638602 674696 644574
rect 674760 641918 674788 647158
rect 675404 645454 675432 645660
rect 675392 645448 675444 645454
rect 675392 645390 675444 645396
rect 675404 644638 675432 645116
rect 675392 644632 675444 644638
rect 675392 644574 675444 644580
rect 675404 644162 675432 644475
rect 675392 644156 675444 644162
rect 675392 644098 675444 644104
rect 675404 643414 675432 643824
rect 675392 643408 675444 643414
rect 675392 643350 675444 643356
rect 675404 642122 675432 642635
rect 675392 642116 675444 642122
rect 675392 642058 675444 642064
rect 674748 641912 674800 641918
rect 674748 641854 674800 641860
rect 675392 641912 675444 641918
rect 675392 641854 675444 641860
rect 674748 641708 674800 641714
rect 674748 641650 674800 641656
rect 674760 638722 674788 641650
rect 675404 641444 675432 641854
rect 675404 640286 675432 640795
rect 675392 640280 675444 640286
rect 675392 640222 675444 640228
rect 674748 638716 674800 638722
rect 674748 638658 674800 638664
rect 675208 638716 675260 638722
rect 675208 638658 675260 638664
rect 674668 638574 674788 638602
rect 674656 638444 674708 638450
rect 674656 638386 674708 638392
rect 674564 624300 674616 624306
rect 674564 624242 674616 624248
rect 674564 603084 674616 603090
rect 674564 603026 674616 603032
rect 674576 596902 674604 603026
rect 674564 596896 674616 596902
rect 674564 596838 674616 596844
rect 674472 596828 674524 596834
rect 674472 596770 674524 596776
rect 674392 596686 674604 596714
rect 674472 596624 674524 596630
rect 674472 596566 674524 596572
rect 674380 595332 674432 595338
rect 674380 595274 674432 595280
rect 674392 583982 674420 595274
rect 674380 583976 674432 583982
rect 674380 583918 674432 583924
rect 674380 583704 674432 583710
rect 674380 583646 674432 583652
rect 674288 531140 674340 531146
rect 674288 531082 674340 531088
rect 674392 529514 674420 583646
rect 674484 576842 674512 596566
rect 674576 593094 674604 596686
rect 674564 593088 674616 593094
rect 674564 593030 674616 593036
rect 674668 583982 674696 638386
rect 674760 638246 674788 638574
rect 674748 638240 674800 638246
rect 674748 638182 674800 638188
rect 675220 637566 675248 638658
rect 675496 638450 675524 638928
rect 675484 638444 675536 638450
rect 675484 638386 675536 638392
rect 675484 638240 675536 638246
rect 675484 638182 675536 638188
rect 675208 637560 675260 637566
rect 675208 637502 675260 637508
rect 675496 608841 675524 638182
rect 675668 638172 675720 638178
rect 675668 638114 675720 638120
rect 675482 608832 675538 608841
rect 675680 608802 675708 638114
rect 679164 637900 679216 637906
rect 679164 637842 679216 637848
rect 679072 637560 679124 637566
rect 679072 637502 679124 637508
rect 678978 626104 679034 626113
rect 678978 626039 679034 626048
rect 676126 625696 676182 625705
rect 676126 625631 676182 625640
rect 676034 625152 676090 625161
rect 676034 625087 676090 625096
rect 676048 624306 676076 625087
rect 676036 624300 676088 624306
rect 676036 624242 676088 624248
rect 676140 624034 676168 625631
rect 676310 625288 676366 625297
rect 676310 625223 676366 625232
rect 676218 624472 676274 624481
rect 676218 624407 676274 624416
rect 676128 624028 676180 624034
rect 676128 623970 676180 623976
rect 676036 623960 676088 623966
rect 676034 623928 676036 623937
rect 676088 623928 676090 623937
rect 676034 623863 676090 623872
rect 676232 623830 676260 624407
rect 676324 623898 676352 625223
rect 678992 624170 679020 626039
rect 679084 624481 679112 637502
rect 679070 624472 679126 624481
rect 679070 624407 679126 624416
rect 678980 624164 679032 624170
rect 678980 624106 679032 624112
rect 676312 623892 676364 623898
rect 676312 623834 676364 623840
rect 676220 623824 676272 623830
rect 676220 623766 676272 623772
rect 676036 623756 676088 623762
rect 676036 623698 676088 623704
rect 676048 621489 676076 623698
rect 679176 623665 679204 637842
rect 708512 627360 708564 627366
rect 704168 627298 704504 627314
rect 708564 627308 708768 627314
rect 708512 627302 708768 627308
rect 704168 627292 704516 627298
rect 704168 627286 704464 627292
rect 704464 627234 704516 627240
rect 708420 627292 708472 627298
rect 708524 627286 708768 627302
rect 708420 627234 708472 627240
rect 704372 627224 704424 627230
rect 703556 627150 703708 627178
rect 707500 627224 707552 627230
rect 704372 627166 704424 627172
rect 703556 626686 703584 627150
rect 704384 626906 704412 627166
rect 704628 627150 704964 627178
rect 705088 627150 705424 627178
rect 705548 627150 705884 627178
rect 706008 627150 706344 627178
rect 704168 626878 704412 626906
rect 704936 626822 704964 627150
rect 705292 627088 705344 627094
rect 705292 627030 705344 627036
rect 705304 626906 705332 627030
rect 705088 626878 705332 626906
rect 705396 626890 705424 627150
rect 705752 627088 705804 627094
rect 705752 627030 705804 627036
rect 705764 626906 705792 627030
rect 705856 627026 705884 627150
rect 706212 627088 706264 627094
rect 706212 627030 706264 627036
rect 705844 627020 705896 627026
rect 705844 626962 705896 626968
rect 706224 626906 706252 627030
rect 706316 626958 706344 627150
rect 706592 627150 706928 627178
rect 707052 627162 707388 627178
rect 707552 627172 707848 627178
rect 707500 627166 707848 627172
rect 707040 627156 707388 627162
rect 706592 627094 706620 627150
rect 707092 627150 707388 627156
rect 707512 627150 707848 627166
rect 708064 627150 708308 627178
rect 707040 627098 707092 627104
rect 706580 627088 706632 627094
rect 706580 627030 706632 627036
rect 705384 626884 705436 626890
rect 705548 626878 705792 626906
rect 706008 626878 706252 626906
rect 706304 626952 706356 626958
rect 706304 626894 706356 626900
rect 706454 626892 706482 627028
rect 707040 627020 707092 627026
rect 707040 626962 707092 626968
rect 706580 626952 706632 626958
rect 707052 626906 707080 626962
rect 706632 626900 706928 626906
rect 706580 626894 706928 626900
rect 706592 626878 706928 626894
rect 707052 626878 707388 626906
rect 707512 626890 707848 626906
rect 708064 626890 708092 627150
rect 708432 626906 708460 627234
rect 708984 627150 709228 627178
rect 707500 626884 707848 626890
rect 705384 626826 705436 626832
rect 707552 626878 707848 626884
rect 708052 626884 708104 626890
rect 707500 626826 707552 626832
rect 708432 626878 708768 626906
rect 708052 626826 708104 626832
rect 704924 626816 704976 626822
rect 704628 626754 704872 626770
rect 704924 626758 704976 626764
rect 707960 626816 708012 626822
rect 708012 626764 708308 626770
rect 707960 626758 708308 626764
rect 704628 626748 704884 626754
rect 704628 626742 704832 626748
rect 707972 626742 708308 626758
rect 708984 626754 709012 627150
rect 708972 626748 709024 626754
rect 704832 626690 704884 626696
rect 708972 626690 709024 626696
rect 703544 626680 703596 626686
rect 708880 626680 708932 626686
rect 703544 626622 703596 626628
rect 703708 626618 704044 626634
rect 708932 626628 709228 626634
rect 708880 626622 709228 626628
rect 703708 626612 704056 626618
rect 703708 626606 704004 626612
rect 708892 626606 709228 626622
rect 704004 626554 704056 626560
rect 679162 623656 679218 623665
rect 679162 623591 679218 623600
rect 678978 623248 679034 623257
rect 678978 623183 679034 623192
rect 676218 622024 676274 622033
rect 676218 621959 676274 621968
rect 676034 621480 676090 621489
rect 676034 621415 676090 621424
rect 676232 621110 676260 621959
rect 676220 621104 676272 621110
rect 676220 621046 676272 621052
rect 678992 621042 679020 623183
rect 678980 621036 679032 621042
rect 678980 620978 679032 620984
rect 676036 620968 676088 620974
rect 676036 620910 676088 620916
rect 676048 619857 676076 620910
rect 676128 620900 676180 620906
rect 676128 620842 676180 620848
rect 676140 620401 676168 620842
rect 676126 620392 676182 620401
rect 676126 620327 676182 620336
rect 676034 619848 676090 619857
rect 676034 619783 676090 619792
rect 676036 618248 676088 618254
rect 676034 618216 676036 618225
rect 676088 618216 676090 618225
rect 676034 618151 676090 618160
rect 676220 617976 676272 617982
rect 676218 617944 676220 617953
rect 676272 617944 676274 617953
rect 676218 617879 676274 617888
rect 676220 616752 676272 616758
rect 676218 616720 676220 616729
rect 676272 616720 676274 616729
rect 676218 616655 676274 616664
rect 679254 615904 679310 615913
rect 679254 615839 679310 615848
rect 679268 615505 679296 615839
rect 678978 615496 679034 615505
rect 678978 615431 679034 615440
rect 679254 615496 679310 615505
rect 679254 615431 679310 615440
rect 678992 615097 679020 615431
rect 678978 615088 679034 615097
rect 678978 615023 679034 615032
rect 679268 614786 679296 615431
rect 679256 614780 679308 614786
rect 679256 614722 679308 614728
rect 675482 608767 675538 608776
rect 675668 608796 675720 608802
rect 675668 608738 675720 608744
rect 675680 607617 675708 608124
rect 675666 607608 675722 607617
rect 675666 607543 675722 607552
rect 675772 607345 675800 607479
rect 675758 607336 675814 607345
rect 675758 607271 675814 607280
rect 675404 606529 675432 606832
rect 675390 606520 675446 606529
rect 675390 606455 675446 606464
rect 675404 604761 675432 604996
rect 675390 604752 675446 604761
rect 675390 604687 675446 604696
rect 675496 604353 675524 604452
rect 675482 604344 675538 604353
rect 675482 604279 675538 604288
rect 675496 603537 675524 603772
rect 675482 603528 675538 603537
rect 675482 603463 675538 603472
rect 675772 602993 675800 603160
rect 675758 602984 675814 602993
rect 675758 602919 675814 602928
rect 675496 600438 675524 600644
rect 675484 600432 675536 600438
rect 675484 600374 675536 600380
rect 675496 599622 675524 600100
rect 674748 599616 674800 599622
rect 674748 599558 674800 599564
rect 675484 599616 675536 599622
rect 675484 599558 675536 599564
rect 674564 583976 674616 583982
rect 674564 583918 674616 583924
rect 674656 583976 674708 583982
rect 674656 583918 674708 583924
rect 674576 583794 674604 583918
rect 674576 583766 674696 583794
rect 674760 583778 674788 599558
rect 675404 599146 675432 599488
rect 675392 599140 675444 599146
rect 675392 599082 675444 599088
rect 675496 598466 675524 598808
rect 675484 598460 675536 598466
rect 675484 598402 675536 598408
rect 675404 597174 675432 597652
rect 675392 597168 675444 597174
rect 675392 597110 675444 597116
rect 675392 596896 675444 596902
rect 675392 596838 675444 596844
rect 675404 596428 675432 596838
rect 675404 595338 675432 595816
rect 675392 595332 675444 595338
rect 675392 595274 675444 595280
rect 675496 593706 675524 593980
rect 675208 593700 675260 593706
rect 675208 593642 675260 593648
rect 675484 593700 675536 593706
rect 675484 593642 675536 593648
rect 674564 583704 674616 583710
rect 674564 583646 674616 583652
rect 674472 576836 674524 576842
rect 674472 576778 674524 576784
rect 674472 548888 674524 548894
rect 674472 548830 674524 548836
rect 674380 529508 674432 529514
rect 674380 529450 674432 529456
rect 674484 487898 674512 548830
rect 674576 529922 674604 583646
rect 674668 574094 674696 583766
rect 674748 583772 674800 583778
rect 674748 583714 674800 583720
rect 675220 583710 675248 593642
rect 675576 593088 675628 593094
rect 675576 593030 675628 593036
rect 675392 583976 675444 583982
rect 675392 583918 675444 583924
rect 675208 583704 675260 583710
rect 675208 583646 675260 583652
rect 675404 574569 675432 583918
rect 675484 583772 675536 583778
rect 675484 583714 675536 583720
rect 675390 574560 675446 574569
rect 675390 574495 675446 574504
rect 674668 574066 674788 574094
rect 674656 548276 674708 548282
rect 674656 548218 674708 548224
rect 674564 529916 674616 529922
rect 674564 529858 674616 529864
rect 674472 487892 674524 487898
rect 674472 487834 674524 487840
rect 674196 487144 674248 487150
rect 674196 487086 674248 487092
rect 674668 485790 674696 548218
rect 674760 532710 674788 574066
rect 675496 564505 675524 583714
rect 675588 575385 675616 593030
rect 678980 587920 679032 587926
rect 678980 587862 679032 587868
rect 676126 580952 676182 580961
rect 676126 580887 676182 580896
rect 676036 580236 676088 580242
rect 676036 580178 676088 580184
rect 676048 579873 676076 580178
rect 676140 579970 676168 580887
rect 676310 580544 676366 580553
rect 676310 580479 676366 580488
rect 676218 580136 676274 580145
rect 676218 580071 676220 580080
rect 676272 580071 676274 580080
rect 676220 580042 676272 580048
rect 676128 579964 676180 579970
rect 676128 579906 676180 579912
rect 676034 579864 676090 579873
rect 676324 579834 676352 580479
rect 676034 579799 676090 579808
rect 676312 579828 676364 579834
rect 676312 579770 676364 579776
rect 678992 579329 679020 587862
rect 703452 584180 703504 584186
rect 703452 584122 703504 584128
rect 709340 584180 709392 584186
rect 709340 584122 709392 584128
rect 703464 581754 703492 584122
rect 709352 582162 709380 584122
rect 703708 582146 704044 582162
rect 703708 582140 704056 582146
rect 703708 582134 704004 582140
rect 704004 582082 704056 582088
rect 708880 582140 708932 582146
rect 709228 582134 709380 582162
rect 708880 582082 708932 582088
rect 708052 582072 708104 582078
rect 704628 582010 704964 582026
rect 708104 582020 708308 582026
rect 708052 582014 708308 582020
rect 704628 582004 704976 582010
rect 704628 581998 704924 582004
rect 704924 581946 704976 581952
rect 707960 582004 708012 582010
rect 708064 581998 708308 582014
rect 707960 581946 708012 581952
rect 704832 581936 704884 581942
rect 704168 581862 704504 581890
rect 707040 581936 707092 581942
rect 704832 581878 704884 581884
rect 703464 581726 703708 581754
rect 704476 581534 704504 581862
rect 704844 581754 704872 581878
rect 705088 581862 705424 581890
rect 705548 581862 705884 581890
rect 706008 581862 706344 581890
rect 704628 581726 704872 581754
rect 705396 581670 705424 581862
rect 705752 581800 705804 581806
rect 705548 581748 705752 581754
rect 705548 581742 705804 581748
rect 705548 581726 705792 581742
rect 705856 581738 705884 581862
rect 706316 581806 706344 581862
rect 706212 581800 706264 581806
rect 706008 581748 706212 581754
rect 706008 581742 706264 581748
rect 706304 581800 706356 581806
rect 706304 581742 706356 581748
rect 705844 581732 705896 581738
rect 706008 581726 706252 581742
rect 706454 581740 706482 581876
rect 706684 581874 706928 581890
rect 707092 581884 707388 581890
rect 707040 581878 707388 581884
rect 706672 581868 706928 581874
rect 706724 581862 706928 581868
rect 707052 581862 707388 581878
rect 707604 581862 707848 581890
rect 706672 581810 706724 581816
rect 706580 581800 706632 581806
rect 706632 581748 706928 581754
rect 706580 581742 706928 581748
rect 706592 581726 706928 581742
rect 707052 581738 707388 581754
rect 707604 581738 707632 581862
rect 707972 581754 708000 581946
rect 708524 581862 708768 581890
rect 707040 581732 707388 581738
rect 705844 581674 705896 581680
rect 707092 581726 707388 581732
rect 707592 581732 707644 581738
rect 707040 581674 707092 581680
rect 707972 581726 708308 581754
rect 707592 581674 707644 581680
rect 705384 581664 705436 581670
rect 705088 581602 705332 581618
rect 705384 581606 705436 581612
rect 707500 581664 707552 581670
rect 707552 581612 707848 581618
rect 707500 581606 707848 581612
rect 705088 581596 705344 581602
rect 705088 581590 705292 581596
rect 707512 581590 707848 581606
rect 708524 581602 708552 581862
rect 708892 581754 708920 582082
rect 708892 581726 709228 581754
rect 708512 581596 708564 581602
rect 705292 581538 705344 581544
rect 708512 581538 708564 581544
rect 704464 581528 704516 581534
rect 704168 581466 704412 581482
rect 704464 581470 704516 581476
rect 708420 581528 708472 581534
rect 708472 581476 708768 581482
rect 708420 581470 708768 581476
rect 704168 581460 704424 581466
rect 704168 581454 704372 581460
rect 708432 581454 708768 581470
rect 704372 581402 704424 581408
rect 676218 579320 676274 579329
rect 676218 579255 676220 579264
rect 676272 579255 676274 579264
rect 678978 579320 679034 579329
rect 678978 579255 679034 579264
rect 676220 579226 676272 579232
rect 676218 578504 676274 578513
rect 676218 578439 676220 578448
rect 676272 578439 676274 578448
rect 676220 578410 676272 578416
rect 676218 577688 676274 577697
rect 676218 577623 676220 577632
rect 676272 577623 676274 577632
rect 676220 577594 676272 577600
rect 676218 577280 676274 577289
rect 676218 577215 676274 577224
rect 676232 577182 676260 577215
rect 676220 577176 676272 577182
rect 676220 577118 676272 577124
rect 676034 577008 676090 577017
rect 676034 576943 676036 576952
rect 676088 576943 676090 576952
rect 676036 576914 676088 576920
rect 676036 576836 676088 576842
rect 676036 576778 676088 576784
rect 676048 576201 676076 576778
rect 676034 576192 676090 576201
rect 676034 576127 676090 576136
rect 676036 576088 676088 576094
rect 676036 576030 676088 576036
rect 675574 575376 675630 575385
rect 675574 575311 675630 575320
rect 676048 574977 676076 576030
rect 676034 574968 676090 574977
rect 676034 574903 676090 574912
rect 676036 573640 676088 573646
rect 676036 573582 676088 573588
rect 676048 572937 676076 573582
rect 676034 572928 676090 572937
rect 676034 572863 676090 572872
rect 676036 572824 676088 572830
rect 676036 572766 676088 572772
rect 676048 572529 676076 572766
rect 676034 572520 676090 572529
rect 676034 572455 676090 572464
rect 676036 572416 676088 572422
rect 676036 572358 676088 572364
rect 676048 572121 676076 572358
rect 676034 572112 676090 572121
rect 676034 572047 676090 572056
rect 678978 570752 679034 570761
rect 678978 570687 679034 570696
rect 678992 570353 679020 570687
rect 678978 570344 679034 570353
rect 678978 570279 679034 570288
rect 684498 570344 684554 570353
rect 684498 570279 684554 570288
rect 678992 568614 679020 570279
rect 684512 569945 684540 570279
rect 684498 569936 684554 569945
rect 684498 569871 684554 569880
rect 678980 568608 679032 568614
rect 678980 568550 679032 568556
rect 675482 564496 675538 564505
rect 675482 564431 675538 564440
rect 675496 562465 675524 562904
rect 675482 562456 675538 562465
rect 675482 562391 675538 562400
rect 675772 562057 675800 562292
rect 675758 562048 675814 562057
rect 675758 561983 675814 561992
rect 675496 561241 675524 561612
rect 675482 561232 675538 561241
rect 675482 561167 675538 561176
rect 675496 559570 675524 559776
rect 675484 559564 675536 559570
rect 675484 559506 675536 559512
rect 675404 558793 675432 559232
rect 675390 558784 675446 558793
rect 675390 558719 675446 558728
rect 675772 558385 675800 558620
rect 675758 558376 675814 558385
rect 675758 558311 675814 558320
rect 675772 557569 675800 557940
rect 675758 557560 675814 557569
rect 675758 557495 675814 557504
rect 675300 556164 675352 556170
rect 675300 556106 675352 556112
rect 675312 551253 675340 556106
rect 675404 555286 675432 555492
rect 675392 555280 675444 555286
rect 675392 555222 675444 555228
rect 675404 554606 675432 554919
rect 675392 554600 675444 554606
rect 675392 554542 675444 554548
rect 675404 553790 675432 554268
rect 675392 553784 675444 553790
rect 675392 553726 675444 553732
rect 675404 553246 675432 553656
rect 675392 553240 675444 553246
rect 675392 553182 675444 553188
rect 675404 551954 675432 552432
rect 675392 551948 675444 551954
rect 675392 551890 675444 551896
rect 675312 551225 675418 551253
rect 675312 550582 675418 550610
rect 675312 548894 675340 550582
rect 675300 548888 675352 548894
rect 675300 548830 675352 548836
rect 675312 548746 675418 548774
rect 675312 548282 675340 548746
rect 675300 548276 675352 548282
rect 675300 548218 675352 548224
rect 679072 546304 679124 546310
rect 679072 546246 679124 546252
rect 676218 535936 676274 535945
rect 676218 535871 676274 535880
rect 676232 535770 676260 535871
rect 676220 535764 676272 535770
rect 676034 535732 676090 535741
rect 676220 535706 676272 535712
rect 676034 535667 676090 535676
rect 676048 535634 676076 535667
rect 676036 535628 676088 535634
rect 676036 535570 676088 535576
rect 678978 535120 679034 535129
rect 678978 535055 679034 535064
rect 676036 534948 676088 534954
rect 676034 534916 676036 534925
rect 676088 534916 676090 534925
rect 676034 534851 676090 534860
rect 676126 534304 676182 534313
rect 676126 534239 676182 534248
rect 676036 533316 676088 533322
rect 676034 533284 676036 533293
rect 676088 533284 676090 533293
rect 676034 533219 676090 533228
rect 675942 532876 675998 532885
rect 675852 532840 675904 532846
rect 676140 532846 676168 534239
rect 678992 532914 679020 535055
rect 679084 534313 679112 546246
rect 703452 537192 703504 537198
rect 703452 537134 703504 537140
rect 703464 536738 703492 537134
rect 703556 537130 703708 537146
rect 708984 537130 709228 537146
rect 703544 537124 703708 537130
rect 703596 537118 703708 537124
rect 708880 537124 708932 537130
rect 703544 537066 703596 537072
rect 708880 537066 708932 537072
rect 708972 537124 709228 537130
rect 709024 537118 709228 537124
rect 708972 537066 709024 537072
rect 708052 537056 708104 537062
rect 704628 536994 704964 537010
rect 708104 537004 708308 537010
rect 708052 536998 708308 537004
rect 704628 536988 704976 536994
rect 704628 536982 704924 536988
rect 704924 536930 704976 536936
rect 707960 536988 708012 536994
rect 708064 536982 708308 536998
rect 707960 536930 708012 536936
rect 704832 536920 704884 536926
rect 704168 536846 704504 536874
rect 707040 536920 707092 536926
rect 704832 536862 704884 536868
rect 703464 536710 703708 536738
rect 704476 536518 704504 536846
rect 704844 536738 704872 536862
rect 705088 536846 705424 536874
rect 705548 536846 705884 536874
rect 706008 536846 706344 536874
rect 704628 536710 704872 536738
rect 705396 536654 705424 536846
rect 705752 536784 705804 536790
rect 705548 536732 705752 536738
rect 705548 536726 705804 536732
rect 705548 536710 705792 536726
rect 705856 536722 705884 536846
rect 706316 536790 706344 536846
rect 706212 536784 706264 536790
rect 706008 536732 706212 536738
rect 706008 536726 706264 536732
rect 706304 536784 706356 536790
rect 706304 536726 706356 536732
rect 705844 536716 705896 536722
rect 706008 536710 706252 536726
rect 706454 536724 706482 536860
rect 706684 536858 706928 536874
rect 707092 536868 707388 536874
rect 707040 536862 707388 536868
rect 706672 536852 706928 536858
rect 706724 536846 706928 536852
rect 707052 536846 707388 536862
rect 707604 536846 707848 536874
rect 706672 536794 706724 536800
rect 706580 536784 706632 536790
rect 706632 536732 706928 536738
rect 706580 536726 706928 536732
rect 706592 536710 706928 536726
rect 707052 536722 707388 536738
rect 707604 536722 707632 536846
rect 707972 536738 708000 536930
rect 708524 536846 708768 536874
rect 707040 536716 707388 536722
rect 705844 536658 705896 536664
rect 707092 536710 707388 536716
rect 707592 536716 707644 536722
rect 707040 536658 707092 536664
rect 707972 536710 708308 536738
rect 707592 536658 707644 536664
rect 705384 536648 705436 536654
rect 705088 536586 705332 536602
rect 705384 536590 705436 536596
rect 707500 536648 707552 536654
rect 707552 536596 707848 536602
rect 707500 536590 707848 536596
rect 705088 536580 705344 536586
rect 705088 536574 705292 536580
rect 707512 536574 707848 536590
rect 708524 536586 708552 536846
rect 708892 536738 708920 537066
rect 708892 536710 709228 536738
rect 708512 536580 708564 536586
rect 705292 536522 705344 536528
rect 708512 536522 708564 536528
rect 704464 536512 704516 536518
rect 704168 536450 704412 536466
rect 704464 536454 704516 536460
rect 708420 536512 708472 536518
rect 708472 536460 708768 536466
rect 708420 536454 708768 536460
rect 704168 536444 704424 536450
rect 704168 536438 704372 536444
rect 708432 536438 708768 536454
rect 704372 536386 704424 536392
rect 679070 534304 679126 534313
rect 679070 534239 679126 534248
rect 679070 533488 679126 533497
rect 679070 533423 679126 533432
rect 678980 532908 679032 532914
rect 678980 532850 679032 532856
rect 675942 532811 675998 532820
rect 676128 532840 676180 532846
rect 675852 532782 675904 532788
rect 674748 532704 674800 532710
rect 674748 532646 674800 532652
rect 675758 532060 675814 532069
rect 675758 531995 675814 532004
rect 675666 488880 675722 488889
rect 675666 488815 675722 488824
rect 675576 488572 675628 488578
rect 675576 488514 675628 488520
rect 675208 488096 675260 488102
rect 675206 488064 675208 488073
rect 675260 488064 675262 488073
rect 675206 487999 675262 488008
rect 674656 485784 674708 485790
rect 674656 485726 674708 485732
rect 674012 485512 674064 485518
rect 674012 485454 674064 485460
rect 673920 483880 673972 483886
rect 673920 483822 673972 483828
rect 673644 482996 673696 483002
rect 673644 482938 673696 482944
rect 673460 482928 673512 482934
rect 673460 482870 673512 482876
rect 675588 478922 675616 488514
rect 675576 478916 675628 478922
rect 675576 478858 675628 478864
rect 675680 419534 675708 488815
rect 675772 488481 675800 531995
rect 675864 490929 675892 532782
rect 675956 496814 675984 532811
rect 676128 532782 676180 532788
rect 676036 532704 676088 532710
rect 676036 532646 676088 532652
rect 676218 532672 676274 532681
rect 676048 531253 676076 532646
rect 676218 532607 676220 532616
rect 676272 532607 676274 532616
rect 676220 532578 676272 532584
rect 676034 531244 676090 531253
rect 676034 531179 676090 531188
rect 676036 531140 676088 531146
rect 676036 531082 676088 531088
rect 676048 530029 676076 531082
rect 676034 530020 676090 530029
rect 676034 529955 676090 529964
rect 676036 529916 676088 529922
rect 676036 529858 676088 529864
rect 676048 529621 676076 529858
rect 676034 529612 676090 529621
rect 676034 529547 676090 529556
rect 676036 529508 676088 529514
rect 676036 529450 676088 529456
rect 676048 527989 676076 529450
rect 676034 527980 676090 527989
rect 676034 527915 676090 527924
rect 676036 527876 676088 527882
rect 676036 527818 676088 527824
rect 676048 527581 676076 527818
rect 676034 527572 676090 527581
rect 676034 527507 676090 527516
rect 676036 527128 676088 527134
rect 676036 527070 676088 527076
rect 676048 526357 676076 527070
rect 676034 526348 676090 526357
rect 676034 526283 676090 526292
rect 678978 525736 679034 525745
rect 678978 525671 679034 525680
rect 678992 525337 679020 525671
rect 678978 525328 679034 525337
rect 678978 525263 679034 525272
rect 678992 524482 679020 525263
rect 678980 524476 679032 524482
rect 678980 524418 679032 524424
rect 679084 524414 679112 533423
rect 684590 525328 684646 525337
rect 684590 525263 684646 525272
rect 684604 524929 684632 525263
rect 684590 524920 684646 524929
rect 684590 524855 684646 524864
rect 677508 524408 677560 524414
rect 677508 524350 677560 524356
rect 679072 524408 679124 524414
rect 679072 524350 679124 524356
rect 675956 496786 676168 496814
rect 676034 492144 676090 492153
rect 676034 492079 676090 492088
rect 675942 491736 675998 491745
rect 676048 491706 676076 492079
rect 675942 491671 675998 491680
rect 676036 491700 676088 491706
rect 675956 491434 675984 491671
rect 676036 491642 676088 491648
rect 676036 491564 676088 491570
rect 676036 491506 676088 491512
rect 675944 491428 675996 491434
rect 675944 491370 675996 491376
rect 676048 491337 676076 491506
rect 676034 491328 676090 491337
rect 676034 491263 676090 491272
rect 675850 490920 675906 490929
rect 675850 490855 675906 490864
rect 675942 490512 675998 490521
rect 675942 490447 675998 490456
rect 675850 489696 675906 489705
rect 675850 489631 675906 489640
rect 675758 488472 675814 488481
rect 675758 488407 675814 488416
rect 675588 419506 675708 419534
rect 674656 401260 674708 401266
rect 674656 401202 674708 401208
rect 674380 399492 674432 399498
rect 674380 399434 674432 399440
rect 673736 397656 673788 397662
rect 673736 397598 673788 397604
rect 673460 396636 673512 396642
rect 673460 396578 673512 396584
rect 672908 392080 672960 392086
rect 672908 392022 672960 392028
rect 672814 278488 672870 278497
rect 672814 278423 672870 278432
rect 672816 256896 672868 256902
rect 672816 256838 672868 256844
rect 672722 148200 672778 148209
rect 672722 148135 672778 148144
rect 672448 130892 672500 130898
rect 672448 130834 672500 130840
rect 672354 117736 672410 117745
rect 672354 117671 672410 117680
rect 672262 109304 672318 109313
rect 672262 109239 672318 109248
rect 672460 105913 672488 130834
rect 672828 127945 672856 256838
rect 672920 143177 672948 392022
rect 673472 372094 673500 396578
rect 673552 395412 673604 395418
rect 673552 395354 673604 395360
rect 673564 376922 673592 395354
rect 673644 394868 673696 394874
rect 673644 394810 673696 394816
rect 673656 378214 673684 394810
rect 673748 379506 673776 397598
rect 674288 397588 674340 397594
rect 674288 397530 674340 397536
rect 673828 394188 673880 394194
rect 673828 394130 673880 394136
rect 673736 379500 673788 379506
rect 673736 379442 673788 379448
rect 673644 378208 673696 378214
rect 673644 378150 673696 378156
rect 673840 378010 673868 394130
rect 674012 392012 674064 392018
rect 674012 391954 674064 391960
rect 673828 378004 673880 378010
rect 673828 377946 673880 377952
rect 674024 376990 674052 391954
rect 674012 376984 674064 376990
rect 674012 376926 674064 376932
rect 673552 376916 673604 376922
rect 673552 376858 673604 376864
rect 674300 373930 674328 397530
rect 674392 382362 674420 399434
rect 674472 398268 674524 398274
rect 674472 398210 674524 398216
rect 674484 385014 674512 398210
rect 674564 390516 674616 390522
rect 674564 390458 674616 390464
rect 674472 385008 674524 385014
rect 674472 384950 674524 384956
rect 674380 382356 674432 382362
rect 674380 382298 674432 382304
rect 674288 373924 674340 373930
rect 674288 373866 674340 373872
rect 673460 372088 673512 372094
rect 673460 372030 673512 372036
rect 674576 370734 674604 390458
rect 674564 370728 674616 370734
rect 674564 370670 674616 370676
rect 674668 361574 674696 401202
rect 675588 401033 675616 419506
rect 675864 401849 675892 489631
rect 675956 488578 675984 490447
rect 676140 490210 676168 496786
rect 677520 491298 677548 524350
rect 704372 493128 704424 493134
rect 704177 493076 704372 493082
rect 704177 493070 704424 493076
rect 704177 493054 704412 493070
rect 708432 493066 708768 493082
rect 704464 493060 704516 493066
rect 704464 493002 704516 493008
rect 708420 493060 708768 493066
rect 708472 493054 708768 493060
rect 708420 493002 708472 493008
rect 703556 492918 703708 492946
rect 703556 492386 703584 492918
rect 704476 492674 704504 493002
rect 705384 492992 705436 492998
rect 704637 492918 704964 492946
rect 705097 492940 705384 492946
rect 708512 492992 708564 492998
rect 705097 492934 705436 492940
rect 705097 492918 705424 492934
rect 705557 492918 705884 492946
rect 706017 492918 706344 492946
rect 704168 492646 704504 492674
rect 704832 492584 704884 492590
rect 703708 492522 703952 492538
rect 704628 492532 704832 492538
rect 704628 492526 704884 492532
rect 703708 492516 703964 492522
rect 703708 492510 703912 492516
rect 704628 492510 704872 492526
rect 703912 492458 703964 492464
rect 704936 492454 704964 492918
rect 705752 492856 705804 492862
rect 705752 492798 705804 492804
rect 705764 492674 705792 492798
rect 705856 492794 705884 492918
rect 706212 492856 706264 492862
rect 706212 492798 706264 492804
rect 705844 492788 705896 492794
rect 705844 492730 705896 492736
rect 706224 492674 706252 492798
rect 706316 492726 706344 492918
rect 706454 492796 706482 492932
rect 706592 492918 706928 492946
rect 707052 492930 707388 492946
rect 707040 492924 707388 492930
rect 706592 492862 706620 492918
rect 707092 492918 707388 492924
rect 707512 492918 707848 492946
rect 707972 492918 708308 492946
rect 708512 492934 708564 492940
rect 707040 492866 707092 492872
rect 706580 492856 706632 492862
rect 706580 492798 706632 492804
rect 707040 492788 707092 492794
rect 707040 492730 707092 492736
rect 705088 492658 705424 492674
rect 705088 492652 705436 492658
rect 705088 492646 705384 492652
rect 705548 492646 705792 492674
rect 706008 492646 706252 492674
rect 706304 492720 706356 492726
rect 706304 492662 706356 492668
rect 706580 492720 706632 492726
rect 707052 492674 707080 492730
rect 706632 492668 706928 492674
rect 706580 492662 706928 492668
rect 706592 492646 706928 492662
rect 707052 492646 707388 492674
rect 707512 492658 707540 492918
rect 707592 492856 707644 492862
rect 707592 492798 707644 492804
rect 707604 492674 707632 492798
rect 707500 492652 707552 492658
rect 705384 492594 705436 492600
rect 707604 492646 707848 492674
rect 707500 492594 707552 492600
rect 707972 492590 708000 492918
rect 708524 492674 708552 492934
rect 708892 492918 709228 492946
rect 708524 492646 708768 492674
rect 707960 492584 708012 492590
rect 707960 492526 708012 492532
rect 708892 492522 708920 492918
rect 708880 492516 708932 492522
rect 708880 492458 708932 492464
rect 704924 492448 704976 492454
rect 704924 492390 704976 492396
rect 707960 492448 708012 492454
rect 708012 492396 708308 492402
rect 707960 492390 708308 492396
rect 703544 492380 703596 492386
rect 707972 492374 708308 492390
rect 708892 492386 709228 492402
rect 708880 492380 709228 492386
rect 703544 492322 703596 492328
rect 708932 492374 709228 492380
rect 708880 492322 708932 492328
rect 676220 491292 676272 491298
rect 676220 491234 676272 491240
rect 677508 491292 677560 491298
rect 677508 491234 677560 491240
rect 676128 490204 676180 490210
rect 676128 490146 676180 490152
rect 676034 490104 676090 490113
rect 676232 490090 676260 491234
rect 676090 490062 676260 490090
rect 676034 490039 676090 490048
rect 676036 490000 676088 490006
rect 676036 489942 676088 489948
rect 676048 489297 676076 489942
rect 676034 489288 676090 489297
rect 676034 489223 676090 489232
rect 675944 488572 675996 488578
rect 675944 488514 675996 488520
rect 676034 488064 676090 488073
rect 676090 488022 676168 488050
rect 676034 487999 676090 488008
rect 676036 487892 676088 487898
rect 676036 487834 676088 487840
rect 675944 487484 675996 487490
rect 675944 487426 675996 487432
rect 675956 486441 675984 487426
rect 676048 487257 676076 487834
rect 676034 487248 676090 487257
rect 676034 487183 676090 487192
rect 676036 487144 676088 487150
rect 676036 487086 676088 487092
rect 675942 486432 675998 486441
rect 675942 486367 675998 486376
rect 676048 486033 676076 487086
rect 676034 486024 676090 486033
rect 676034 485959 676090 485968
rect 676036 485784 676088 485790
rect 676036 485726 676088 485732
rect 676048 485625 676076 485726
rect 676034 485616 676090 485625
rect 676034 485551 676090 485560
rect 676036 485512 676088 485518
rect 676036 485454 676088 485460
rect 676048 483993 676076 485454
rect 676034 483984 676090 483993
rect 676034 483919 676090 483928
rect 676036 483880 676088 483886
rect 676036 483822 676088 483828
rect 676048 483585 676076 483822
rect 676034 483576 676090 483585
rect 676034 483511 676090 483520
rect 676036 482996 676088 483002
rect 676036 482938 676088 482944
rect 675944 482928 675996 482934
rect 675944 482870 675996 482876
rect 675956 482769 675984 482870
rect 675942 482760 675998 482769
rect 675942 482695 675998 482704
rect 676048 482361 676076 482938
rect 676034 482352 676090 482361
rect 676034 482287 676090 482296
rect 676034 481944 676090 481953
rect 676034 481879 676090 481888
rect 675942 481536 675998 481545
rect 675942 481471 675998 481480
rect 675956 480729 675984 481471
rect 676048 481166 676076 481879
rect 676036 481160 676088 481166
rect 676034 481128 676036 481137
rect 676088 481128 676090 481137
rect 676034 481063 676090 481072
rect 675942 480720 675998 480729
rect 675942 480655 675998 480664
rect 676140 480254 676168 488022
rect 676048 480226 676168 480254
rect 675942 403472 675998 403481
rect 675942 403407 675944 403416
rect 675996 403407 675998 403416
rect 675944 403378 675996 403384
rect 675944 403164 675996 403170
rect 675944 403106 675996 403112
rect 675956 403073 675984 403106
rect 675942 403064 675998 403073
rect 675942 402999 675998 403008
rect 675850 401840 675906 401849
rect 675850 401775 675906 401784
rect 675666 401432 675722 401441
rect 675666 401367 675722 401376
rect 675574 401024 675630 401033
rect 675574 400959 675630 400968
rect 674932 397520 674984 397526
rect 674932 397462 674984 397468
rect 674748 390584 674800 390590
rect 674748 390526 674800 390532
rect 674760 370802 674788 390526
rect 674944 383178 674972 397462
rect 675298 396944 675354 396953
rect 675298 396879 675354 396888
rect 675116 395004 675168 395010
rect 675116 394946 675168 394952
rect 675024 394800 675076 394806
rect 675024 394742 675076 394748
rect 674932 383172 674984 383178
rect 674932 383114 674984 383120
rect 675036 381954 675064 394742
rect 675128 382498 675156 394946
rect 675208 394732 675260 394738
rect 675208 394674 675260 394680
rect 675220 384130 675248 394674
rect 675312 385098 675340 396879
rect 675680 390522 675708 401367
rect 675758 400616 675814 400625
rect 675758 400551 675814 400560
rect 675772 390590 675800 400551
rect 676048 400217 676076 480226
rect 676128 478916 676180 478922
rect 676128 478858 676180 478864
rect 676140 402937 676168 478858
rect 703708 404938 704044 404954
rect 708984 404938 709228 404954
rect 703544 404932 703596 404938
rect 703708 404932 704056 404938
rect 703708 404926 704004 404932
rect 703544 404874 703596 404880
rect 704004 404874 704056 404880
rect 708880 404932 708932 404938
rect 708880 404874 708932 404880
rect 708972 404932 709228 404938
rect 709024 404926 709228 404932
rect 708972 404874 709024 404880
rect 703556 404546 703584 404874
rect 708052 404864 708104 404870
rect 704628 404802 704964 404818
rect 708104 404812 708308 404818
rect 708052 404806 708308 404812
rect 704628 404796 704976 404802
rect 704628 404790 704924 404796
rect 704924 404738 704976 404744
rect 707960 404796 708012 404802
rect 708064 404790 708308 404806
rect 707960 404738 708012 404744
rect 704832 404728 704884 404734
rect 704168 404654 704504 404682
rect 707040 404728 707092 404734
rect 704832 404670 704884 404676
rect 703556 404518 703708 404546
rect 704476 404326 704504 404654
rect 704844 404546 704872 404670
rect 705088 404654 705424 404682
rect 705548 404654 705884 404682
rect 706008 404654 706344 404682
rect 704628 404518 704872 404546
rect 705396 404462 705424 404654
rect 705752 404592 705804 404598
rect 705548 404540 705752 404546
rect 705548 404534 705804 404540
rect 705548 404518 705792 404534
rect 705856 404530 705884 404654
rect 706316 404598 706344 404654
rect 706212 404592 706264 404598
rect 706008 404540 706212 404546
rect 706008 404534 706264 404540
rect 706304 404592 706356 404598
rect 706304 404534 706356 404540
rect 705844 404524 705896 404530
rect 706008 404518 706252 404534
rect 706454 404532 706482 404668
rect 706684 404666 706928 404682
rect 707092 404676 707388 404682
rect 707040 404670 707388 404676
rect 706672 404660 706928 404666
rect 706724 404654 706928 404660
rect 707052 404654 707388 404670
rect 707604 404654 707848 404682
rect 706672 404602 706724 404608
rect 706580 404592 706632 404598
rect 706632 404540 706928 404546
rect 706580 404534 706928 404540
rect 706592 404518 706928 404534
rect 707052 404530 707388 404546
rect 707604 404530 707632 404654
rect 707972 404546 708000 404738
rect 708524 404654 708768 404682
rect 707040 404524 707388 404530
rect 705844 404466 705896 404472
rect 707092 404518 707388 404524
rect 707592 404524 707644 404530
rect 707040 404466 707092 404472
rect 707972 404518 708308 404546
rect 707592 404466 707644 404472
rect 705384 404456 705436 404462
rect 705088 404394 705332 404410
rect 705384 404398 705436 404404
rect 707500 404456 707552 404462
rect 707552 404404 707848 404410
rect 707500 404398 707848 404404
rect 705088 404388 705344 404394
rect 705088 404382 705292 404388
rect 707512 404382 707848 404398
rect 708524 404394 708552 404654
rect 708892 404546 708920 404874
rect 708892 404518 709228 404546
rect 708512 404388 708564 404394
rect 705292 404330 705344 404336
rect 708512 404330 708564 404336
rect 704464 404320 704516 404326
rect 704168 404258 704412 404274
rect 704464 404262 704516 404268
rect 708420 404320 708472 404326
rect 708472 404268 708768 404274
rect 708420 404262 708768 404268
rect 704168 404252 704424 404258
rect 704168 404246 704372 404252
rect 708432 404246 708768 404262
rect 704372 404194 704424 404200
rect 676218 403744 676274 403753
rect 676218 403679 676274 403688
rect 676232 403306 676260 403679
rect 676220 403300 676272 403306
rect 676220 403242 676272 403248
rect 676126 402928 676182 402937
rect 676126 402863 676182 402872
rect 676126 402112 676182 402121
rect 676126 402047 676182 402056
rect 676140 401266 676168 402047
rect 676128 401260 676180 401266
rect 676128 401202 676180 401208
rect 676034 400208 676090 400217
rect 676034 400143 676090 400152
rect 676034 399800 676090 399809
rect 676034 399735 676090 399744
rect 676048 399498 676076 399735
rect 676036 399492 676088 399498
rect 676036 399434 676088 399440
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 675850 398576 675906 398585
rect 675850 398511 675906 398520
rect 675760 390584 675812 390590
rect 675760 390526 675812 390532
rect 675668 390516 675720 390522
rect 675668 390458 675720 390464
rect 675864 390402 675892 398511
rect 676048 398274 676076 399327
rect 676126 398848 676182 398857
rect 676126 398783 676182 398792
rect 676036 398268 676088 398274
rect 676036 398210 676088 398216
rect 676034 398168 676090 398177
rect 676034 398103 676090 398112
rect 675942 397760 675998 397769
rect 675942 397695 675998 397704
rect 675956 397662 675984 397695
rect 675944 397656 675996 397662
rect 675944 397598 675996 397604
rect 676048 397526 676076 398103
rect 676140 397594 676168 398783
rect 676128 397588 676180 397594
rect 676128 397530 676180 397536
rect 676036 397520 676088 397526
rect 676036 397462 676088 397468
rect 676034 397352 676090 397361
rect 676034 397287 676090 397296
rect 676048 396642 676076 397287
rect 676036 396636 676088 396642
rect 676036 396578 676088 396584
rect 676034 396536 676090 396545
rect 676034 396471 676090 396480
rect 675942 395720 675998 395729
rect 675942 395655 675998 395664
rect 675956 395418 675984 395655
rect 675944 395412 675996 395418
rect 675944 395354 675996 395360
rect 675942 395312 675998 395321
rect 675942 395247 675998 395256
rect 675956 394874 675984 395247
rect 676048 395010 676076 396471
rect 676126 395992 676182 396001
rect 676126 395927 676182 395936
rect 676036 395004 676088 395010
rect 676036 394946 676088 394952
rect 676034 394904 676090 394913
rect 675944 394868 675996 394874
rect 676034 394839 676090 394848
rect 675944 394810 675996 394816
rect 676048 394738 676076 394839
rect 676140 394806 676168 395927
rect 676128 394800 676180 394806
rect 676128 394742 676180 394748
rect 676036 394732 676088 394738
rect 676036 394674 676088 394680
rect 676034 394496 676090 394505
rect 676034 394431 676090 394440
rect 676048 394194 676076 394431
rect 676036 394188 676088 394194
rect 676036 394130 676088 394136
rect 676034 394088 676090 394097
rect 676034 394023 676090 394032
rect 676048 392018 676076 394023
rect 678978 393544 679034 393553
rect 678978 393479 679034 393488
rect 678992 393145 679020 393479
rect 678978 393136 679034 393145
rect 678978 393071 679034 393080
rect 684498 393136 684554 393145
rect 684498 393071 684554 393080
rect 678992 392086 679020 393071
rect 684512 392737 684540 393071
rect 684498 392728 684554 392737
rect 684498 392663 684554 392672
rect 678980 392080 679032 392086
rect 678980 392022 679032 392028
rect 676036 392012 676088 392018
rect 676036 391954 676088 391960
rect 675772 390374 675892 390402
rect 675772 386442 675800 390374
rect 675760 386436 675812 386442
rect 675760 386378 675812 386384
rect 675760 386164 675812 386170
rect 675760 386106 675812 386112
rect 675772 385696 675800 386106
rect 675312 385070 675418 385098
rect 675300 385008 675352 385014
rect 675300 384950 675352 384956
rect 675312 384449 675340 384950
rect 675312 384421 675418 384449
rect 675208 384124 675260 384130
rect 675208 384066 675260 384072
rect 675300 383920 675352 383926
rect 675300 383862 675352 383868
rect 675116 382492 675168 382498
rect 675116 382434 675168 382440
rect 675116 382356 675168 382362
rect 675116 382298 675168 382304
rect 675024 381948 675076 381954
rect 675024 381890 675076 381896
rect 675128 374134 675156 382298
rect 675312 380894 675340 383862
rect 675392 383172 675444 383178
rect 675392 383114 675444 383120
rect 675404 382568 675432 383114
rect 675392 382492 675444 382498
rect 675392 382434 675444 382440
rect 675404 382024 675432 382434
rect 675392 381948 675444 381954
rect 675392 381890 675444 381896
rect 675404 381412 675432 381890
rect 675312 380866 675432 380894
rect 675404 380732 675432 380866
rect 675300 379500 675352 379506
rect 675300 379442 675352 379448
rect 675312 378298 675340 379442
rect 675312 378270 675418 378298
rect 675300 378208 675352 378214
rect 675300 378150 675352 378156
rect 675312 377074 675340 378150
rect 675484 378004 675536 378010
rect 675484 377946 675536 377952
rect 675496 377740 675524 377946
rect 675312 377046 675418 377074
rect 675484 376984 675536 376990
rect 675484 376926 675536 376932
rect 675300 376916 675352 376922
rect 675300 376858 675352 376864
rect 675312 375238 675340 376858
rect 675496 376448 675524 376926
rect 675312 375210 675418 375238
rect 675116 374128 675168 374134
rect 675116 374070 675168 374076
rect 675300 374128 675352 374134
rect 675300 374070 675352 374076
rect 675312 372910 675340 374070
rect 675392 373924 675444 373930
rect 675392 373866 675444 373872
rect 675404 373388 675432 373866
rect 675300 372904 675352 372910
rect 675300 372846 675352 372852
rect 675300 372700 675352 372706
rect 675300 372642 675352 372648
rect 674748 370796 674800 370802
rect 674748 370738 674800 370744
rect 674668 361546 674788 361574
rect 674760 357513 674788 361546
rect 674746 357504 674802 357513
rect 674746 357439 674802 357448
rect 673276 357060 673328 357066
rect 673276 357002 673328 357008
rect 673288 356114 673316 357002
rect 673368 356176 673420 356182
rect 673368 356118 673420 356124
rect 673000 356108 673052 356114
rect 673000 356050 673052 356056
rect 673276 356108 673328 356114
rect 673276 356050 673328 356056
rect 673012 343641 673040 356050
rect 673184 355428 673236 355434
rect 673184 355370 673236 355376
rect 673092 353524 673144 353530
rect 673092 353466 673144 353472
rect 672998 343632 673054 343641
rect 672998 343567 673054 343576
rect 673000 342440 673052 342446
rect 673000 342382 673052 342388
rect 672906 143168 672962 143177
rect 672906 143103 672962 143112
rect 673012 138145 673040 342382
rect 673104 310078 673132 353466
rect 673196 353394 673224 355370
rect 673276 354612 673328 354618
rect 673276 354554 673328 354560
rect 673288 353530 673316 354554
rect 673276 353524 673328 353530
rect 673276 353466 673328 353472
rect 673184 353388 673236 353394
rect 673184 353330 673236 353336
rect 673196 353294 673224 353330
rect 673196 353266 673316 353294
rect 673182 343632 673238 343641
rect 673182 343567 673238 343576
rect 673196 312526 673224 343567
rect 673184 312520 673236 312526
rect 673184 312462 673236 312468
rect 673288 310894 673316 353266
rect 673380 311710 673408 356118
rect 675312 355065 675340 372642
rect 675392 372088 675444 372094
rect 675392 372030 675444 372036
rect 675404 371552 675432 372030
rect 675760 370796 675812 370802
rect 675760 370738 675812 370744
rect 675668 370728 675720 370734
rect 675668 370670 675720 370676
rect 675574 357096 675630 357105
rect 675574 357031 675576 357040
rect 675628 357031 675630 357040
rect 675576 357002 675628 357008
rect 675680 356697 675708 370670
rect 675666 356688 675722 356697
rect 675666 356623 675722 356632
rect 675772 355881 675800 370738
rect 703452 361752 703504 361758
rect 703452 361694 703504 361700
rect 709340 361752 709392 361758
rect 709340 361694 709392 361700
rect 703464 359258 703492 361694
rect 709352 359802 709380 361694
rect 709228 359774 709380 359802
rect 708512 359712 708564 359718
rect 704168 359650 704504 359666
rect 708564 359660 708768 359666
rect 708512 359654 708768 359660
rect 704168 359644 704516 359650
rect 704168 359638 704464 359644
rect 704464 359586 704516 359592
rect 708420 359644 708472 359650
rect 708524 359638 708768 359654
rect 708420 359586 708472 359592
rect 704372 359576 704424 359582
rect 703708 359502 703860 359530
rect 707500 359576 707552 359582
rect 704372 359518 704424 359524
rect 703464 359230 703708 359258
rect 703832 358902 703860 359502
rect 704384 359258 704412 359518
rect 704628 359502 704964 359530
rect 705088 359502 705424 359530
rect 705548 359502 705884 359530
rect 706008 359502 706344 359530
rect 704168 359230 704412 359258
rect 704936 359174 704964 359502
rect 705292 359440 705344 359446
rect 705292 359382 705344 359388
rect 705304 359258 705332 359382
rect 705088 359230 705332 359258
rect 705396 359242 705424 359502
rect 705752 359440 705804 359446
rect 705752 359382 705804 359388
rect 705764 359258 705792 359382
rect 705856 359378 705884 359502
rect 706212 359440 706264 359446
rect 706212 359382 706264 359388
rect 705844 359372 705896 359378
rect 705844 359314 705896 359320
rect 706224 359258 706252 359382
rect 706316 359310 706344 359502
rect 706454 359380 706482 359516
rect 706592 359502 706928 359530
rect 707052 359514 707388 359530
rect 707552 359524 707848 359530
rect 707500 359518 707848 359524
rect 707040 359508 707388 359514
rect 706592 359446 706620 359502
rect 707092 359502 707388 359508
rect 707512 359502 707848 359518
rect 708064 359502 708308 359530
rect 707040 359450 707092 359456
rect 706580 359440 706632 359446
rect 706580 359382 706632 359388
rect 707040 359372 707092 359378
rect 707040 359314 707092 359320
rect 705384 359236 705436 359242
rect 705548 359230 705792 359258
rect 706008 359230 706252 359258
rect 706304 359304 706356 359310
rect 706304 359246 706356 359252
rect 706580 359304 706632 359310
rect 707052 359258 707080 359314
rect 706632 359252 706928 359258
rect 706580 359246 706928 359252
rect 706592 359230 706928 359246
rect 707052 359230 707388 359258
rect 707512 359242 707848 359258
rect 708064 359242 708092 359502
rect 708432 359258 708460 359586
rect 707500 359236 707848 359242
rect 705384 359178 705436 359184
rect 707552 359230 707848 359236
rect 708052 359236 708104 359242
rect 707500 359178 707552 359184
rect 708432 359230 708768 359258
rect 708052 359178 708104 359184
rect 704924 359168 704976 359174
rect 704628 359106 704872 359122
rect 704924 359110 704976 359116
rect 707960 359168 708012 359174
rect 708012 359116 708308 359122
rect 707960 359110 708308 359116
rect 704628 359100 704884 359106
rect 704628 359094 704832 359100
rect 707972 359094 708308 359110
rect 704832 359042 704884 359048
rect 703820 358896 703872 358902
rect 703820 358838 703872 358844
rect 708880 358896 708932 358902
rect 708932 358844 709228 358850
rect 708880 358838 709228 358844
rect 708892 358822 709228 358838
rect 675850 358728 675906 358737
rect 675850 358663 675906 358672
rect 675864 356250 675892 358663
rect 675942 358320 675998 358329
rect 675942 358255 675998 358264
rect 675956 356386 675984 358255
rect 676034 357912 676090 357921
rect 676034 357847 676090 357856
rect 676048 356522 676076 357847
rect 676036 356516 676088 356522
rect 676036 356458 676088 356464
rect 675944 356380 675996 356386
rect 675944 356322 675996 356328
rect 676034 356280 676090 356289
rect 675852 356244 675904 356250
rect 676034 356215 676090 356224
rect 675852 356186 675904 356192
rect 676048 356182 676076 356215
rect 676036 356176 676088 356182
rect 676036 356118 676088 356124
rect 675758 355872 675814 355881
rect 675758 355807 675814 355816
rect 676034 355464 676090 355473
rect 676034 355399 676036 355408
rect 676088 355399 676090 355408
rect 676036 355370 676088 355376
rect 675298 355056 675354 355065
rect 675298 354991 675354 355000
rect 676034 354648 676090 354657
rect 676034 354583 676036 354592
rect 676088 354583 676090 354592
rect 676036 354554 676088 354560
rect 676034 354240 676090 354249
rect 676034 354175 676090 354184
rect 676048 353530 676076 354175
rect 673552 353524 673604 353530
rect 673552 353466 673604 353472
rect 676036 353524 676088 353530
rect 676036 353466 676088 353472
rect 673460 351076 673512 351082
rect 673460 351018 673512 351024
rect 673472 333606 673500 351018
rect 673564 339794 673592 353466
rect 676034 353424 676090 353433
rect 676034 353359 676090 353368
rect 676048 353326 676076 353359
rect 674012 353320 674064 353326
rect 674012 353262 674064 353268
rect 676036 353320 676088 353326
rect 676036 353262 676088 353268
rect 673736 349852 673788 349858
rect 673736 349794 673788 349800
rect 673552 339788 673604 339794
rect 673552 339730 673604 339736
rect 673460 333600 673512 333606
rect 673460 333542 673512 333548
rect 673748 332246 673776 349794
rect 673828 347948 673880 347954
rect 673828 347890 673880 347896
rect 673736 332240 673788 332246
rect 673736 332182 673788 332188
rect 673840 331634 673868 347890
rect 673920 347880 673972 347886
rect 673920 347822 673972 347828
rect 673932 332994 673960 347822
rect 674024 341018 674052 353262
rect 676034 353016 676090 353025
rect 676034 352951 676090 352960
rect 675942 352608 675998 352617
rect 675942 352543 675998 352552
rect 675298 351792 675354 351801
rect 675298 351727 675354 351736
rect 674564 351484 674616 351490
rect 674564 351426 674616 351432
rect 674012 341012 674064 341018
rect 674012 340954 674064 340960
rect 674576 337958 674604 351426
rect 674656 350668 674708 350674
rect 674656 350610 674708 350616
rect 674564 337952 674616 337958
rect 674564 337894 674616 337900
rect 674668 336598 674696 350610
rect 674748 350600 674800 350606
rect 674748 350542 674800 350548
rect 674760 337074 674788 350542
rect 674840 347812 674892 347818
rect 674840 347754 674892 347760
rect 674748 337068 674800 337074
rect 674748 337010 674800 337016
rect 674656 336592 674708 336598
rect 674656 336534 674708 336540
rect 674852 336122 674880 347754
rect 675312 339878 675340 351727
rect 675956 351082 675984 352543
rect 676048 351490 676076 352951
rect 676036 351484 676088 351490
rect 676036 351426 676088 351432
rect 676034 351384 676090 351393
rect 676034 351319 676090 351328
rect 675944 351076 675996 351082
rect 675944 351018 675996 351024
rect 675942 350976 675998 350985
rect 675942 350911 675998 350920
rect 675956 350674 675984 350911
rect 675944 350668 675996 350674
rect 675944 350610 675996 350616
rect 676048 350606 676076 351319
rect 676036 350600 676088 350606
rect 676036 350542 676088 350548
rect 676034 350160 676090 350169
rect 676034 350095 676090 350104
rect 676048 349858 676076 350095
rect 676036 349852 676088 349858
rect 676036 349794 676088 349800
rect 676034 349752 676090 349761
rect 676034 349687 676090 349696
rect 675942 349344 675998 349353
rect 675942 349279 675998 349288
rect 675850 348936 675906 348945
rect 675850 348871 675906 348880
rect 675758 348528 675814 348537
rect 675758 348463 675814 348472
rect 675666 348120 675722 348129
rect 675666 348055 675722 348064
rect 675680 347313 675708 348055
rect 675772 347721 675800 348463
rect 675864 347954 675892 348871
rect 675852 347948 675904 347954
rect 675852 347890 675904 347896
rect 675956 347886 675984 349279
rect 675944 347880 675996 347886
rect 675944 347822 675996 347828
rect 676048 347818 676076 349687
rect 676036 347812 676088 347818
rect 676036 347754 676088 347760
rect 675758 347712 675814 347721
rect 675758 347647 675814 347656
rect 675666 347304 675722 347313
rect 675666 347239 675722 347248
rect 675772 342446 675800 347647
rect 675760 342440 675812 342446
rect 675760 342382 675812 342388
rect 675484 341012 675536 341018
rect 675484 340954 675536 340960
rect 675496 340544 675524 340954
rect 675312 339850 675418 339878
rect 675484 339788 675536 339794
rect 675484 339730 675536 339736
rect 675496 339252 675524 339730
rect 675484 337952 675536 337958
rect 675484 337894 675536 337900
rect 675496 337416 675524 337894
rect 675392 337068 675444 337074
rect 675392 337010 675444 337016
rect 675404 336843 675432 337010
rect 675392 336592 675444 336598
rect 675392 336534 675444 336540
rect 675404 336192 675432 336534
rect 674840 336116 674892 336122
rect 674840 336058 674892 336064
rect 675484 336116 675536 336122
rect 675484 336058 675536 336064
rect 675496 335580 675524 336058
rect 675392 333600 675444 333606
rect 675392 333542 675444 333548
rect 675404 333064 675432 333542
rect 673920 332988 673972 332994
rect 673920 332930 673972 332936
rect 675392 332988 675444 332994
rect 675392 332930 675444 332936
rect 675404 332520 675432 332930
rect 675392 332240 675444 332246
rect 675392 332182 675444 332188
rect 675404 331875 675432 332182
rect 673828 331628 673880 331634
rect 673828 331570 673880 331576
rect 675392 331628 675444 331634
rect 675392 331570 675444 331576
rect 675404 331228 675432 331570
rect 675666 330576 675722 330585
rect 675666 330511 675722 330520
rect 675680 330035 675708 330511
rect 675758 328400 675814 328409
rect 675758 328335 675814 328344
rect 675772 328168 675800 328335
rect 675758 326904 675814 326913
rect 675758 326839 675814 326848
rect 675772 326332 675800 326839
rect 704004 314764 704056 314770
rect 704004 314706 704056 314712
rect 708880 314764 708932 314770
rect 708880 314706 708932 314712
rect 703556 314486 703708 314514
rect 703556 314022 703584 314486
rect 704016 314242 704044 314706
rect 708512 314696 708564 314702
rect 704168 314634 704504 314650
rect 708892 314650 708920 314706
rect 708564 314644 708768 314650
rect 708512 314638 708768 314644
rect 704168 314628 704516 314634
rect 704168 314622 704464 314628
rect 704464 314570 704516 314576
rect 708420 314628 708472 314634
rect 708524 314622 708768 314638
rect 708892 314622 709228 314650
rect 708420 314570 708472 314576
rect 704372 314560 704424 314566
rect 707500 314560 707552 314566
rect 704372 314502 704424 314508
rect 704384 314242 704412 314502
rect 704628 314486 704964 314514
rect 705088 314486 705424 314514
rect 705548 314486 705884 314514
rect 706008 314486 706344 314514
rect 703708 314214 704044 314242
rect 704168 314214 704412 314242
rect 704936 314158 704964 314486
rect 705292 314424 705344 314430
rect 705292 314366 705344 314372
rect 705304 314242 705332 314366
rect 705088 314214 705332 314242
rect 705396 314226 705424 314486
rect 705752 314424 705804 314430
rect 705752 314366 705804 314372
rect 705764 314242 705792 314366
rect 705856 314362 705884 314486
rect 706212 314424 706264 314430
rect 706212 314366 706264 314372
rect 705844 314356 705896 314362
rect 705844 314298 705896 314304
rect 706224 314242 706252 314366
rect 706316 314294 706344 314486
rect 706454 314364 706482 314500
rect 706592 314486 706928 314514
rect 707052 314498 707388 314514
rect 707552 314508 707848 314514
rect 707500 314502 707848 314508
rect 707040 314492 707388 314498
rect 706592 314430 706620 314486
rect 707092 314486 707388 314492
rect 707512 314486 707848 314502
rect 708064 314486 708308 314514
rect 707040 314434 707092 314440
rect 706580 314424 706632 314430
rect 706580 314366 706632 314372
rect 707040 314356 707092 314362
rect 707040 314298 707092 314304
rect 705384 314220 705436 314226
rect 705548 314214 705792 314242
rect 706008 314214 706252 314242
rect 706304 314288 706356 314294
rect 706304 314230 706356 314236
rect 706580 314288 706632 314294
rect 707052 314242 707080 314298
rect 706632 314236 706928 314242
rect 706580 314230 706928 314236
rect 706592 314214 706928 314230
rect 707052 314214 707388 314242
rect 707512 314226 707848 314242
rect 708064 314226 708092 314486
rect 708432 314242 708460 314570
rect 707500 314220 707848 314226
rect 705384 314162 705436 314168
rect 707552 314214 707848 314220
rect 708052 314220 708104 314226
rect 707500 314162 707552 314168
rect 708432 314214 708768 314242
rect 708052 314162 708104 314168
rect 704924 314152 704976 314158
rect 704628 314090 704872 314106
rect 704924 314094 704976 314100
rect 707960 314152 708012 314158
rect 708012 314100 708308 314106
rect 707960 314094 708308 314100
rect 704628 314084 704884 314090
rect 704628 314078 704832 314084
rect 707972 314078 708308 314094
rect 704832 314026 704884 314032
rect 703544 314016 703596 314022
rect 703544 313958 703596 313964
rect 708880 314016 708932 314022
rect 708932 313964 709228 313970
rect 708880 313958 709228 313964
rect 708892 313942 709228 313958
rect 676218 313576 676274 313585
rect 676218 313511 676274 313520
rect 676036 313336 676088 313342
rect 676034 313304 676036 313313
rect 676088 313304 676090 313313
rect 676034 313239 676090 313248
rect 676036 312928 676088 312934
rect 676034 312896 676036 312905
rect 676088 312896 676090 312905
rect 676034 312831 676090 312840
rect 676036 312520 676088 312526
rect 676034 312488 676036 312497
rect 676088 312488 676090 312497
rect 676034 312423 676090 312432
rect 676036 312112 676088 312118
rect 676034 312080 676036 312089
rect 676088 312080 676090 312089
rect 676232 312050 676260 313511
rect 676034 312015 676090 312024
rect 676220 312044 676272 312050
rect 676220 311986 676272 311992
rect 673368 311704 673420 311710
rect 676036 311704 676088 311710
rect 673368 311646 673420 311652
rect 676034 311672 676036 311681
rect 676088 311672 676090 311681
rect 676034 311607 676090 311616
rect 676034 311264 676090 311273
rect 676034 311199 676090 311208
rect 676048 311030 676076 311199
rect 674748 311024 674800 311030
rect 674748 310966 674800 310972
rect 676036 311024 676088 311030
rect 676036 310966 676088 310972
rect 673276 310888 673328 310894
rect 673276 310830 673328 310836
rect 673092 310072 673144 310078
rect 673092 310014 673144 310020
rect 673184 309664 673236 309670
rect 673184 309606 673236 309612
rect 673092 300892 673144 300898
rect 673092 300834 673144 300840
rect 672998 138136 673054 138145
rect 672998 138071 673054 138080
rect 673104 132977 673132 300834
rect 673196 264994 673224 309606
rect 674196 309188 674248 309194
rect 674196 309130 674248 309136
rect 673552 308100 673604 308106
rect 673552 308042 673604 308048
rect 673460 306536 673512 306542
rect 673460 306478 673512 306484
rect 673472 281926 673500 306478
rect 673564 283762 673592 308042
rect 673920 306468 673972 306474
rect 673920 306410 673972 306416
rect 673736 305108 673788 305114
rect 673736 305050 673788 305056
rect 673644 303816 673696 303822
rect 673644 303758 673696 303764
rect 673656 286618 673684 303758
rect 673644 286612 673696 286618
rect 673644 286554 673696 286560
rect 673748 285598 673776 305050
rect 673828 304292 673880 304298
rect 673828 304234 673880 304240
rect 673840 287230 673868 304234
rect 673932 288590 673960 306410
rect 674012 303748 674064 303754
rect 674012 303690 674064 303696
rect 673920 288584 673972 288590
rect 673920 288526 673972 288532
rect 674024 287978 674052 303690
rect 674208 294574 674236 309130
rect 674472 306876 674524 306882
rect 674472 306818 674524 306824
rect 674196 294568 674248 294574
rect 674196 294510 674248 294516
rect 674484 292942 674512 306818
rect 674656 304836 674708 304842
rect 674656 304778 674708 304784
rect 674564 303680 674616 303686
rect 674564 303622 674616 303628
rect 674472 292936 674524 292942
rect 674472 292878 674524 292884
rect 674576 291106 674604 303622
rect 674668 291582 674696 304778
rect 674656 291576 674708 291582
rect 674656 291518 674708 291524
rect 674564 291100 674616 291106
rect 674564 291042 674616 291048
rect 674012 287972 674064 287978
rect 674012 287914 674064 287920
rect 673828 287224 673880 287230
rect 673828 287166 673880 287172
rect 673736 285592 673788 285598
rect 673736 285534 673788 285540
rect 673552 283756 673604 283762
rect 673552 283698 673604 283704
rect 673460 281920 673512 281926
rect 673460 281862 673512 281868
rect 674760 267714 674788 310966
rect 676036 310888 676088 310894
rect 676034 310856 676036 310865
rect 676088 310856 676090 310865
rect 676034 310791 676090 310800
rect 676036 310480 676088 310486
rect 676034 310448 676036 310457
rect 676088 310448 676090 310457
rect 676034 310383 676090 310392
rect 676036 310072 676088 310078
rect 676034 310040 676036 310049
rect 676088 310040 676090 310049
rect 676034 309975 676090 309984
rect 676036 309664 676088 309670
rect 676034 309632 676036 309641
rect 676088 309632 676090 309641
rect 676034 309567 676090 309576
rect 676034 309224 676090 309233
rect 676034 309159 676036 309168
rect 676088 309159 676090 309168
rect 676036 309130 676088 309136
rect 676034 308816 676090 308825
rect 676034 308751 676090 308760
rect 675758 308408 675814 308417
rect 675758 308343 675814 308352
rect 675116 306264 675168 306270
rect 675116 306206 675168 306212
rect 675128 301050 675156 306206
rect 675128 301022 675248 301050
rect 675220 295118 675248 301022
rect 675772 296206 675800 308343
rect 676048 308106 676076 308751
rect 676036 308100 676088 308106
rect 676036 308042 676088 308048
rect 676034 308000 676090 308009
rect 676034 307935 676090 307944
rect 675942 307184 675998 307193
rect 675942 307119 675998 307128
rect 675956 306542 675984 307119
rect 676048 306882 676076 307935
rect 676126 307456 676182 307465
rect 676126 307391 676182 307400
rect 676036 306876 676088 306882
rect 676036 306818 676088 306824
rect 676034 306776 676090 306785
rect 676034 306711 676090 306720
rect 675944 306536 675996 306542
rect 675944 306478 675996 306484
rect 676048 306406 676076 306711
rect 676140 306474 676168 307391
rect 676128 306468 676180 306474
rect 676128 306410 676180 306416
rect 676036 306400 676088 306406
rect 676036 306342 676088 306348
rect 676034 305960 676090 305969
rect 676034 305895 676090 305904
rect 676048 304842 676076 305895
rect 676126 305416 676182 305425
rect 676126 305351 676182 305360
rect 676140 305114 676168 305351
rect 676128 305108 676180 305114
rect 676128 305050 676180 305056
rect 676126 305008 676182 305017
rect 676126 304943 676182 304952
rect 676036 304836 676088 304842
rect 676036 304778 676088 304784
rect 676034 304736 676090 304745
rect 676034 304671 676090 304680
rect 675942 303920 675998 303929
rect 675942 303855 675998 303864
rect 675956 303822 675984 303855
rect 675944 303816 675996 303822
rect 675944 303758 675996 303764
rect 676048 303686 676076 304671
rect 676140 304298 676168 304943
rect 676128 304292 676180 304298
rect 676128 304234 676180 304240
rect 676126 304192 676182 304201
rect 676126 304127 676182 304136
rect 676140 303754 676168 304127
rect 676128 303748 676180 303754
rect 676128 303690 676180 303696
rect 676036 303680 676088 303686
rect 676036 303622 676088 303628
rect 679070 303376 679126 303385
rect 679070 303311 679126 303320
rect 679084 302977 679112 303311
rect 679070 302968 679126 302977
rect 679070 302903 679126 302912
rect 684498 302968 684554 302977
rect 684498 302903 684554 302912
rect 679084 300898 679112 302903
rect 684512 302569 684540 302903
rect 684498 302560 684554 302569
rect 684498 302495 684554 302504
rect 679072 300892 679124 300898
rect 679072 300834 679124 300840
rect 675760 296200 675812 296206
rect 675760 296142 675812 296148
rect 675760 295996 675812 296002
rect 675760 295938 675812 295944
rect 675772 295528 675800 295938
rect 675208 295112 675260 295118
rect 675208 295054 675260 295060
rect 675392 295112 675444 295118
rect 675392 295054 675444 295060
rect 675404 294879 675432 295054
rect 675392 294568 675444 294574
rect 675392 294510 675444 294516
rect 675404 294236 675432 294510
rect 675392 292936 675444 292942
rect 675392 292878 675444 292884
rect 675404 292400 675432 292878
rect 675758 292224 675814 292233
rect 675758 292159 675814 292168
rect 675772 291856 675800 292159
rect 675392 291576 675444 291582
rect 675392 291518 675444 291524
rect 675404 291176 675432 291518
rect 675392 291100 675444 291106
rect 675392 291042 675444 291048
rect 675404 290564 675432 291042
rect 675392 288584 675444 288590
rect 675392 288526 675444 288532
rect 675404 288048 675432 288526
rect 675392 287972 675444 287978
rect 675392 287914 675444 287920
rect 675404 287504 675432 287914
rect 675484 287224 675536 287230
rect 675484 287166 675536 287172
rect 675496 286892 675524 287166
rect 675392 286612 675444 286618
rect 675392 286554 675444 286560
rect 675404 286212 675432 286554
rect 675484 285592 675536 285598
rect 675484 285534 675536 285540
rect 675496 285056 675524 285534
rect 675484 283756 675536 283762
rect 675484 283698 675536 283704
rect 675496 283220 675524 283698
rect 675392 281920 675444 281926
rect 675392 281862 675444 281868
rect 675404 281355 675432 281862
rect 703708 269754 704044 269770
rect 708984 269754 709228 269770
rect 703544 269748 703596 269754
rect 703708 269748 704056 269754
rect 703708 269742 704004 269748
rect 703544 269690 703596 269696
rect 704004 269690 704056 269696
rect 708880 269748 708932 269754
rect 708880 269690 708932 269696
rect 708972 269748 709228 269754
rect 709024 269742 709228 269748
rect 708972 269690 709024 269696
rect 703556 269362 703584 269690
rect 708052 269680 708104 269686
rect 704628 269618 704964 269634
rect 708104 269628 708308 269634
rect 708052 269622 708308 269628
rect 704628 269612 704976 269618
rect 704628 269606 704924 269612
rect 704924 269554 704976 269560
rect 707960 269612 708012 269618
rect 708064 269606 708308 269622
rect 707960 269554 708012 269560
rect 704832 269544 704884 269550
rect 704168 269470 704504 269498
rect 707040 269544 707092 269550
rect 704832 269486 704884 269492
rect 703556 269334 703708 269362
rect 704476 269142 704504 269470
rect 704844 269362 704872 269486
rect 705088 269470 705424 269498
rect 705548 269470 705884 269498
rect 706008 269470 706344 269498
rect 704628 269334 704872 269362
rect 705396 269278 705424 269470
rect 705752 269408 705804 269414
rect 705548 269356 705752 269362
rect 705548 269350 705804 269356
rect 705548 269334 705792 269350
rect 705856 269346 705884 269470
rect 706316 269414 706344 269470
rect 706212 269408 706264 269414
rect 706008 269356 706212 269362
rect 706008 269350 706264 269356
rect 706304 269408 706356 269414
rect 706304 269350 706356 269356
rect 705844 269340 705896 269346
rect 706008 269334 706252 269350
rect 706454 269348 706482 269484
rect 706684 269482 706928 269498
rect 707092 269492 707388 269498
rect 707040 269486 707388 269492
rect 706672 269476 706928 269482
rect 706724 269470 706928 269476
rect 707052 269470 707388 269486
rect 707604 269470 707848 269498
rect 706672 269418 706724 269424
rect 706580 269408 706632 269414
rect 706632 269356 706928 269362
rect 706580 269350 706928 269356
rect 706592 269334 706928 269350
rect 707052 269346 707388 269362
rect 707604 269346 707632 269470
rect 707972 269362 708000 269554
rect 708524 269470 708768 269498
rect 707040 269340 707388 269346
rect 705844 269282 705896 269288
rect 707092 269334 707388 269340
rect 707592 269340 707644 269346
rect 707040 269282 707092 269288
rect 707972 269334 708308 269362
rect 707592 269282 707644 269288
rect 705384 269272 705436 269278
rect 705088 269210 705332 269226
rect 705384 269214 705436 269220
rect 707500 269272 707552 269278
rect 707552 269220 707848 269226
rect 707500 269214 707848 269220
rect 705088 269204 705344 269210
rect 705088 269198 705292 269204
rect 707512 269198 707848 269214
rect 708524 269210 708552 269470
rect 708892 269362 708920 269690
rect 708892 269334 709228 269362
rect 708512 269204 708564 269210
rect 705292 269146 705344 269152
rect 708512 269146 708564 269152
rect 704464 269136 704516 269142
rect 704168 269074 704412 269090
rect 704464 269078 704516 269084
rect 708420 269136 708472 269142
rect 708472 269084 708768 269090
rect 708420 269078 708768 269084
rect 704168 269068 704424 269074
rect 704168 269062 704372 269068
rect 708432 269062 708768 269078
rect 704372 269010 704424 269016
rect 676126 268560 676182 268569
rect 676126 268495 676182 268504
rect 676036 267980 676088 267986
rect 676036 267922 676088 267928
rect 676048 267889 676076 267922
rect 676034 267880 676090 267889
rect 676034 267815 676090 267824
rect 676140 267782 676168 268495
rect 676218 268152 676274 268161
rect 676218 268087 676220 268096
rect 676272 268087 676274 268096
rect 676220 268058 676272 268064
rect 676128 267776 676180 267782
rect 676128 267718 676180 267724
rect 674748 267708 674800 267714
rect 674748 267650 674800 267656
rect 676036 267708 676088 267714
rect 676036 267650 676088 267656
rect 675944 267504 675996 267510
rect 675942 267472 675944 267481
rect 675996 267472 675998 267481
rect 675942 267407 675998 267416
rect 675758 267064 675814 267073
rect 675758 266999 675814 267008
rect 675668 266348 675720 266354
rect 675668 266290 675720 266296
rect 675680 265441 675708 266290
rect 675666 265432 675722 265441
rect 674748 265396 674800 265402
rect 675666 265367 675722 265376
rect 674748 265338 674800 265344
rect 673184 264988 673236 264994
rect 674760 264974 674788 265338
rect 673184 264930 673236 264936
rect 674576 264946 674788 264974
rect 674196 263084 674248 263090
rect 674196 263026 674248 263032
rect 673736 262404 673788 262410
rect 673736 262346 673788 262352
rect 673460 260228 673512 260234
rect 673460 260170 673512 260176
rect 673472 240582 673500 260170
rect 673552 259752 673604 259758
rect 673552 259694 673604 259700
rect 673564 242214 673592 259694
rect 673644 256828 673696 256834
rect 673644 256770 673696 256776
rect 673552 242208 673604 242214
rect 673552 242150 673604 242156
rect 673656 241602 673684 256770
rect 673748 243642 673776 262346
rect 674012 262336 674064 262342
rect 674012 262278 674064 262284
rect 673828 256760 673880 256766
rect 673828 256702 673880 256708
rect 673736 243636 673788 243642
rect 673736 243578 673788 243584
rect 673840 242962 673868 256702
rect 674024 247178 674052 262278
rect 674104 261860 674156 261866
rect 674104 261802 674156 261808
rect 674012 247172 674064 247178
rect 674012 247114 674064 247120
rect 674116 245654 674144 261802
rect 674208 249626 674236 263026
rect 674288 262268 674340 262274
rect 674288 262210 674340 262216
rect 674196 249620 674248 249626
rect 674196 249562 674248 249568
rect 674300 247926 674328 262210
rect 674472 259684 674524 259690
rect 674472 259626 674524 259632
rect 674380 259616 674432 259622
rect 674380 259558 674432 259564
rect 674288 247920 674340 247926
rect 674288 247862 674340 247868
rect 674392 246566 674420 259558
rect 674484 247314 674512 259626
rect 674472 247308 674524 247314
rect 674472 247250 674524 247256
rect 674472 247172 674524 247178
rect 674472 247114 674524 247120
rect 674380 246560 674432 246566
rect 674380 246502 674432 246508
rect 674116 245626 674420 245654
rect 673828 242956 673880 242962
rect 673828 242898 673880 242904
rect 673644 241596 673696 241602
rect 673644 241538 673696 241544
rect 673460 240576 673512 240582
rect 673460 240518 673512 240524
rect 674392 236910 674420 245626
rect 674484 241942 674512 247114
rect 674472 241936 674524 241942
rect 674472 241878 674524 241884
rect 674380 236904 674432 236910
rect 674380 236846 674432 236852
rect 674576 222222 674604 264946
rect 675574 260536 675630 260545
rect 675574 260471 675630 260480
rect 675588 260234 675616 260471
rect 675576 260228 675628 260234
rect 675576 260170 675628 260176
rect 675574 260128 675630 260137
rect 675574 260063 675630 260072
rect 675588 259758 675616 260063
rect 675576 259752 675628 259758
rect 675576 259694 675628 259700
rect 675024 259548 675076 259554
rect 675024 259490 675076 259496
rect 674748 255332 674800 255338
rect 674748 255274 674800 255280
rect 674656 255264 674708 255270
rect 674656 255206 674708 255212
rect 674668 235550 674696 255206
rect 674760 235618 674788 255274
rect 675036 247602 675064 259490
rect 675208 259480 675260 259486
rect 675208 259422 675260 259428
rect 675220 250442 675248 259422
rect 675680 255338 675708 265367
rect 675772 265062 675800 266999
rect 676048 266665 676076 267650
rect 676034 266656 676090 266665
rect 676034 266591 676090 266600
rect 676034 266248 676090 266257
rect 676034 266183 676090 266192
rect 676048 265402 676076 266183
rect 676220 266144 676272 266150
rect 676218 266112 676220 266121
rect 676272 266112 676274 266121
rect 676218 266047 676274 266056
rect 676036 265396 676088 265402
rect 676036 265338 676088 265344
rect 675760 265056 675812 265062
rect 675760 264998 675812 265004
rect 675668 255332 675720 255338
rect 675668 255274 675720 255280
rect 675772 255270 675800 264998
rect 676220 264988 676272 264994
rect 676220 264930 676272 264936
rect 676232 264897 676260 264930
rect 676218 264888 676274 264897
rect 676218 264823 676274 264832
rect 676034 264208 676090 264217
rect 676034 264143 676090 264152
rect 675850 263392 675906 263401
rect 675850 263327 675906 263336
rect 675760 255264 675812 255270
rect 675760 255206 675812 255212
rect 675864 255082 675892 263327
rect 676048 263090 676076 264143
rect 676126 263664 676182 263673
rect 676126 263599 676182 263608
rect 676036 263084 676088 263090
rect 676036 263026 676088 263032
rect 676034 262984 676090 262993
rect 676034 262919 676090 262928
rect 675942 262576 675998 262585
rect 675942 262511 675998 262520
rect 675956 262410 675984 262511
rect 675944 262404 675996 262410
rect 675944 262346 675996 262352
rect 676048 262274 676076 262919
rect 676140 262342 676168 263599
rect 676128 262336 676180 262342
rect 676128 262278 676180 262284
rect 676036 262268 676088 262274
rect 676036 262210 676088 262216
rect 676034 262168 676090 262177
rect 676034 262103 676090 262112
rect 676048 261866 676076 262103
rect 676036 261860 676088 261866
rect 676036 261802 676088 261808
rect 676034 261760 676090 261769
rect 676034 261695 676090 261704
rect 675942 260944 675998 260953
rect 675942 260879 675998 260888
rect 675956 259622 675984 260879
rect 675944 259616 675996 259622
rect 675944 259558 675996 259564
rect 676048 259486 676076 261695
rect 676126 261216 676182 261225
rect 676126 261151 676182 261160
rect 676140 259690 676168 261151
rect 676128 259684 676180 259690
rect 676128 259626 676180 259632
rect 676126 259584 676182 259593
rect 676126 259519 676128 259528
rect 676180 259519 676182 259528
rect 676128 259490 676180 259496
rect 676036 259480 676088 259486
rect 676036 259422 676088 259428
rect 676034 259312 676090 259321
rect 676034 259247 676090 259256
rect 676048 256766 676076 259247
rect 676126 258768 676182 258777
rect 676126 258703 676182 258712
rect 676140 256834 676168 258703
rect 678978 258360 679034 258369
rect 678978 258295 679034 258304
rect 678992 257961 679020 258295
rect 678978 257952 679034 257961
rect 678978 257887 679034 257896
rect 684498 257952 684554 257961
rect 684498 257887 684554 257896
rect 678992 256902 679020 257887
rect 684512 257553 684540 257887
rect 684498 257544 684554 257553
rect 684498 257479 684554 257488
rect 678980 256896 679032 256902
rect 678980 256838 679032 256844
rect 676128 256828 676180 256834
rect 676128 256770 676180 256776
rect 676036 256760 676088 256766
rect 676036 256702 676088 256708
rect 675772 255054 675892 255082
rect 675772 251258 675800 255054
rect 675760 251252 675812 251258
rect 675760 251194 675812 251200
rect 675760 250980 675812 250986
rect 675760 250922 675812 250928
rect 675772 250512 675800 250922
rect 675208 250436 675260 250442
rect 675208 250378 675260 250384
rect 675484 250436 675536 250442
rect 675484 250378 675536 250384
rect 675496 249900 675524 250378
rect 675392 249620 675444 249626
rect 675392 249562 675444 249568
rect 675404 249220 675432 249562
rect 675484 247920 675536 247926
rect 675484 247862 675536 247868
rect 675036 247574 675156 247602
rect 675128 246090 675156 247574
rect 675496 247384 675524 247862
rect 675392 247308 675444 247314
rect 675392 247250 675444 247256
rect 675404 246840 675432 247250
rect 675392 246560 675444 246566
rect 675392 246502 675444 246508
rect 675404 246199 675432 246502
rect 675116 246084 675168 246090
rect 675116 246026 675168 246032
rect 675392 246084 675444 246090
rect 675392 246026 675444 246032
rect 675404 245548 675432 246026
rect 675300 243636 675352 243642
rect 675300 243578 675352 243584
rect 675312 243085 675340 243578
rect 675312 243057 675418 243085
rect 675300 242956 675352 242962
rect 675300 242898 675352 242904
rect 675312 242533 675340 242898
rect 675312 242505 675418 242533
rect 675392 242208 675444 242214
rect 675392 242150 675444 242156
rect 675300 241936 675352 241942
rect 675300 241878 675352 241884
rect 675312 238218 675340 241878
rect 675404 241876 675432 242150
rect 675392 241596 675444 241602
rect 675392 241538 675444 241544
rect 675404 241231 675432 241538
rect 675392 240576 675444 240582
rect 675392 240518 675444 240524
rect 675404 240040 675432 240518
rect 675312 238190 675418 238218
rect 675392 236904 675444 236910
rect 675392 236846 675444 236852
rect 675404 236368 675432 236846
rect 674748 235612 674800 235618
rect 674748 235554 674800 235560
rect 675668 235612 675720 235618
rect 675668 235554 675720 235560
rect 674656 235544 674708 235550
rect 674656 235486 674708 235492
rect 674564 222216 674616 222222
rect 674564 222158 674616 222164
rect 674656 222148 674708 222154
rect 674656 222090 674708 222096
rect 675576 222148 675628 222154
rect 675576 222090 675628 222096
rect 673920 218340 673972 218346
rect 673920 218282 673972 218288
rect 673460 218136 673512 218142
rect 673460 218078 673512 218084
rect 673184 212492 673236 212498
rect 673184 212434 673236 212440
rect 673090 132968 673146 132977
rect 673090 132903 673146 132912
rect 672814 127936 672870 127945
rect 672814 127871 672870 127880
rect 673196 122913 673224 212434
rect 673472 193526 673500 218078
rect 673828 216300 673880 216306
rect 673828 216242 673880 216248
rect 673552 215892 673604 215898
rect 673552 215834 673604 215840
rect 673564 202450 673592 215834
rect 673644 214668 673696 214674
rect 673644 214610 673696 214616
rect 673656 202638 673684 214610
rect 673736 213852 673788 213858
rect 673736 213794 673788 213800
rect 673644 202632 673696 202638
rect 673644 202574 673696 202580
rect 673564 202422 673684 202450
rect 673552 202360 673604 202366
rect 673552 202302 673604 202308
rect 673460 193520 673512 193526
rect 673460 193462 673512 193468
rect 673564 191690 673592 202302
rect 673656 198422 673684 202422
rect 673644 198416 673696 198422
rect 673644 198358 673696 198364
rect 673748 197606 673776 213794
rect 673840 202774 673868 216242
rect 673932 205222 673960 218282
rect 674380 218068 674432 218074
rect 674380 218010 674432 218016
rect 674012 216708 674064 216714
rect 674012 216650 674064 216656
rect 673920 205216 673972 205222
rect 673920 205158 673972 205164
rect 673828 202768 673880 202774
rect 673828 202710 673880 202716
rect 673828 202632 673880 202638
rect 673828 202574 673880 202580
rect 673736 197600 673788 197606
rect 673736 197542 673788 197548
rect 673840 197062 673868 202574
rect 674024 198734 674052 216650
rect 674104 215484 674156 215490
rect 674104 215426 674156 215432
rect 674116 201958 674144 215426
rect 674196 215416 674248 215422
rect 674196 215358 674248 215364
rect 674104 201952 674156 201958
rect 674104 201894 674156 201900
rect 674208 201550 674236 215358
rect 674288 208412 674340 208418
rect 674288 208354 674340 208360
rect 674196 201544 674248 201550
rect 674196 201486 674248 201492
rect 674300 200818 674328 208354
rect 674392 205562 674420 218010
rect 674668 212906 674696 222090
rect 675588 221921 675616 222090
rect 675574 221912 675630 221921
rect 675574 221847 675630 221856
rect 675680 220697 675708 235554
rect 675760 235544 675812 235550
rect 675760 235486 675812 235492
rect 675772 222329 675800 235486
rect 704004 224528 704056 224534
rect 703717 224476 704004 224482
rect 708880 224528 708932 224534
rect 703717 224470 704056 224476
rect 703717 224454 704044 224470
rect 704177 224466 704504 224482
rect 708880 224470 708932 224476
rect 704177 224460 704516 224466
rect 704177 224454 704464 224460
rect 704464 224402 704516 224408
rect 708420 224460 708472 224466
rect 708420 224402 708472 224408
rect 707500 224392 707552 224398
rect 704002 224360 704058 224369
rect 704637 224318 704964 224346
rect 705097 224318 705424 224346
rect 705557 224318 705884 224346
rect 706017 224318 706344 224346
rect 704002 224295 704058 224304
rect 704016 224074 704044 224295
rect 704462 224224 704518 224233
rect 704462 224159 704518 224168
rect 704476 224074 704504 224159
rect 703708 224046 704044 224074
rect 704168 224046 704504 224074
rect 704936 223990 704964 224318
rect 705292 224256 705344 224262
rect 705292 224198 705344 224204
rect 705304 224074 705332 224198
rect 705088 224046 705332 224074
rect 705396 224058 705424 224318
rect 705752 224256 705804 224262
rect 705752 224198 705804 224204
rect 705764 224074 705792 224198
rect 705856 224194 705884 224318
rect 706212 224256 706264 224262
rect 706212 224198 706264 224204
rect 705844 224188 705896 224194
rect 705844 224130 705896 224136
rect 706224 224074 706252 224198
rect 706316 224126 706344 224318
rect 706454 224196 706482 224332
rect 706592 224318 706928 224346
rect 707052 224330 707388 224346
rect 707552 224340 707848 224346
rect 707500 224334 707848 224340
rect 707040 224324 707388 224330
rect 706592 224262 706620 224318
rect 707092 224318 707388 224324
rect 707512 224318 707848 224334
rect 708064 224318 708308 224346
rect 707040 224266 707092 224272
rect 706580 224256 706632 224262
rect 706580 224198 706632 224204
rect 707040 224188 707092 224194
rect 707040 224130 707092 224136
rect 705384 224052 705436 224058
rect 705548 224046 705792 224074
rect 706008 224046 706252 224074
rect 706304 224120 706356 224126
rect 706304 224062 706356 224068
rect 706580 224120 706632 224126
rect 707052 224074 707080 224130
rect 706632 224068 706928 224074
rect 706580 224062 706928 224068
rect 706592 224046 706928 224062
rect 707052 224046 707388 224074
rect 707512 224058 707848 224074
rect 708064 224058 708092 224318
rect 708432 224074 708460 224402
rect 708524 224318 708768 224346
rect 708524 224233 708552 224318
rect 708510 224224 708566 224233
rect 708510 224159 708566 224168
rect 708892 224074 708920 224470
rect 708970 224360 709026 224369
rect 709026 224318 709228 224346
rect 708970 224295 709026 224304
rect 707500 224052 707848 224058
rect 705384 223994 705436 224000
rect 707552 224046 707848 224052
rect 708052 224052 708104 224058
rect 707500 223994 707552 224000
rect 708432 224046 708768 224074
rect 708892 224046 709228 224074
rect 708052 223994 708104 224000
rect 704924 223984 704976 223990
rect 704628 223922 704872 223938
rect 704924 223926 704976 223932
rect 707960 223984 708012 223990
rect 708012 223932 708308 223938
rect 707960 223926 708308 223932
rect 704628 223916 704884 223922
rect 704628 223910 704832 223916
rect 707972 223910 708308 223926
rect 704832 223858 704884 223864
rect 676034 223544 676090 223553
rect 676034 223479 676090 223488
rect 675850 223136 675906 223145
rect 675850 223071 675906 223080
rect 675758 222320 675814 222329
rect 675758 222255 675814 222264
rect 675760 222216 675812 222222
rect 675760 222158 675812 222164
rect 675772 221513 675800 222158
rect 675758 221504 675814 221513
rect 675758 221439 675814 221448
rect 675758 221096 675814 221105
rect 675864 221066 675892 223071
rect 675942 222728 675998 222737
rect 675942 222663 675998 222672
rect 675758 221031 675814 221040
rect 675852 221060 675904 221066
rect 675666 220688 675722 220697
rect 675666 220623 675722 220632
rect 675576 220176 675628 220182
rect 675576 220118 675628 220124
rect 674840 220108 674892 220114
rect 674840 220050 674892 220056
rect 674852 218054 674880 220050
rect 674760 218026 674880 218054
rect 674656 212900 674708 212906
rect 674656 212842 674708 212848
rect 674760 212786 674788 218026
rect 675208 215348 675260 215354
rect 675208 215290 675260 215296
rect 674576 212758 674788 212786
rect 674472 212560 674524 212566
rect 674472 212502 674524 212508
rect 674380 205556 674432 205562
rect 674380 205498 674432 205504
rect 674380 205420 674432 205426
rect 674380 205362 674432 205368
rect 674392 202366 674420 205362
rect 674380 202360 674432 202366
rect 674380 202302 674432 202308
rect 674484 200938 674512 212502
rect 674472 200932 674524 200938
rect 674472 200874 674524 200880
rect 674300 200790 674512 200818
rect 674024 198706 674420 198734
rect 673828 197056 673880 197062
rect 673828 196998 673880 197004
rect 674392 195226 674420 198706
rect 674484 196450 674512 200790
rect 674472 196444 674524 196450
rect 674472 196386 674524 196392
rect 674380 195220 674432 195226
rect 674380 195162 674432 195168
rect 673552 191684 673604 191690
rect 673552 191626 673604 191632
rect 673276 176928 673328 176934
rect 673276 176870 673328 176876
rect 673288 132326 673316 176870
rect 674576 176390 674604 212758
rect 674748 212696 674800 212702
rect 674748 212638 674800 212644
rect 674656 212628 674708 212634
rect 674656 212570 674708 212576
rect 674668 196586 674696 212570
rect 674656 196580 674708 196586
rect 674656 196522 674708 196528
rect 674656 196444 674708 196450
rect 674656 196386 674708 196392
rect 674564 176384 674616 176390
rect 674564 176326 674616 176332
rect 673368 176044 673420 176050
rect 673368 175986 673420 175992
rect 673276 132320 673328 132326
rect 673276 132262 673328 132268
rect 673380 131510 673408 175986
rect 674668 175574 674696 196386
rect 674760 179382 674788 212638
rect 675220 208350 675248 215290
rect 675390 212528 675446 212537
rect 675390 212463 675392 212472
rect 675444 212463 675446 212472
rect 675392 212434 675444 212440
rect 675588 208418 675616 220118
rect 675666 217016 675722 217025
rect 675666 216951 675722 216960
rect 675576 208412 675628 208418
rect 675576 208354 675628 208360
rect 674840 208344 674892 208350
rect 674840 208286 674892 208292
rect 675208 208344 675260 208350
rect 675208 208286 675260 208292
rect 674852 202094 674880 208286
rect 675680 206038 675708 216951
rect 675772 216714 675800 221031
rect 675852 221002 675904 221008
rect 675956 220998 675984 222663
rect 676048 221202 676076 223479
rect 676036 221196 676088 221202
rect 676036 221138 676088 221144
rect 675944 220992 675996 220998
rect 675944 220934 675996 220940
rect 675942 220280 675998 220289
rect 675942 220215 675998 220224
rect 675956 220114 675984 220215
rect 676036 220176 676088 220182
rect 676036 220118 676088 220124
rect 675944 220108 675996 220114
rect 675944 220050 675996 220056
rect 676048 219473 676076 220118
rect 676034 219464 676090 219473
rect 676034 219399 676090 219408
rect 676034 219056 676090 219065
rect 676034 218991 676090 219000
rect 675942 218648 675998 218657
rect 675942 218583 675998 218592
rect 675956 218142 675984 218583
rect 676048 218346 676076 218991
rect 676036 218340 676088 218346
rect 676036 218282 676088 218288
rect 676034 218240 676090 218249
rect 676034 218175 676090 218184
rect 675944 218136 675996 218142
rect 675944 218078 675996 218084
rect 676048 218074 676076 218175
rect 676036 218068 676088 218074
rect 676036 218010 676088 218016
rect 676034 217832 676090 217841
rect 676034 217767 676090 217776
rect 675942 217424 675998 217433
rect 675942 217359 675998 217368
rect 675760 216708 675812 216714
rect 675760 216650 675812 216656
rect 675758 216608 675814 216617
rect 675758 216543 675814 216552
rect 675772 206038 675800 216543
rect 675956 215898 675984 217359
rect 676048 216306 676076 217767
rect 676036 216300 676088 216306
rect 676036 216242 676088 216248
rect 676034 216200 676090 216209
rect 676034 216135 676090 216144
rect 675944 215892 675996 215898
rect 675944 215834 675996 215840
rect 675942 215792 675998 215801
rect 675942 215727 675998 215736
rect 675852 215484 675904 215490
rect 675852 215426 675904 215432
rect 675864 215393 675892 215426
rect 675956 215422 675984 215727
rect 675944 215416 675996 215422
rect 675850 215384 675906 215393
rect 675944 215358 675996 215364
rect 676048 215354 676076 216135
rect 675850 215319 675906 215328
rect 676036 215348 676088 215354
rect 676036 215290 676088 215296
rect 676034 214976 676090 214985
rect 676034 214911 676090 214920
rect 676048 214674 676076 214911
rect 676036 214668 676088 214674
rect 676036 214610 676088 214616
rect 676034 214568 676090 214577
rect 676034 214503 676090 214512
rect 675942 214160 675998 214169
rect 675942 214095 675998 214104
rect 675956 213858 675984 214095
rect 675944 213852 675996 213858
rect 675944 213794 675996 213800
rect 675942 213752 675998 213761
rect 675942 213687 675998 213696
rect 675850 212936 675906 212945
rect 675850 212871 675906 212880
rect 675864 212129 675892 212871
rect 675956 212634 675984 213687
rect 675944 212628 675996 212634
rect 675944 212570 675996 212576
rect 676048 212566 676076 214503
rect 676036 212560 676088 212566
rect 676036 212502 676088 212508
rect 675850 212120 675906 212129
rect 675850 212055 675906 212064
rect 675668 206032 675720 206038
rect 675668 205974 675720 205980
rect 675760 206032 675812 206038
rect 675760 205974 675812 205980
rect 675300 205556 675352 205562
rect 675300 205498 675352 205504
rect 675312 205337 675340 205498
rect 675312 205309 675418 205337
rect 675300 205216 675352 205222
rect 675300 205158 675352 205164
rect 675312 204049 675340 205158
rect 675760 205012 675812 205018
rect 675760 204954 675812 204960
rect 675772 204680 675800 204954
rect 675312 204021 675418 204049
rect 675484 202768 675536 202774
rect 675484 202710 675536 202716
rect 675496 202195 675524 202710
rect 674840 202088 674892 202094
rect 674840 202030 674892 202036
rect 675392 202088 675444 202094
rect 675392 202030 675444 202036
rect 674840 201952 674892 201958
rect 674840 201894 674892 201900
rect 674852 195362 674880 201894
rect 675404 201620 675432 202030
rect 675392 201544 675444 201550
rect 675392 201486 675444 201492
rect 675404 201008 675432 201486
rect 675392 200932 675444 200938
rect 675392 200874 675444 200880
rect 675404 200328 675432 200874
rect 675392 198416 675444 198422
rect 675392 198358 675444 198364
rect 675404 197880 675432 198358
rect 675484 197600 675536 197606
rect 675484 197542 675536 197548
rect 675496 197336 675524 197542
rect 675392 197056 675444 197062
rect 675392 196998 675444 197004
rect 675404 196656 675432 196998
rect 675392 196580 675444 196586
rect 675392 196522 675444 196528
rect 675404 196044 675432 196522
rect 674840 195356 674892 195362
rect 674840 195298 674892 195304
rect 675392 195356 675444 195362
rect 675392 195298 675444 195304
rect 674840 195220 674892 195226
rect 674840 195162 674892 195168
rect 674748 179376 674800 179382
rect 674748 179318 674800 179324
rect 674852 176662 674880 195162
rect 675404 194820 675432 195298
rect 675392 193520 675444 193526
rect 675392 193462 675444 193468
rect 675404 192984 675432 193462
rect 675392 191684 675444 191690
rect 675392 191626 675444 191632
rect 675404 191148 675432 191626
rect 708512 179512 708564 179518
rect 704168 179450 704504 179466
rect 708564 179460 708768 179466
rect 708512 179454 708768 179460
rect 704168 179444 704516 179450
rect 704168 179438 704464 179444
rect 704464 179386 704516 179392
rect 708420 179444 708472 179450
rect 708524 179438 708768 179454
rect 708892 179438 709228 179466
rect 708420 179386 708472 179392
rect 675852 179376 675904 179382
rect 704372 179376 704424 179382
rect 703910 179344 703966 179353
rect 675852 179318 675904 179324
rect 675758 178528 675814 178537
rect 675758 178463 675814 178472
rect 675772 176866 675800 178463
rect 675864 177313 675892 179318
rect 703708 179302 703910 179330
rect 707500 179376 707552 179382
rect 704372 179318 704424 179324
rect 703910 179279 703966 179288
rect 704384 179058 704412 179318
rect 704628 179302 704964 179330
rect 705088 179302 705424 179330
rect 705548 179302 705884 179330
rect 706008 179302 706344 179330
rect 704168 179030 704412 179058
rect 704936 178974 704964 179302
rect 705292 179240 705344 179246
rect 705292 179182 705344 179188
rect 705304 179058 705332 179182
rect 705088 179030 705332 179058
rect 705396 179042 705424 179302
rect 705752 179240 705804 179246
rect 705752 179182 705804 179188
rect 705764 179058 705792 179182
rect 705856 179110 705884 179302
rect 706212 179240 706264 179246
rect 706212 179182 706264 179188
rect 705384 179036 705436 179042
rect 705548 179030 705792 179058
rect 705844 179104 705896 179110
rect 706224 179058 706252 179182
rect 706316 179178 706344 179302
rect 706454 179180 706482 179316
rect 706684 179302 706928 179330
rect 707052 179314 707388 179330
rect 707552 179324 707848 179330
rect 707500 179318 707848 179324
rect 707040 179308 707388 179314
rect 706684 179246 706712 179302
rect 707092 179302 707388 179308
rect 707512 179302 707848 179318
rect 708064 179302 708308 179330
rect 707040 179250 707092 179256
rect 706672 179240 706724 179246
rect 706672 179182 706724 179188
rect 706304 179172 706356 179178
rect 706304 179114 706356 179120
rect 706580 179172 706632 179178
rect 706580 179114 706632 179120
rect 705844 179046 705896 179052
rect 706008 179030 706252 179058
rect 706592 179058 706620 179114
rect 707040 179104 707092 179110
rect 706592 179030 706928 179058
rect 707092 179052 707388 179058
rect 707040 179046 707388 179052
rect 707052 179030 707388 179046
rect 707512 179042 707848 179058
rect 708064 179042 708092 179302
rect 708432 179058 708460 179386
rect 707500 179036 707848 179042
rect 705384 178978 705436 178984
rect 707552 179030 707848 179036
rect 708052 179036 708104 179042
rect 707500 178978 707552 178984
rect 708432 179030 708768 179058
rect 708052 178978 708104 178984
rect 704924 178968 704976 178974
rect 704628 178906 704872 178922
rect 704924 178910 704976 178916
rect 707960 178968 708012 178974
rect 708012 178916 708308 178922
rect 707960 178910 708308 178916
rect 704628 178900 704884 178906
rect 704628 178894 704832 178900
rect 707972 178894 708308 178910
rect 704832 178842 704884 178848
rect 708892 178838 708920 179438
rect 709062 179344 709118 179353
rect 709062 179279 709118 179288
rect 709076 179058 709104 179279
rect 709076 179030 709228 179058
rect 704004 178832 704056 178838
rect 703708 178780 704004 178786
rect 703708 178774 704056 178780
rect 708880 178832 708932 178838
rect 708880 178774 708932 178780
rect 703708 178758 704044 178774
rect 675942 178120 675998 178129
rect 675942 178055 675998 178064
rect 675850 177304 675906 177313
rect 675850 177239 675906 177248
rect 675956 177138 675984 178055
rect 676034 177712 676090 177721
rect 676034 177647 676090 177656
rect 675944 177132 675996 177138
rect 675944 177074 675996 177080
rect 676048 177002 676076 177647
rect 676036 176996 676088 177002
rect 676036 176938 676088 176944
rect 675944 176928 675996 176934
rect 675942 176896 675944 176905
rect 675996 176896 675998 176905
rect 675760 176860 675812 176866
rect 675942 176831 675998 176840
rect 675760 176802 675812 176808
rect 674840 176656 674892 176662
rect 674840 176598 674892 176604
rect 676036 176656 676088 176662
rect 676036 176598 676088 176604
rect 676048 176497 676076 176598
rect 676034 176488 676090 176497
rect 676034 176423 676090 176432
rect 676036 176384 676088 176390
rect 676036 176326 676088 176332
rect 675942 176080 675998 176089
rect 675942 176015 675944 176024
rect 675996 176015 675998 176024
rect 675944 175986 675996 175992
rect 676048 175681 676076 176326
rect 676034 175672 676090 175681
rect 676034 175607 676090 175616
rect 674656 175568 674708 175574
rect 674656 175510 674708 175516
rect 676036 175568 676088 175574
rect 676036 175510 676088 175516
rect 675944 175296 675996 175302
rect 675942 175264 675944 175273
rect 675996 175264 675998 175273
rect 675942 175199 675998 175208
rect 676048 174865 676076 175510
rect 676034 174856 676090 174865
rect 676034 174791 676090 174800
rect 676036 174480 676088 174486
rect 676034 174448 676036 174457
rect 676088 174448 676090 174457
rect 676034 174383 676090 174392
rect 676034 174040 676090 174049
rect 676034 173975 676090 173984
rect 676048 173942 676076 173975
rect 674104 173936 674156 173942
rect 674104 173878 674156 173884
rect 676036 173936 676088 173942
rect 676036 173878 676088 173884
rect 673460 171352 673512 171358
rect 673460 171294 673512 171300
rect 673472 153406 673500 171294
rect 673552 170060 673604 170066
rect 673552 170002 673604 170008
rect 673460 153400 673512 153406
rect 673460 153342 673512 153348
rect 673564 150414 673592 170002
rect 673736 169244 673788 169250
rect 673736 169186 673788 169192
rect 673644 168564 673696 168570
rect 673644 168506 673696 168512
rect 673656 151434 673684 168506
rect 673748 152046 673776 169186
rect 674012 168768 674064 168774
rect 674012 168710 674064 168716
rect 674024 152794 674052 168710
rect 674116 159390 674144 173878
rect 675758 173224 675814 173233
rect 675758 173159 675814 173168
rect 674840 171692 674892 171698
rect 674840 171634 674892 171640
rect 674564 171216 674616 171222
rect 674564 171158 674616 171164
rect 674104 159384 674156 159390
rect 674104 159326 674156 159332
rect 674576 156942 674604 171158
rect 674656 169652 674708 169658
rect 674656 169594 674708 169600
rect 674564 156936 674616 156942
rect 674564 156878 674616 156884
rect 674668 156534 674696 169594
rect 674748 168700 674800 168706
rect 674748 168642 674800 168648
rect 674656 156528 674708 156534
rect 674656 156470 674708 156476
rect 674760 155922 674788 168642
rect 674852 157758 674880 171634
rect 675208 171012 675260 171018
rect 675208 170954 675260 170960
rect 675220 160070 675248 170954
rect 675772 161022 675800 173159
rect 676034 172816 676090 172825
rect 676034 172751 676090 172760
rect 675942 172408 675998 172417
rect 675942 172343 675998 172352
rect 675956 171358 675984 172343
rect 676048 171698 676076 172751
rect 676036 171692 676088 171698
rect 676036 171634 676088 171640
rect 676034 171592 676090 171601
rect 676034 171527 676090 171536
rect 675944 171352 675996 171358
rect 675944 171294 675996 171300
rect 675944 171216 675996 171222
rect 675942 171184 675944 171193
rect 675996 171184 675998 171193
rect 676048 171154 676076 171527
rect 675942 171119 675998 171128
rect 676036 171148 676088 171154
rect 676036 171090 676088 171096
rect 676034 170776 676090 170785
rect 676034 170711 676090 170720
rect 675942 170368 675998 170377
rect 675942 170303 675998 170312
rect 675956 170066 675984 170303
rect 675944 170060 675996 170066
rect 675944 170002 675996 170008
rect 675942 169960 675998 169969
rect 675942 169895 675998 169904
rect 675956 169250 675984 169895
rect 676048 169658 676076 170711
rect 676036 169652 676088 169658
rect 676036 169594 676088 169600
rect 676034 169552 676090 169561
rect 676034 169487 676090 169496
rect 675944 169244 675996 169250
rect 675944 169186 675996 169192
rect 675942 169144 675998 169153
rect 675942 169079 675998 169088
rect 675956 168774 675984 169079
rect 675944 168768 675996 168774
rect 675850 168736 675906 168745
rect 675944 168710 675996 168716
rect 676048 168706 676076 169487
rect 675850 168671 675906 168680
rect 676036 168700 676088 168706
rect 675864 168570 675892 168671
rect 676036 168642 676088 168648
rect 675852 168564 675904 168570
rect 675852 168506 675904 168512
rect 676034 168328 676090 168337
rect 676034 168263 676036 168272
rect 676088 168263 676090 168272
rect 676036 168234 676088 168240
rect 676034 167920 676090 167929
rect 676034 167855 676036 167864
rect 676088 167855 676090 167864
rect 676036 167826 676088 167832
rect 676034 167512 676090 167521
rect 676034 167447 676036 167456
rect 676088 167447 676090 167456
rect 676036 167418 676088 167424
rect 675760 161016 675812 161022
rect 675760 160958 675812 160964
rect 675760 160812 675812 160818
rect 675760 160754 675812 160760
rect 675772 160344 675800 160754
rect 675208 160064 675260 160070
rect 675208 160006 675260 160012
rect 675392 160064 675444 160070
rect 675392 160006 675444 160012
rect 675404 159664 675432 160006
rect 675484 159384 675536 159390
rect 675484 159326 675536 159332
rect 675496 159052 675524 159326
rect 674840 157752 674892 157758
rect 674840 157694 674892 157700
rect 675484 157752 675536 157758
rect 675484 157694 675536 157700
rect 675496 157216 675524 157694
rect 675392 156936 675444 156942
rect 675392 156878 675444 156884
rect 675404 156643 675432 156878
rect 675392 156528 675444 156534
rect 675392 156470 675444 156476
rect 675404 155992 675432 156470
rect 674748 155916 674800 155922
rect 674748 155858 674800 155864
rect 675484 155916 675536 155922
rect 675484 155858 675536 155864
rect 675496 155380 675524 155858
rect 675392 153400 675444 153406
rect 675392 153342 675444 153348
rect 675404 152864 675432 153342
rect 674012 152788 674064 152794
rect 674012 152730 674064 152736
rect 675392 152788 675444 152794
rect 675392 152730 675444 152736
rect 675404 152320 675432 152730
rect 673736 152040 673788 152046
rect 673736 151982 673788 151988
rect 675392 152040 675444 152046
rect 675392 151982 675444 151988
rect 675404 151675 675432 151982
rect 673644 151428 673696 151434
rect 673644 151370 673696 151376
rect 675392 151428 675444 151434
rect 675392 151370 675444 151376
rect 675404 151028 675432 151370
rect 673552 150408 673604 150414
rect 673552 150350 673604 150356
rect 675392 150408 675444 150414
rect 675392 150350 675444 150356
rect 675404 149835 675432 150350
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675758 146296 675814 146305
rect 675758 146231 675814 146240
rect 675772 146132 675800 146231
rect 704372 134360 704424 134366
rect 704168 134308 704372 134314
rect 704168 134302 704424 134308
rect 704168 134286 704412 134302
rect 708432 134298 708768 134314
rect 704464 134292 704516 134298
rect 704464 134234 704516 134240
rect 708420 134292 708768 134298
rect 708472 134286 708768 134292
rect 708892 134286 709228 134314
rect 708420 134234 708472 134240
rect 703818 134192 703874 134201
rect 703708 134150 703818 134178
rect 703818 134127 703874 134136
rect 704476 133906 704504 134234
rect 707500 134224 707552 134230
rect 704628 134150 704872 134178
rect 705088 134150 705424 134178
rect 705548 134150 705884 134178
rect 706008 134150 706344 134178
rect 704168 133878 704504 133906
rect 704844 133890 704872 134150
rect 705292 134088 705344 134094
rect 705292 134030 705344 134036
rect 705304 133906 705332 134030
rect 704832 133884 704884 133890
rect 705088 133878 705332 133906
rect 705396 133890 705424 134150
rect 705752 134088 705804 134094
rect 705752 134030 705804 134036
rect 705764 133906 705792 134030
rect 705856 134026 705884 134150
rect 706212 134088 706264 134094
rect 706212 134030 706264 134036
rect 705844 134020 705896 134026
rect 705844 133962 705896 133968
rect 706224 133906 706252 134030
rect 706316 133958 706344 134150
rect 706592 134150 706928 134178
rect 707052 134162 707388 134178
rect 708512 134224 708564 134230
rect 707552 134172 707848 134178
rect 707500 134166 707848 134172
rect 707040 134156 707388 134162
rect 706592 134094 706620 134150
rect 707092 134150 707388 134156
rect 707512 134150 707848 134166
rect 707972 134150 708308 134178
rect 708512 134166 708564 134172
rect 707040 134098 707092 134104
rect 706580 134088 706632 134094
rect 706580 134030 706632 134036
rect 705384 133884 705436 133890
rect 704832 133826 704884 133832
rect 705548 133878 705792 133906
rect 706008 133878 706252 133906
rect 706304 133952 706356 133958
rect 706304 133894 706356 133900
rect 706454 133892 706482 134028
rect 707040 134020 707092 134026
rect 707040 133962 707092 133968
rect 706580 133952 706632 133958
rect 707052 133906 707080 133962
rect 706632 133900 706928 133906
rect 706580 133894 706928 133900
rect 706592 133878 706928 133894
rect 707052 133878 707388 133906
rect 707512 133890 707848 133906
rect 707500 133884 707848 133890
rect 705384 133826 705436 133832
rect 707552 133878 707848 133884
rect 707500 133826 707552 133832
rect 707972 133822 708000 134150
rect 708524 133906 708552 134166
rect 708524 133878 708768 133906
rect 704924 133816 704976 133822
rect 704628 133764 704924 133770
rect 704628 133758 704976 133764
rect 707960 133816 708012 133822
rect 707960 133758 708012 133764
rect 704628 133742 704964 133758
rect 708064 133754 708308 133770
rect 708052 133748 708308 133754
rect 708104 133742 708308 133748
rect 708052 133690 708104 133696
rect 708892 133686 708920 134286
rect 709062 134192 709118 134201
rect 709062 134127 709118 134136
rect 709076 133906 709104 134127
rect 709076 133878 709228 133906
rect 704004 133680 704056 133686
rect 703708 133628 704004 133634
rect 703708 133622 704056 133628
rect 708880 133680 708932 133686
rect 708880 133622 708932 133628
rect 703708 133606 704044 133622
rect 676126 133104 676182 133113
rect 676126 133039 676182 133048
rect 676034 132968 676090 132977
rect 676034 132903 676090 132912
rect 676048 132666 676076 132903
rect 676140 132802 676168 133039
rect 676220 132932 676272 132938
rect 676220 132874 676272 132880
rect 676128 132796 676180 132802
rect 676128 132738 676180 132744
rect 676232 132705 676260 132874
rect 676218 132696 676274 132705
rect 676036 132660 676088 132666
rect 676218 132631 676274 132640
rect 676036 132602 676088 132608
rect 676220 132320 676272 132326
rect 676218 132288 676220 132297
rect 676272 132288 676274 132297
rect 676218 132223 676274 132232
rect 676034 131744 676090 131753
rect 676034 131679 676036 131688
rect 676088 131679 676090 131688
rect 676036 131650 676088 131656
rect 673368 131504 673420 131510
rect 676220 131504 676272 131510
rect 673368 131446 673420 131452
rect 676218 131472 676220 131481
rect 676272 131472 676274 131481
rect 676218 131407 676274 131416
rect 676034 130928 676090 130937
rect 676034 130863 676036 130872
rect 676088 130863 676090 130872
rect 676036 130834 676088 130840
rect 676220 130688 676272 130694
rect 676218 130656 676220 130665
rect 676272 130656 676274 130665
rect 676218 130591 676274 130600
rect 676034 130112 676090 130121
rect 676034 130047 676036 130056
rect 676088 130047 676090 130056
rect 676036 130018 676088 130024
rect 676036 129736 676088 129742
rect 676034 129704 676036 129713
rect 676088 129704 676090 129713
rect 676034 129639 676090 129648
rect 676220 129464 676272 129470
rect 676218 129432 676220 129441
rect 676272 129432 676274 129441
rect 676218 129367 676274 129376
rect 676034 128888 676090 128897
rect 676034 128823 676090 128832
rect 675758 128072 675814 128081
rect 675758 128007 675814 128016
rect 674472 127764 674524 127770
rect 674472 127706 674524 127712
rect 673644 127084 673696 127090
rect 673644 127026 673696 127032
rect 673460 124908 673512 124914
rect 673460 124850 673512 124856
rect 673182 122904 673238 122913
rect 673182 122839 673238 122848
rect 672908 122732 672960 122738
rect 672908 122674 672960 122680
rect 672920 110945 672948 122674
rect 672906 110936 672962 110945
rect 672906 110871 672962 110880
rect 672446 105904 672502 105913
rect 672446 105839 672502 105848
rect 673472 105194 673500 124850
rect 673552 124432 673604 124438
rect 673552 124374 673604 124380
rect 673564 107030 673592 124374
rect 673656 108254 673684 127026
rect 673828 123276 673880 123282
rect 673828 123218 673880 123224
rect 673736 121508 673788 121514
rect 673736 121450 673788 121456
rect 673644 108248 673696 108254
rect 673644 108190 673696 108196
rect 673552 107024 673604 107030
rect 673552 106966 673604 106972
rect 673748 106418 673776 121450
rect 673840 107574 673868 123218
rect 674484 114238 674512 127706
rect 674564 127016 674616 127022
rect 674564 126958 674616 126964
rect 674472 114232 674524 114238
rect 674472 114174 674524 114180
rect 674576 112402 674604 126958
rect 674748 124500 674800 124506
rect 674748 124442 674800 124448
rect 674656 124364 674708 124370
rect 674656 124306 674708 124312
rect 674564 112396 674616 112402
rect 674564 112338 674616 112344
rect 674668 111178 674696 124306
rect 674760 111926 674788 124442
rect 675116 124296 675168 124302
rect 675116 124238 675168 124244
rect 674748 111920 674800 111926
rect 674748 111862 674800 111868
rect 674656 111172 674708 111178
rect 674656 111114 674708 111120
rect 675128 110702 675156 124238
rect 675208 124228 675260 124234
rect 675208 124170 675260 124176
rect 675220 115054 675248 124170
rect 675772 115802 675800 128007
rect 676048 127770 676076 128823
rect 676036 127764 676088 127770
rect 676036 127706 676088 127712
rect 676034 127664 676090 127673
rect 676034 127599 676090 127608
rect 675942 127256 675998 127265
rect 675942 127191 675998 127200
rect 675956 127090 675984 127191
rect 675944 127084 675996 127090
rect 675944 127026 675996 127032
rect 676048 127022 676076 127599
rect 676036 127016 676088 127022
rect 676036 126958 676088 126964
rect 676034 126440 676090 126449
rect 676034 126375 676090 126384
rect 675942 126032 675998 126041
rect 675942 125967 675998 125976
rect 675850 125216 675906 125225
rect 675850 125151 675906 125160
rect 675864 124914 675892 125151
rect 675852 124908 675904 124914
rect 675852 124850 675904 124856
rect 675850 124808 675906 124817
rect 675850 124743 675906 124752
rect 675864 124438 675892 124743
rect 675956 124506 675984 125967
rect 675944 124500 675996 124506
rect 675944 124442 675996 124448
rect 675852 124432 675904 124438
rect 675852 124374 675904 124380
rect 675942 124400 675998 124409
rect 675942 124335 675998 124344
rect 675956 124302 675984 124335
rect 675944 124296 675996 124302
rect 675944 124238 675996 124244
rect 676048 124234 676076 126375
rect 676126 125352 676182 125361
rect 676126 125287 676182 125296
rect 676140 124370 676168 125287
rect 676128 124364 676180 124370
rect 676128 124306 676180 124312
rect 676036 124228 676088 124234
rect 676036 124170 676088 124176
rect 676034 123992 676090 124001
rect 676034 123927 676090 123936
rect 675942 123584 675998 123593
rect 675942 123519 675998 123528
rect 675956 121514 675984 123519
rect 676048 123282 676076 123927
rect 676036 123276 676088 123282
rect 676036 123218 676088 123224
rect 676034 123176 676090 123185
rect 676034 123111 676036 123120
rect 676088 123111 676090 123120
rect 676036 123082 676088 123088
rect 676034 122768 676090 122777
rect 676034 122703 676036 122712
rect 676088 122703 676090 122712
rect 676036 122674 676088 122680
rect 676034 122360 676090 122369
rect 676034 122295 676036 122304
rect 676088 122295 676090 122304
rect 676036 122266 676088 122272
rect 675944 121508 675996 121514
rect 675944 121450 675996 121456
rect 675760 115796 675812 115802
rect 675760 115738 675812 115744
rect 675760 115592 675812 115598
rect 675760 115534 675812 115540
rect 675772 115124 675800 115534
rect 675208 115048 675260 115054
rect 675208 114990 675260 114996
rect 675392 115048 675444 115054
rect 675392 114990 675444 114996
rect 675404 114479 675432 114990
rect 675392 114232 675444 114238
rect 675392 114174 675444 114180
rect 675404 113832 675432 114174
rect 675392 112396 675444 112402
rect 675392 112338 675444 112344
rect 675404 111996 675432 112338
rect 675392 111920 675444 111926
rect 675392 111862 675444 111868
rect 675404 111452 675432 111862
rect 675392 111172 675444 111178
rect 675392 111114 675444 111120
rect 675404 110772 675432 111114
rect 675116 110696 675168 110702
rect 675116 110638 675168 110644
rect 675392 110696 675444 110702
rect 675392 110638 675444 110644
rect 675404 110160 675432 110638
rect 675484 108248 675536 108254
rect 675484 108190 675536 108196
rect 675496 107644 675524 108190
rect 673828 107568 673880 107574
rect 673828 107510 673880 107516
rect 675392 107568 675444 107574
rect 675392 107510 675444 107516
rect 675404 107100 675432 107510
rect 675392 107024 675444 107030
rect 675392 106966 675444 106972
rect 675404 106488 675432 106966
rect 673736 106412 673788 106418
rect 673736 106354 673788 106360
rect 675392 106412 675444 106418
rect 675392 106354 675444 106360
rect 675404 105808 675432 106354
rect 673460 105188 673512 105194
rect 673460 105130 673512 105136
rect 675484 105188 675536 105194
rect 675484 105130 675536 105136
rect 675496 104652 675524 105130
rect 675758 103320 675814 103329
rect 675758 103255 675814 103264
rect 675772 102816 675800 103255
rect 671986 102504 672042 102513
rect 671986 102439 672042 102448
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 670882 100872 670938 100881
rect 670882 100807 670938 100816
rect 646320 46912 646372 46918
rect 646320 46854 646372 46860
rect 666560 46912 666612 46918
rect 666560 46854 666612 46860
rect 646332 45121 646360 46854
rect 646318 45112 646374 45121
rect 646318 45047 646374 45056
rect 642638 41304 642694 41313
rect 642638 41239 642694 41248
rect 475660 38548 475712 38554
rect 475660 38490 475712 38496
rect 514024 38548 514076 38554
rect 514024 38490 514076 38496
rect 231030 15192 231086 15201
rect 231030 15127 231086 15136
rect 230938 12200 230994 12209
rect 230938 12135 230994 12144
rect 230662 9208 230718 9217
rect 230662 9143 230718 9152
rect 230570 7712 230626 7721
rect 230570 7647 230626 7656
rect 230386 6216 230442 6225
rect 230386 6151 230442 6160
<< via2 >>
rect 425978 1006052 426034 1006088
rect 425978 1006032 425980 1006052
rect 425980 1006032 426032 1006052
rect 426032 1006032 426034 1006052
rect 424322 1005916 424378 1005952
rect 424322 1005896 424324 1005916
rect 424324 1005896 424376 1005916
rect 424376 1005896 424378 1005916
rect 423862 1005796 423864 1005816
rect 423864 1005796 423916 1005816
rect 423916 1005796 423918 1005816
rect 423862 1005760 423918 1005796
rect 356058 1005644 356114 1005680
rect 356058 1005624 356060 1005644
rect 356060 1005624 356112 1005644
rect 356112 1005624 356114 1005644
rect 356886 1005524 356888 1005544
rect 356888 1005524 356940 1005544
rect 356940 1005524 356942 1005544
rect 356886 1005488 356942 1005524
rect 160282 1005388 160284 1005408
rect 160284 1005388 160336 1005408
rect 160336 1005388 160338 1005408
rect 86590 995696 86646 995752
rect 87786 995560 87842 995616
rect 81622 995424 81678 995480
rect 81990 995288 82046 995344
rect 85302 995424 85358 995480
rect 80702 995152 80758 995208
rect 84474 995152 84530 995208
rect 80150 993792 80206 993848
rect 78310 993656 78366 993712
rect 106462 1005236 106518 1005272
rect 106462 1005216 106464 1005236
rect 106464 1005216 106516 1005236
rect 106516 1005216 106518 1005236
rect 109314 1005252 109316 1005272
rect 109316 1005252 109368 1005272
rect 109368 1005252 109370 1005272
rect 109314 1005216 109370 1005252
rect 105634 1005116 105636 1005136
rect 105636 1005116 105688 1005136
rect 105688 1005116 105690 1005136
rect 105634 1005080 105690 1005116
rect 108026 1004844 108028 1004864
rect 108028 1004844 108080 1004864
rect 108080 1004844 108082 1004864
rect 108026 1004808 108082 1004844
rect 109682 1004844 109684 1004864
rect 109684 1004844 109736 1004864
rect 109736 1004844 109738 1004864
rect 109682 1004808 109738 1004844
rect 114650 1004828 114706 1004864
rect 114650 1004808 114652 1004828
rect 114652 1004808 114704 1004828
rect 114704 1004808 114706 1004828
rect 98274 1004672 98330 1004728
rect 98642 1004672 98698 1004728
rect 99470 1004708 99472 1004728
rect 99472 1004708 99524 1004728
rect 99524 1004708 99526 1004728
rect 99470 1004672 99526 1004708
rect 108854 1004692 108910 1004728
rect 108854 1004672 108856 1004692
rect 108856 1004672 108908 1004692
rect 108908 1004672 108910 1004692
rect 92754 995016 92810 995072
rect 41786 968768 41842 968824
rect 41786 965096 41842 965152
rect 41786 963328 41842 963384
rect 35806 949456 35862 949512
rect 41510 943880 41566 943936
rect 41786 943084 41842 943120
rect 41786 943064 41788 943084
rect 41788 943064 41840 943084
rect 41840 943064 41842 943084
rect 41786 942692 41788 942712
rect 41788 942692 41840 942712
rect 41840 942692 41842 942712
rect 41786 942656 41842 942692
rect 41878 942248 41934 942304
rect 41786 941468 41788 941488
rect 41788 941468 41840 941488
rect 41840 941468 41842 941488
rect 41786 941432 41842 941468
rect 41694 940480 41750 940536
rect 41970 941840 42026 941896
rect 41878 941024 41934 941080
rect 41786 936536 41842 936592
rect 35806 934904 35862 934960
rect 35714 934496 35770 934552
rect 35622 934088 35678 934144
rect 41970 940208 42026 940264
rect 41970 938440 42026 938496
rect 42338 938984 42394 939040
rect 42246 938168 42302 938224
rect 41510 921984 41566 922040
rect 41786 933272 41842 933328
rect 41786 932476 41842 932512
rect 41786 932456 41788 932476
rect 41788 932456 41840 932476
rect 41840 932456 41842 932476
rect 41786 817672 41842 817728
rect 41786 817300 41788 817320
rect 41788 817300 41840 817320
rect 41840 817300 41842 817320
rect 41786 817264 41842 817300
rect 42798 938576 42854 938632
rect 42982 939800 43038 939856
rect 42890 933680 42946 933736
rect 42798 921984 42854 922040
rect 41970 816448 42026 816504
rect 41694 815768 41750 815824
rect 41142 814238 41198 814294
rect 42706 816040 42762 816096
rect 41970 814136 42026 814192
rect 41878 814000 41934 814056
rect 42338 814000 42394 814056
rect 41786 813592 41842 813648
rect 41786 811552 41842 811608
rect 41970 811144 42026 811200
rect 41786 808288 41842 808344
rect 41878 807900 41934 807936
rect 41878 807880 41880 807900
rect 41880 807880 41932 807900
rect 41932 807880 41934 807900
rect 41786 807472 41842 807528
rect 41786 806676 41842 806712
rect 41786 806656 41788 806676
rect 41788 806656 41840 806676
rect 41840 806656 41842 806676
rect 42614 809512 42670 809568
rect 41510 774732 41512 774752
rect 41512 774732 41564 774752
rect 41564 774732 41566 774752
rect 41510 774696 41566 774732
rect 41786 774016 41842 774072
rect 41510 773916 41512 773936
rect 41512 773916 41564 773936
rect 41564 773916 41566 773936
rect 41510 773880 41566 773916
rect 41510 773472 41566 773528
rect 42154 771976 42210 772032
rect 41878 767896 41934 767952
rect 41510 764088 41566 764144
rect 30378 763680 30434 763736
rect 30378 763272 30434 763328
rect 41510 763292 41566 763328
rect 41510 763272 41512 763292
rect 41512 763272 41564 763292
rect 41564 763272 41566 763292
rect 42062 766672 42118 766728
rect 42430 770752 42486 770808
rect 42706 769936 42762 769992
rect 41970 757016 42026 757072
rect 42062 754024 42118 754080
rect 41786 731348 41788 731368
rect 41788 731348 41840 731368
rect 41840 731348 41842 731368
rect 41786 731312 41842 731348
rect 39394 731040 39450 731096
rect 41510 731076 41512 731096
rect 41512 731076 41564 731096
rect 41564 731076 41566 731096
rect 41510 731040 41566 731076
rect 41510 730668 41512 730688
rect 41512 730668 41564 730688
rect 41564 730668 41566 730688
rect 41510 730632 41566 730668
rect 39394 729816 39450 729872
rect 43074 937352 43130 937408
rect 43258 937760 43314 937816
rect 43166 936128 43222 936184
rect 43350 935720 43406 935776
rect 43994 927152 44050 927208
rect 43534 815224 43590 815280
rect 43442 814816 43498 814872
rect 43350 813184 43406 813240
rect 42890 812776 42946 812832
rect 42982 812368 43038 812424
rect 43074 811960 43130 812016
rect 43258 809104 43314 809160
rect 43810 810736 43866 810792
rect 43626 808696 43682 808752
rect 42890 771160 42946 771216
rect 43074 769528 43130 769584
rect 42890 764632 42946 764688
rect 42798 730088 42854 730144
rect 41510 729408 41566 729464
rect 43166 768304 43222 768360
rect 43258 767488 43314 767544
rect 43166 766264 43222 766320
rect 43442 772384 43498 772440
rect 43902 809920 43958 809976
rect 44086 810328 44142 810384
rect 43534 770344 43590 770400
rect 43718 769120 43774 769176
rect 43534 765856 43590 765912
rect 43442 765040 43498 765096
rect 44086 768712 44142 768768
rect 44086 767080 44142 767136
rect 43994 765448 44050 765504
rect 44178 730088 44234 730144
rect 43350 729680 43406 729736
rect 41786 728884 41842 728920
rect 41786 728864 41788 728884
rect 41788 728864 41840 728884
rect 41840 728864 41842 728884
rect 39394 728184 39450 728240
rect 43718 728456 43774 728512
rect 42522 727232 42578 727288
rect 43626 726824 43682 726880
rect 43074 726416 43130 726472
rect 41878 724784 41934 724840
rect 41326 723696 41382 723752
rect 30378 720432 30434 720488
rect 30378 720024 30434 720080
rect 41510 720840 41566 720896
rect 41510 720044 41566 720080
rect 41510 720024 41512 720044
rect 41512 720024 41564 720044
rect 41564 720024 41566 720044
rect 42890 724376 42946 724432
rect 42798 723152 42854 723208
rect 42982 723560 43038 723616
rect 43166 726008 43222 726064
rect 43534 725600 43590 725656
rect 43350 725192 43406 725248
rect 43258 721520 43314 721576
rect 41510 688372 41512 688392
rect 41512 688372 41564 688392
rect 41564 688372 41566 688392
rect 41510 688336 41566 688372
rect 41786 687692 41788 687712
rect 41788 687692 41840 687712
rect 41840 687692 41842 687712
rect 41786 687656 41842 687692
rect 41694 687520 41750 687576
rect 42798 685208 42854 685264
rect 43442 722744 43498 722800
rect 43902 722336 43958 722392
rect 44086 721928 44142 721984
rect 44178 686432 44234 686488
rect 44362 727640 44418 727696
rect 44270 686024 44326 686080
rect 43442 685616 43498 685672
rect 43166 684800 43222 684856
rect 41694 681808 41750 681864
rect 41878 681536 41934 681592
rect 41786 678680 41842 678736
rect 41786 677864 41842 677920
rect 41786 677068 41842 677104
rect 41786 677048 41788 677068
rect 41788 677048 41840 677068
rect 41840 677048 41842 677068
rect 41970 678272 42026 678328
rect 41510 645124 41512 645144
rect 41512 645124 41564 645144
rect 41564 645124 41566 645144
rect 41510 645088 41566 645124
rect 41510 644716 41512 644736
rect 41512 644716 41564 644736
rect 41564 644716 41566 644736
rect 41510 644680 41566 644716
rect 41510 644272 41566 644328
rect 41510 643476 41566 643512
rect 41510 643456 41512 643476
rect 41512 643456 41564 643476
rect 41564 643456 41566 643476
rect 42890 684392 42946 684448
rect 43350 683576 43406 683632
rect 42982 682760 43038 682816
rect 43166 680720 43222 680776
rect 42798 641824 42854 641880
rect 44362 683984 44418 684040
rect 43994 683168 44050 683224
rect 43810 682352 43866 682408
rect 43718 681128 43774 681184
rect 43626 680312 43682 680368
rect 43534 679496 43590 679552
rect 43902 679904 43958 679960
rect 44086 679088 44142 679144
rect 43442 643048 43498 643104
rect 44270 641960 44326 642016
rect 42890 641008 42946 641064
rect 43074 640328 43130 640384
rect 42798 639376 42854 639432
rect 41786 638356 41842 638412
rect 33046 634888 33102 634944
rect 30378 634072 30434 634128
rect 30378 633664 30434 633720
rect 41510 634480 41566 634536
rect 41510 633684 41566 633720
rect 41510 633664 41512 633684
rect 41512 633664 41564 633684
rect 41564 633664 41566 633684
rect 42982 637744 43038 637800
rect 42890 636520 42946 636576
rect 43534 639784 43590 639840
rect 43166 638968 43222 639024
rect 43442 638560 43498 638616
rect 43350 636112 43406 636168
rect 43258 635296 43314 635352
rect 43718 637608 43774 637664
rect 43626 635704 43682 635760
rect 43810 636928 43866 636984
rect 41510 601876 41512 601896
rect 41512 601876 41564 601896
rect 41564 601876 41566 601896
rect 41510 601840 41566 601876
rect 41510 601468 41512 601488
rect 41512 601468 41564 601488
rect 41564 601468 41566 601488
rect 41510 601432 41566 601468
rect 43074 600480 43130 600536
rect 41510 599836 41512 599856
rect 41512 599836 41564 599856
rect 41564 599836 41566 599856
rect 41510 599800 41566 599836
rect 41510 599004 41566 599040
rect 41510 598984 41512 599004
rect 41512 598984 41564 599004
rect 41564 598984 41566 599004
rect 42430 598032 42486 598088
rect 41878 595176 41934 595232
rect 41326 594088 41382 594144
rect 29918 591232 29974 591288
rect 29918 590824 29974 590880
rect 30378 590824 30434 590880
rect 30378 590416 30434 590472
rect 42890 596808 42946 596864
rect 42798 593544 42854 593600
rect 42706 591912 42762 591968
rect 42982 593952 43038 594008
rect 41510 558764 41512 558784
rect 41512 558764 41564 558784
rect 41564 558764 41566 558784
rect 41510 558728 41566 558764
rect 41786 558048 41842 558104
rect 41510 557912 41566 557968
rect 43258 596400 43314 596456
rect 43166 594768 43222 594824
rect 43258 592320 43314 592376
rect 43074 556824 43130 556880
rect 44454 642232 44510 642288
rect 44362 600072 44418 600128
rect 44638 641416 44694 641472
rect 44270 598440 44326 598496
rect 44638 597624 44694 597680
rect 43810 597216 43866 597272
rect 43442 595584 43498 595640
rect 43626 593136 43682 593192
rect 43718 592728 43774 592784
rect 43902 595992 43958 596048
rect 43350 556416 43406 556472
rect 43166 554376 43222 554432
rect 43534 553968 43590 554024
rect 42706 553560 42762 553616
rect 41786 551928 41842 551984
rect 41602 548936 41658 548992
rect 41510 548528 41566 548584
rect 41418 548120 41474 548176
rect 30470 547712 30526 547768
rect 30470 547304 30526 547360
rect 41418 547324 41474 547360
rect 41418 547304 41420 547324
rect 41420 547304 41472 547324
rect 41472 547304 41474 547324
rect 43350 553152 43406 553208
rect 42982 552744 43038 552800
rect 42890 550296 42946 550352
rect 43166 552336 43222 552392
rect 43074 551112 43130 551168
rect 43442 549888 43498 549944
rect 43626 551520 43682 551576
rect 43718 550704 43774 550760
rect 43810 549480 43866 549536
rect 44086 540912 44142 540968
rect 43994 540776 44050 540832
rect 41786 430888 41842 430944
rect 43534 429664 43590 429720
rect 41786 426808 41842 426864
rect 43258 426400 43314 426456
rect 42798 425992 42854 426048
rect 41878 424360 41934 424416
rect 41786 421504 41842 421560
rect 42522 421096 42578 421152
rect 42890 425584 42946 425640
rect 42798 411212 42854 411268
rect 41510 387948 41512 387968
rect 41512 387948 41564 387968
rect 41564 387948 41566 387968
rect 41510 387912 41566 387948
rect 41786 387232 41842 387288
rect 41510 387132 41512 387152
rect 41512 387132 41564 387152
rect 41564 387132 41566 387152
rect 41510 387096 41566 387132
rect 43166 425176 43222 425232
rect 42982 422728 43038 422784
rect 43442 424768 43498 424824
rect 43350 422320 43406 422376
rect 43994 429256 44050 429312
rect 43718 428440 43774 428496
rect 43626 423136 43682 423192
rect 43534 411440 43590 411496
rect 42798 386008 42854 386064
rect 43902 423952 43958 424008
rect 43810 423544 43866 423600
rect 43994 421912 44050 421968
rect 43718 385600 43774 385656
rect 43534 385192 43590 385248
rect 42982 383152 43038 383208
rect 42706 382744 42762 382800
rect 42338 381112 42394 381168
rect 41510 377712 41566 377768
rect 41418 377304 41474 377360
rect 30470 376896 30526 376952
rect 30470 376488 30526 376544
rect 41418 376508 41474 376544
rect 41418 376488 41420 376508
rect 41420 376488 41472 376508
rect 41472 376488 41474 376508
rect 42890 381928 42946 381984
rect 42798 381520 42854 381576
rect 43074 379480 43130 379536
rect 43258 379072 43314 379128
rect 43166 378256 43222 378312
rect 43442 378664 43498 378720
rect 41786 355680 41842 355736
rect 33046 351872 33102 351928
rect 41510 344276 41566 344312
rect 41510 344256 41512 344276
rect 41512 344256 41564 344276
rect 41564 344256 41566 344276
rect 41786 344156 41788 344176
rect 41788 344156 41840 344176
rect 41840 344156 41842 344176
rect 41786 344120 41842 344156
rect 43626 380704 43682 380760
rect 43718 380296 43774 380352
rect 43810 379888 43866 379944
rect 33046 343032 33102 343088
rect 41602 343884 41604 343904
rect 41604 343884 41656 343904
rect 41656 343884 41658 343904
rect 41602 343848 41658 343884
rect 41786 343340 41788 343360
rect 41788 343340 41840 343360
rect 41840 343340 41842 343360
rect 41786 343304 41842 343340
rect 41510 342624 41566 342680
rect 43258 342080 43314 342136
rect 32678 339768 32734 339824
rect 32586 338544 32642 338600
rect 30378 333648 30434 333704
rect 30378 333240 30434 333296
rect 32770 338136 32826 338192
rect 33046 337728 33102 337784
rect 32954 336096 33010 336152
rect 32862 335688 32918 335744
rect 32770 329840 32826 329896
rect 43074 335552 43130 335608
rect 42982 335144 43038 335200
rect 41510 334056 41566 334112
rect 41510 333260 41566 333296
rect 41510 333240 41512 333260
rect 41512 333240 41564 333260
rect 41564 333240 41566 333260
rect 32586 329704 32642 329760
rect 41786 319912 41842 319968
rect 43166 334736 43222 334792
rect 41970 316920 42026 316976
rect 42154 315968 42210 316024
rect 42154 315424 42210 315480
rect 42154 313792 42210 313848
rect 41786 313112 41842 313168
rect 41786 312296 41842 312352
rect 41510 301588 41512 301608
rect 41512 301588 41564 301608
rect 41564 301588 41566 301608
rect 41510 301552 41566 301588
rect 41786 300908 41788 300928
rect 41788 300908 41840 300928
rect 41840 300908 41842 300928
rect 41786 300872 41842 300908
rect 44270 341672 44326 341728
rect 44178 340856 44234 340912
rect 43258 299240 43314 299296
rect 43534 298832 43590 298888
rect 32770 296792 32826 296848
rect 32586 295976 32642 296032
rect 32678 294752 32734 294808
rect 32586 285640 32642 285696
rect 35806 296384 35862 296440
rect 32862 295160 32918 295216
rect 32770 285776 32826 285832
rect 33046 294344 33102 294400
rect 32954 293936 33010 293992
rect 42890 293528 42946 293584
rect 33046 285912 33102 285968
rect 42982 293120 43038 293176
rect 43166 292712 43222 292768
rect 43074 292304 43130 292360
rect 43350 291488 43406 291544
rect 41970 272312 42026 272368
rect 42154 270408 42210 270464
rect 42154 270000 42210 270056
rect 42154 269184 42210 269240
rect 41510 258340 41512 258360
rect 41512 258340 41564 258360
rect 41564 258340 41566 258360
rect 41510 258304 41566 258340
rect 41786 257624 41842 257680
rect 41510 257524 41512 257544
rect 41512 257524 41564 257544
rect 41564 257524 41566 257544
rect 41510 257488 41566 257524
rect 41786 256844 41788 256864
rect 41788 256844 41840 256864
rect 41840 256844 41842 256864
rect 41786 256808 41842 256844
rect 44270 340040 44326 340096
rect 44362 299648 44418 299704
rect 44270 298016 44326 298072
rect 44178 297200 44234 297256
rect 43626 291896 43682 291952
rect 43534 255992 43590 256048
rect 43442 255584 43498 255640
rect 42706 253544 42762 253600
rect 31666 253000 31722 253056
rect 33046 251776 33102 251832
rect 32770 250552 32826 250608
rect 32862 250144 32918 250200
rect 32954 249736 33010 249792
rect 38290 248104 38346 248160
rect 41510 247716 41566 247752
rect 41510 247696 41512 247716
rect 41512 247696 41564 247716
rect 41564 247696 41566 247716
rect 41510 247308 41566 247344
rect 41510 247288 41512 247308
rect 41512 247288 41564 247308
rect 41564 247288 41566 247308
rect 41510 246900 41566 246936
rect 41510 246880 41512 246900
rect 41512 246880 41564 246900
rect 41564 246880 41566 246900
rect 42890 252320 42946 252376
rect 43258 249464 43314 249520
rect 43074 248648 43130 248704
rect 43350 249056 43406 249112
rect 41970 225936 42026 225992
rect 41510 215056 41566 215112
rect 41418 214648 41474 214704
rect 41602 214240 41658 214296
rect 41510 213868 41512 213888
rect 41512 213868 41564 213888
rect 41564 213868 41566 213888
rect 41510 213832 41566 213868
rect 43718 251504 43774 251560
rect 43810 251096 43866 251152
rect 41510 213016 41566 213072
rect 45926 255176 45982 255232
rect 45742 254360 45798 254416
rect 46202 340856 46258 340912
rect 46110 298424 46166 298480
rect 46110 291080 46166 291136
rect 46478 641416 46534 641472
rect 46478 600072 46534 600128
rect 46386 340040 46442 340096
rect 46386 290672 46442 290728
rect 46570 598440 46626 598496
rect 46662 419872 46718 419928
rect 58438 975976 58494 976032
rect 57978 962920 58034 962976
rect 58438 949864 58494 949920
rect 58438 936944 58494 937000
rect 58438 923752 58494 923808
rect 58070 910696 58126 910752
rect 48318 300056 48374 300112
rect 48226 297608 48282 297664
rect 46846 290264 46902 290320
rect 48870 590688 48926 590744
rect 58530 897776 58586 897832
rect 58438 884720 58494 884776
rect 58438 871664 58494 871720
rect 58438 858608 58494 858664
rect 58438 845552 58494 845608
rect 57978 832496 58034 832552
rect 53838 816856 53894 816912
rect 59174 819440 59230 819496
rect 58438 806520 58494 806576
rect 58070 793464 58126 793520
rect 58438 780408 58494 780464
rect 58438 767372 58494 767408
rect 58438 767352 58440 767372
rect 58440 767352 58492 767372
rect 58492 767352 58494 767372
rect 58346 754296 58402 754352
rect 58438 741240 58494 741296
rect 58438 728184 58494 728240
rect 58438 715264 58494 715320
rect 58162 702208 58218 702264
rect 58438 689152 58494 689208
rect 58438 676096 58494 676152
rect 58438 663040 58494 663096
rect 59174 649984 59230 650040
rect 58438 637064 58494 637120
rect 58438 624008 58494 624064
rect 58438 610952 58494 611008
rect 53838 600888 53894 600944
rect 59174 597896 59230 597952
rect 58438 584840 58494 584896
rect 58438 571784 58494 571840
rect 57978 558728 58034 558784
rect 59174 545808 59230 545864
rect 51262 430480 51318 430536
rect 59266 532752 59322 532808
rect 58438 519696 58494 519752
rect 58438 506640 58494 506696
rect 57978 493584 58034 493640
rect 58438 480528 58494 480584
rect 58622 467472 58678 467528
rect 53838 430072 53894 430128
rect 59174 454552 59230 454608
rect 58438 441496 58494 441552
rect 57978 428440 58034 428496
rect 58438 415384 58494 415440
rect 58438 402328 58494 402384
rect 57978 389272 58034 389328
rect 62118 386280 62174 386336
rect 62026 383424 62082 383480
rect 62302 939392 62358 939448
rect 62210 383016 62266 383072
rect 58438 376216 58494 376272
rect 58438 363296 58494 363352
rect 58438 350240 58494 350296
rect 58438 337184 58494 337240
rect 58162 324128 58218 324184
rect 53838 300464 53894 300520
rect 46938 212472 46994 212528
rect 45650 212064 45706 212120
rect 45466 211248 45522 211304
rect 32954 209752 33010 209808
rect 31850 204856 31906 204912
rect 31666 204040 31722 204096
rect 33046 208120 33102 208176
rect 42890 206760 42946 206816
rect 42798 205128 42854 205184
rect 43074 206352 43130 206408
rect 42982 205536 43038 205592
rect 48226 204312 48282 204368
rect 42154 190168 42210 190224
rect 41878 187584 41934 187640
rect 41970 187040 42026 187096
rect 42062 186360 42118 186416
rect 42154 185816 42210 185872
rect 42154 184184 42210 184240
rect 41786 183640 41842 183696
rect 41786 182688 41842 182744
rect 62026 316104 62082 316160
rect 59266 311072 59322 311128
rect 56874 224848 56930 224904
rect 59358 298152 59414 298208
rect 59450 285096 59506 285152
rect 62486 938440 62542 938496
rect 62394 596128 62450 596184
rect 62302 278296 62358 278352
rect 62578 684256 62634 684312
rect 62486 278160 62542 278216
rect 102782 999796 102838 999832
rect 102782 999776 102784 999796
rect 102784 999776 102836 999796
rect 102836 999776 102838 999796
rect 104346 999812 104348 999832
rect 104348 999812 104400 999832
rect 104400 999812 104402 999832
rect 104346 999776 104402 999812
rect 102322 999660 102378 999696
rect 102322 999640 102324 999660
rect 102324 999640 102376 999660
rect 102376 999640 102378 999660
rect 101954 999524 102010 999560
rect 101954 999504 101956 999524
rect 101956 999504 102008 999524
rect 102008 999504 102010 999524
rect 103150 999404 103152 999424
rect 103152 999404 103204 999424
rect 103204 999404 103206 999424
rect 96526 996412 96528 996432
rect 96528 996412 96580 996432
rect 96580 996412 96582 996432
rect 96526 996376 96582 996412
rect 96434 995832 96490 995888
rect 96526 995288 96582 995344
rect 103150 999368 103206 999404
rect 107658 997212 107714 997248
rect 107658 997192 107660 997212
rect 107660 997192 107712 997212
rect 107712 997192 107714 997212
rect 115938 997212 115994 997248
rect 115938 997192 115940 997212
rect 115940 997192 115992 997212
rect 115992 997192 115994 997212
rect 101126 996412 101128 996432
rect 101128 996412 101180 996432
rect 101180 996412 101182 996432
rect 101126 996376 101182 996412
rect 100298 996124 100354 996160
rect 100298 996104 100300 996124
rect 100300 996104 100352 996124
rect 100352 996104 100354 996124
rect 100758 996104 100814 996160
rect 101494 996104 101550 996160
rect 108486 996104 108542 996160
rect 108854 996124 108910 996160
rect 108854 996104 108856 996124
rect 108856 996104 108908 996124
rect 108908 996104 108910 996124
rect 110418 995832 110474 995888
rect 100206 995560 100262 995616
rect 104162 995560 104218 995616
rect 104346 995560 104402 995616
rect 99286 995152 99342 995208
rect 100206 993792 100262 993848
rect 104346 993656 104402 993712
rect 110786 995696 110842 995752
rect 110602 995560 110658 995616
rect 142802 995696 142858 995752
rect 137374 995560 137430 995616
rect 144274 997192 144330 997248
rect 133694 995424 133750 995480
rect 141054 995424 141110 995480
rect 160282 1005352 160338 1005388
rect 209226 1005372 209282 1005408
rect 356518 1005388 356520 1005408
rect 356520 1005388 356572 1005408
rect 356572 1005388 356574 1005408
rect 209226 1005352 209228 1005372
rect 209228 1005352 209280 1005372
rect 209280 1005352 209282 1005372
rect 356518 1005352 356574 1005388
rect 361026 1005372 361082 1005408
rect 361026 1005352 361028 1005372
rect 361028 1005352 361080 1005372
rect 361080 1005352 361082 1005372
rect 150898 1004980 150900 1005000
rect 150900 1004980 150952 1005000
rect 150952 1004980 150954 1005000
rect 150898 1004944 150954 1004980
rect 157798 1004964 157854 1005000
rect 157798 1004944 157800 1004964
rect 157800 1004944 157852 1004964
rect 157852 1004944 157854 1004964
rect 156970 1004828 157026 1004864
rect 156970 1004808 156972 1004828
rect 156972 1004808 157024 1004828
rect 157024 1004808 157026 1004828
rect 149702 1004672 149758 1004728
rect 150070 1004672 150126 1004728
rect 148874 996412 148876 996432
rect 148876 996412 148928 996432
rect 148928 996412 148930 996432
rect 148874 996376 148930 996412
rect 151726 996396 151782 996432
rect 151726 996376 151728 996396
rect 151728 996376 151780 996396
rect 151780 996376 151782 996396
rect 154118 996412 154120 996432
rect 154120 996412 154172 996432
rect 154172 996412 154174 996432
rect 154118 996376 154174 996412
rect 153750 996260 153806 996296
rect 153750 996240 153752 996260
rect 153752 996240 153804 996260
rect 153804 996240 153806 996260
rect 150898 996104 150954 996160
rect 151266 996104 151322 996160
rect 152554 996104 152610 996160
rect 152922 996104 152978 996160
rect 153382 996104 153438 996160
rect 146206 995288 146262 995344
rect 154946 1004692 155002 1004728
rect 154946 1004672 154948 1004692
rect 154948 1004672 155000 1004692
rect 155000 1004672 155002 1004692
rect 159454 1004708 159456 1004728
rect 159456 1004708 159508 1004728
rect 159508 1004708 159510 1004728
rect 159454 1004672 159510 1004708
rect 160650 1004692 160706 1004728
rect 160650 1004672 160652 1004692
rect 160652 1004672 160704 1004692
rect 160704 1004672 160706 1004692
rect 155774 999540 155776 999560
rect 155776 999540 155828 999560
rect 155828 999540 155830 999560
rect 155774 999504 155830 999540
rect 159086 999524 159142 999560
rect 159086 999504 159088 999524
rect 159088 999504 159140 999524
rect 159140 999504 159142 999524
rect 158258 999116 158314 999152
rect 158258 999096 158260 999116
rect 158260 999096 158312 999116
rect 158312 999096 158314 999116
rect 156142 997756 156198 997792
rect 156142 997736 156144 997756
rect 156144 997736 156196 997756
rect 156196 997736 156198 997756
rect 154578 996104 154634 996160
rect 156970 996104 157026 996160
rect 157798 996124 157854 996160
rect 157798 996104 157800 996124
rect 157800 996104 157852 996124
rect 157852 996104 157854 996124
rect 159454 996140 159456 996160
rect 159456 996140 159508 996160
rect 159508 996140 159510 996160
rect 159454 996104 159510 996140
rect 162858 997056 162914 997112
rect 168378 995832 168434 995888
rect 162950 995696 163006 995752
rect 162858 995560 162914 995616
rect 195150 997192 195206 997248
rect 187606 995696 187662 995752
rect 201498 1005100 201554 1005136
rect 201498 1005080 201500 1005100
rect 201500 1005080 201552 1005100
rect 201552 1005080 201554 1005100
rect 202326 1005100 202382 1005136
rect 202326 1005080 202328 1005100
rect 202328 1005080 202380 1005100
rect 202380 1005080 202382 1005100
rect 209594 1005116 209596 1005136
rect 209596 1005116 209648 1005136
rect 209648 1005116 209650 1005136
rect 209594 1005080 209650 1005116
rect 210882 1005116 210884 1005136
rect 210884 1005116 210936 1005136
rect 210936 1005116 210938 1005136
rect 210882 1005080 210938 1005116
rect 208398 1004964 208454 1005000
rect 208398 1004944 208400 1004964
rect 208400 1004944 208452 1004964
rect 208452 1004944 208454 1004964
rect 195334 997056 195390 997112
rect 192482 995560 192538 995616
rect 205178 1004692 205234 1004728
rect 205178 1004672 205180 1004692
rect 205180 1004672 205232 1004692
rect 205232 1004672 205234 1004692
rect 205914 1004672 205970 1004728
rect 206374 1004708 206376 1004728
rect 206376 1004708 206428 1004728
rect 206428 1004708 206430 1004728
rect 206374 1004672 206430 1004708
rect 218058 1004672 218114 1004728
rect 205546 999660 205602 999696
rect 205546 999640 205548 999660
rect 205548 999640 205600 999660
rect 205600 999640 205602 999660
rect 203522 999540 203524 999560
rect 203524 999540 203576 999560
rect 203576 999540 203578 999560
rect 203522 999504 203578 999540
rect 203890 999524 203946 999560
rect 203890 999504 203892 999524
rect 203892 999504 203944 999524
rect 203944 999504 203946 999524
rect 202326 999404 202328 999424
rect 202328 999404 202380 999424
rect 202380 999404 202382 999424
rect 202326 999368 202382 999404
rect 204718 999388 204774 999424
rect 204718 999368 204720 999388
rect 204720 999368 204772 999388
rect 204772 999368 204774 999388
rect 202694 999252 202750 999288
rect 202694 999232 202696 999252
rect 202696 999232 202748 999252
rect 202748 999232 202750 999252
rect 204350 999268 204352 999288
rect 204352 999268 204404 999288
rect 204404 999268 204406 999288
rect 204350 999232 204406 999268
rect 203062 999132 203064 999152
rect 203064 999132 203116 999152
rect 203116 999132 203118 999152
rect 203062 999096 203118 999132
rect 210422 997212 210478 997248
rect 210422 997192 210424 997212
rect 210424 997192 210476 997212
rect 210476 997192 210478 997212
rect 215298 997212 215354 997248
rect 215298 997192 215300 997212
rect 215300 997192 215352 997212
rect 215352 997192 215354 997212
rect 208766 996140 208768 996160
rect 208768 996140 208820 996160
rect 208820 996140 208822 996160
rect 208766 996104 208822 996140
rect 209594 996104 209650 996160
rect 211250 996104 211306 996160
rect 211618 996124 211674 996160
rect 211618 996104 211620 996124
rect 211620 996104 211672 996124
rect 211672 996104 211674 996124
rect 191838 993656 191894 993712
rect 207018 995832 207074 995888
rect 207754 995560 207810 995616
rect 216586 995832 216642 995888
rect 259826 1005252 259828 1005272
rect 259828 1005252 259880 1005272
rect 259880 1005252 259882 1005272
rect 259826 1005216 259882 1005252
rect 260194 1005236 260250 1005272
rect 260194 1005216 260196 1005236
rect 260196 1005216 260248 1005236
rect 260248 1005216 260250 1005236
rect 261022 1005100 261078 1005136
rect 261022 1005080 261024 1005100
rect 261024 1005080 261076 1005100
rect 261076 1005080 261078 1005100
rect 263046 1005116 263048 1005136
rect 263048 1005116 263100 1005136
rect 263100 1005116 263102 1005136
rect 263046 1005080 263102 1005116
rect 264334 1005116 264336 1005136
rect 264336 1005116 264388 1005136
rect 264388 1005116 264390 1005136
rect 264334 1005080 264390 1005116
rect 252834 1004980 252836 1005000
rect 252836 1004980 252888 1005000
rect 252888 1004980 252890 1005000
rect 252834 1004944 252890 1004980
rect 253294 1004980 253296 1005000
rect 253296 1004980 253348 1005000
rect 253348 1004980 253350 1005000
rect 253294 1004944 253350 1004980
rect 260654 1004980 260656 1005000
rect 260656 1004980 260708 1005000
rect 260708 1004980 260710 1005000
rect 260654 1004944 260710 1004980
rect 262678 1004964 262734 1005000
rect 262678 1004944 262680 1004964
rect 262680 1004944 262732 1004964
rect 262732 1004944 262734 1004964
rect 264334 1004964 264390 1005000
rect 264334 1004944 264336 1004964
rect 264336 1004944 264388 1004964
rect 264388 1004944 264390 1004964
rect 261850 1004844 261852 1004864
rect 261852 1004844 261904 1004864
rect 261904 1004844 261906 1004864
rect 261850 1004808 261906 1004844
rect 252466 1004672 252522 1004728
rect 252834 1004672 252890 1004728
rect 261482 1004692 261538 1004728
rect 261482 1004672 261484 1004692
rect 261484 1004672 261536 1004692
rect 261536 1004672 261538 1004692
rect 262218 1004708 262220 1004728
rect 262220 1004708 262272 1004728
rect 262272 1004708 262274 1004728
rect 262218 1004672 262274 1004708
rect 263506 1004672 263562 1004728
rect 263874 1004672 263930 1004728
rect 258630 999932 258686 999968
rect 258630 999912 258632 999932
rect 258632 999912 258684 999932
rect 258684 999912 258686 999932
rect 246578 997192 246634 997248
rect 234526 995696 234582 995752
rect 240046 995696 240102 995752
rect 256974 999796 257030 999832
rect 256974 999776 256976 999796
rect 256976 999776 257028 999796
rect 257028 999776 257030 999796
rect 257342 999812 257344 999832
rect 257344 999812 257396 999832
rect 257396 999812 257398 999832
rect 257342 999776 257398 999812
rect 257802 999676 257804 999696
rect 257804 999676 257856 999696
rect 257856 999676 257858 999696
rect 257802 999640 257858 999676
rect 256514 999252 256570 999288
rect 256514 999232 256516 999252
rect 256516 999232 256568 999252
rect 256568 999232 256570 999252
rect 253662 996104 253718 996160
rect 246946 995968 247002 996024
rect 242070 995560 242126 995616
rect 232226 994064 232282 994120
rect 235906 995424 235962 995480
rect 236228 995288 236284 995344
rect 234940 995152 234996 995208
rect 232870 993928 232926 993984
rect 258538 999132 258540 999152
rect 258540 999132 258592 999152
rect 258592 999132 258594 999152
rect 258538 999096 258594 999132
rect 254122 996104 254178 996160
rect 254490 996104 254546 996160
rect 254490 995288 254546 995344
rect 253846 994064 253902 994120
rect 243266 993792 243322 993848
rect 248326 993656 248382 993712
rect 269210 1005080 269266 1005136
rect 267830 1004944 267886 1005000
rect 267738 1004672 267794 1004728
rect 266266 997192 266322 997248
rect 269026 1004808 269082 1004864
rect 360198 1005236 360254 1005272
rect 360198 1005216 360200 1005236
rect 360200 1005216 360252 1005236
rect 360252 1005216 360254 1005236
rect 350262 1004944 350318 1005000
rect 353666 1004944 353722 1005000
rect 358174 1004980 358176 1005000
rect 358176 1004980 358228 1005000
rect 358228 1004980 358230 1005000
rect 358174 1004944 358230 1004980
rect 304078 1004672 304134 1004728
rect 304446 1004672 304502 1004728
rect 315118 1004692 315174 1004728
rect 315118 1004672 315120 1004692
rect 315120 1004672 315172 1004692
rect 315172 1004672 315174 1004692
rect 321466 1004672 321522 1004728
rect 311438 999796 311494 999832
rect 311438 999776 311440 999796
rect 311440 999776 311492 999796
rect 311492 999776 311494 999796
rect 312174 999812 312176 999832
rect 312176 999812 312228 999832
rect 312228 999812 312230 999832
rect 312174 999776 312230 999812
rect 310150 999660 310206 999696
rect 310150 999640 310152 999660
rect 310152 999640 310204 999660
rect 310204 999640 310206 999660
rect 313830 999676 313832 999696
rect 313832 999676 313884 999696
rect 313884 999676 313886 999696
rect 313830 999640 313886 999676
rect 313002 999540 313004 999560
rect 313004 999540 313056 999560
rect 313056 999540 313058 999560
rect 313002 999504 313058 999540
rect 314658 999524 314714 999560
rect 314658 999504 314660 999524
rect 314660 999504 314712 999524
rect 314712 999504 314714 999524
rect 309782 999404 309784 999424
rect 309784 999404 309836 999424
rect 309836 999404 309838 999424
rect 309782 999368 309838 999404
rect 312634 999388 312690 999424
rect 312634 999368 312636 999388
rect 312636 999368 312688 999388
rect 312688 999368 312690 999388
rect 310978 999268 310980 999288
rect 310980 999268 311032 999288
rect 311032 999268 311034 999288
rect 310978 999232 311034 999268
rect 311806 999252 311862 999288
rect 311806 999232 311808 999252
rect 311808 999232 311860 999252
rect 311860 999232 311862 999252
rect 314290 999132 314292 999152
rect 314292 999132 314344 999152
rect 314344 999132 314346 999152
rect 314290 999096 314346 999132
rect 298742 997192 298798 997248
rect 308126 996276 308128 996296
rect 308128 996276 308180 996296
rect 308180 996276 308182 996296
rect 288070 995696 288126 995752
rect 292486 995696 292542 995752
rect 300766 995832 300822 995888
rect 290646 995560 290702 995616
rect 300214 995560 300270 995616
rect 291106 995424 291162 995480
rect 297270 995424 297326 995480
rect 294510 993656 294566 993712
rect 308126 996240 308182 996276
rect 308954 996260 309010 996296
rect 308954 996240 308956 996260
rect 308956 996240 309008 996260
rect 309008 996240 309010 996260
rect 305274 996104 305330 996160
rect 305734 996104 305790 996160
rect 306470 996104 306526 996160
rect 306930 996104 306986 996160
rect 307298 996104 307354 996160
rect 307758 996104 307814 996160
rect 310150 996104 310206 996160
rect 305274 995560 305330 995616
rect 305734 995288 305790 995344
rect 316774 993792 316830 993848
rect 354494 1004672 354550 1004728
rect 354862 1004672 354918 1004728
rect 358542 1004708 358544 1004728
rect 358544 1004708 358596 1004728
rect 358596 1004708 358598 1004728
rect 358542 1004672 358598 1004708
rect 359738 1004692 359794 1004728
rect 359738 1004672 359740 1004692
rect 359740 1004672 359792 1004692
rect 359792 1004672 359794 1004692
rect 360566 1000748 360622 1000784
rect 360566 1000728 360568 1000748
rect 360568 1000728 360620 1000748
rect 360620 1000728 360622 1000748
rect 361394 1000628 361396 1000648
rect 361396 1000628 361448 1000648
rect 361448 1000628 361450 1000648
rect 361394 1000592 361450 1000628
rect 358910 1000492 358912 1000512
rect 358912 1000492 358964 1000512
rect 358964 1000492 358966 1000512
rect 358910 1000456 358966 1000492
rect 357346 999252 357402 999288
rect 357346 999232 357348 999252
rect 357348 999232 357400 999252
rect 357400 999232 357402 999252
rect 357714 999132 357716 999152
rect 357716 999132 357768 999152
rect 357768 999132 357770 999152
rect 357714 999096 357770 999132
rect 425150 1005388 425152 1005408
rect 425152 1005388 425204 1005408
rect 425204 1005388 425206 1005408
rect 425150 1005352 425206 1005388
rect 428370 1005372 428426 1005408
rect 428370 1005352 428372 1005372
rect 428372 1005352 428424 1005372
rect 428424 1005352 428426 1005372
rect 427542 1005116 427544 1005136
rect 427544 1005116 427596 1005136
rect 427596 1005116 427598 1005136
rect 427542 1005080 427598 1005116
rect 428830 1005100 428886 1005136
rect 428830 1005080 428832 1005100
rect 428832 1005080 428884 1005100
rect 428884 1005080 428886 1005100
rect 363418 997212 363474 997248
rect 363418 997192 363420 997212
rect 363420 997192 363472 997212
rect 363472 997192 363474 997212
rect 367098 997212 367154 997248
rect 367098 997192 367100 997212
rect 367100 997192 367152 997212
rect 367152 997192 367154 997212
rect 365442 996260 365498 996296
rect 365442 996240 365444 996260
rect 365444 996240 365496 996260
rect 365496 996240 365498 996260
rect 362590 996104 362646 996160
rect 364246 996140 364248 996160
rect 364248 996140 364300 996160
rect 364300 996140 364302 996160
rect 364246 996104 364302 996140
rect 364706 996124 364762 996160
rect 364706 996104 364708 996124
rect 364708 996104 364760 996124
rect 364760 996104 364762 996124
rect 365074 996104 365130 996160
rect 353666 995832 353722 995888
rect 367098 995832 367154 995888
rect 359186 995560 359242 995616
rect 366178 993656 366234 993712
rect 367190 995696 367246 995752
rect 367466 995560 367522 995616
rect 371514 996104 371570 996160
rect 381726 996376 381782 996432
rect 425518 1004964 425574 1005000
rect 425518 1004944 425520 1004964
rect 425520 1004944 425572 1004964
rect 425572 1004944 425574 1004964
rect 426806 1004980 426808 1005000
rect 426808 1004980 426860 1005000
rect 426860 1004980 426862 1005000
rect 426806 1004944 426862 1004980
rect 423494 1004828 423550 1004864
rect 423494 1004808 423496 1004828
rect 423496 1004808 423548 1004828
rect 423548 1004808 423550 1004828
rect 427174 1004844 427176 1004864
rect 427176 1004844 427228 1004864
rect 427228 1004844 427230 1004864
rect 427174 1004808 427230 1004844
rect 422298 1004692 422354 1004728
rect 422298 1004672 422300 1004692
rect 422300 1004672 422352 1004692
rect 422352 1004672 422354 1004692
rect 422666 1004672 422722 1004728
rect 424690 1004708 424692 1004728
rect 424692 1004708 424744 1004728
rect 424744 1004708 424746 1004728
rect 424690 1004672 424746 1004708
rect 399942 997192 399998 997248
rect 388166 995696 388222 995752
rect 378138 993792 378194 993848
rect 374458 993656 374514 993712
rect 396998 993792 397054 993848
rect 395158 993656 395214 993712
rect 428002 1000612 428058 1000648
rect 428002 1000592 428004 1000612
rect 428004 1000592 428056 1000612
rect 428056 1000592 428058 1000612
rect 426346 1000492 426348 1000512
rect 426348 1000492 426400 1000512
rect 426400 1000492 426402 1000512
rect 426346 1000456 426402 1000492
rect 430854 999796 430910 999832
rect 430854 999776 430856 999796
rect 430856 999776 430908 999796
rect 430908 999776 430910 999796
rect 429198 999660 429254 999696
rect 429198 999640 429200 999660
rect 429200 999640 429252 999660
rect 429252 999640 429254 999660
rect 431682 999676 431684 999696
rect 431684 999676 431736 999696
rect 431736 999676 431738 999696
rect 431682 999640 431738 999676
rect 430026 999540 430028 999560
rect 430028 999540 430080 999560
rect 430080 999540 430082 999560
rect 430026 999504 430082 999540
rect 431222 999524 431278 999560
rect 431222 999504 431224 999524
rect 431224 999504 431276 999524
rect 431276 999504 431278 999524
rect 429658 999404 429660 999424
rect 429660 999404 429712 999424
rect 429712 999404 429714 999424
rect 429658 999368 429714 999404
rect 432510 999388 432566 999424
rect 432510 999368 432512 999388
rect 432512 999368 432564 999388
rect 432564 999368 432566 999388
rect 432050 999252 432106 999288
rect 432050 999232 432052 999252
rect 432052 999232 432104 999252
rect 432104 999232 432106 999252
rect 432878 999268 432880 999288
rect 432880 999268 432932 999288
rect 432932 999268 432934 999288
rect 432878 999232 432934 999268
rect 430394 999132 430396 999152
rect 430396 999132 430448 999152
rect 430448 999132 430450 999152
rect 430394 999096 430450 999132
rect 437754 999096 437810 999152
rect 438122 997056 438178 997112
rect 447138 995696 447194 995752
rect 504546 1005660 504548 1005680
rect 504548 1005660 504600 1005680
rect 504600 1005660 504602 1005680
rect 504546 1005624 504602 1005660
rect 505006 1005644 505062 1005680
rect 505006 1005624 505008 1005644
rect 505008 1005624 505060 1005644
rect 505060 1005624 505062 1005644
rect 502982 1005508 503038 1005544
rect 502982 1005488 502984 1005508
rect 502984 1005488 503036 1005508
rect 503036 1005488 503038 1005508
rect 505374 1005524 505376 1005544
rect 505376 1005524 505428 1005544
rect 505428 1005524 505430 1005544
rect 505374 1005488 505430 1005524
rect 461030 996376 461086 996432
rect 447322 993656 447378 993712
rect 505834 1005372 505890 1005408
rect 505834 1005352 505836 1005372
rect 505836 1005352 505888 1005372
rect 505888 1005352 505890 1005372
rect 502522 1005100 502578 1005136
rect 502522 1005080 502524 1005100
rect 502524 1005080 502576 1005100
rect 502576 1005080 502578 1005100
rect 504178 1004980 504180 1005000
rect 504180 1004980 504232 1005000
rect 504232 1004980 504234 1005000
rect 504178 1004944 504234 1004980
rect 499302 1004692 499358 1004728
rect 499302 1004672 499304 1004692
rect 499304 1004672 499356 1004692
rect 499356 1004672 499358 1004692
rect 499670 1004672 499726 1004728
rect 501694 1004708 501696 1004728
rect 501696 1004708 501748 1004728
rect 501748 1004708 501750 1004728
rect 501694 1004672 501750 1004708
rect 502154 1004692 502210 1004728
rect 502154 1004672 502156 1004692
rect 502156 1004672 502208 1004692
rect 502208 1004672 502210 1004692
rect 469402 995288 469458 995344
rect 489458 997056 489514 997112
rect 481454 995696 481510 995752
rect 471702 995560 471758 995616
rect 477682 995560 477738 995616
rect 476486 995424 476542 995480
rect 481086 995288 481142 995344
rect 478602 993656 478658 993712
rect 503350 999948 503352 999968
rect 503352 999948 503404 999968
rect 503404 999948 503406 999968
rect 503350 999912 503406 999948
rect 508686 999796 508742 999832
rect 508686 999776 508688 999796
rect 508688 999776 508740 999796
rect 508740 999776 508742 999796
rect 506202 999676 506204 999696
rect 506204 999676 506256 999696
rect 506256 999676 506258 999696
rect 506202 999640 506258 999676
rect 507030 999660 507086 999696
rect 507030 999640 507032 999660
rect 507032 999640 507084 999660
rect 507084 999640 507086 999660
rect 507858 999524 507914 999560
rect 507858 999504 507860 999524
rect 507860 999504 507912 999524
rect 507912 999504 507914 999524
rect 508226 999540 508228 999560
rect 508228 999540 508280 999560
rect 508280 999540 508282 999560
rect 508226 999504 508282 999540
rect 500498 999388 500554 999424
rect 500498 999368 500500 999388
rect 500500 999368 500552 999388
rect 500552 999368 500554 999388
rect 506570 999404 506572 999424
rect 506572 999404 506624 999424
rect 506624 999404 506626 999424
rect 506570 999368 506626 999404
rect 509054 999388 509110 999424
rect 509054 999368 509056 999388
rect 509056 999368 509108 999388
rect 509108 999368 509110 999388
rect 500866 999252 500922 999288
rect 500866 999232 500868 999252
rect 500868 999232 500920 999252
rect 500920 999232 500922 999252
rect 507398 999252 507454 999288
rect 507398 999232 507400 999252
rect 507400 999232 507452 999252
rect 507452 999232 507454 999252
rect 501326 997756 501382 997792
rect 501326 997736 501328 997756
rect 501328 997736 501380 997756
rect 501380 997736 501382 997756
rect 503626 995560 503682 995616
rect 516046 999948 516048 999968
rect 516048 999948 516100 999968
rect 516100 999948 516102 999968
rect 516046 999912 516102 999948
rect 509514 999268 509516 999288
rect 509516 999268 509568 999288
rect 509568 999268 509570 999288
rect 509514 999232 509570 999268
rect 509882 999132 509884 999152
rect 509884 999132 509936 999152
rect 509936 999132 509938 999152
rect 509882 999096 509938 999132
rect 515034 999096 515090 999152
rect 519082 999096 519138 999152
rect 519542 996376 519598 996432
rect 521566 995560 521622 995616
rect 521290 995288 521346 995344
rect 546314 1004944 546370 1005000
rect 549442 1004944 549498 1005000
rect 552754 1004964 552810 1005000
rect 552754 1004944 552756 1004964
rect 552756 1004944 552808 1004964
rect 552808 1004944 552810 1004964
rect 523774 999096 523830 999152
rect 523774 996512 523830 996568
rect 524050 999912 524106 999968
rect 523866 995696 523922 995752
rect 527914 995696 527970 995752
rect 532238 995696 532294 995752
rect 530122 995560 530178 995616
rect 526166 995424 526222 995480
rect 533986 995288 534042 995344
rect 521658 995152 521714 995208
rect 537390 995288 537446 995344
rect 553122 1004828 553178 1004864
rect 553122 1004808 553124 1004828
rect 553124 1004808 553176 1004828
rect 553176 1004808 553178 1004828
rect 550270 1004672 550326 1004728
rect 550638 1004672 550694 1004728
rect 551926 1004708 551928 1004728
rect 551928 1004708 551980 1004728
rect 551980 1004708 551982 1004728
rect 551926 1004672 551982 1004708
rect 554318 1004692 554374 1004728
rect 554318 1004672 554320 1004692
rect 554320 1004672 554372 1004692
rect 554372 1004672 554374 1004692
rect 553950 1003892 553952 1003912
rect 553952 1003892 554004 1003912
rect 554004 1003892 554006 1003912
rect 553950 1003856 554006 1003892
rect 555514 1003332 555570 1003368
rect 555514 1003312 555516 1003332
rect 555516 1003312 555568 1003332
rect 555568 1003312 555570 1003332
rect 554778 1003212 554780 1003232
rect 554780 1003212 554832 1003232
rect 554832 1003212 554834 1003232
rect 554778 1003176 554834 1003212
rect 561310 1004692 561366 1004728
rect 561310 1004672 561312 1004692
rect 561312 1004672 561364 1004692
rect 561364 1004672 561366 1004692
rect 567290 1004672 567346 1004728
rect 560850 999796 560906 999832
rect 560850 999776 560852 999796
rect 560852 999776 560904 999796
rect 560904 999776 560906 999796
rect 560482 999660 560538 999696
rect 560482 999640 560484 999660
rect 560484 999640 560536 999660
rect 560536 999640 560538 999660
rect 552294 999132 552296 999152
rect 552296 999132 552348 999152
rect 552348 999132 552350 999152
rect 552294 999096 552350 999132
rect 553490 997756 553546 997792
rect 553490 997736 553492 997756
rect 553492 997736 553544 997756
rect 553544 997736 553546 997756
rect 556342 997636 556344 997656
rect 556344 997636 556396 997656
rect 556396 997636 556398 997656
rect 556342 997600 556398 997636
rect 557170 997484 557226 997520
rect 557170 997464 557172 997484
rect 557172 997464 557224 997484
rect 557224 997464 557226 997484
rect 558458 996124 558514 996160
rect 558458 996104 558460 996124
rect 558460 996104 558512 996124
rect 558512 996104 558514 996124
rect 559286 996140 559288 996160
rect 559288 996140 559340 996160
rect 559340 996140 559342 996160
rect 559286 996104 559342 996140
rect 549442 995832 549498 995888
rect 557722 995696 557778 995752
rect 558550 995696 558606 995752
rect 564346 995696 564402 995752
rect 555054 995560 555110 995616
rect 561678 995560 561734 995616
rect 561494 995424 561550 995480
rect 561310 995288 561366 995344
rect 561310 993792 561366 993848
rect 561494 993656 561550 993712
rect 561678 985632 561734 985688
rect 564714 995832 564770 995888
rect 564438 985768 564494 985824
rect 568670 994200 568726 994256
rect 568578 994064 568634 994120
rect 570142 993928 570198 993984
rect 629666 993792 629722 993848
rect 634818 994200 634874 994256
rect 638544 995152 638600 995208
rect 637026 994064 637082 994120
rect 635186 993928 635242 993984
rect 638866 993656 638922 993712
rect 641166 995152 641222 995208
rect 62854 814136 62910 814192
rect 62762 427896 62818 427952
rect 62670 278024 62726 278080
rect 63222 729816 63278 729872
rect 62854 277888 62910 277944
rect 63038 277752 63094 277808
rect 63314 383832 63370 383888
rect 63222 277616 63278 277672
rect 70582 271768 70638 271824
rect 69386 269048 69442 269104
rect 76470 271904 76526 271960
rect 78862 269320 78918 269376
rect 83554 272040 83610 272096
rect 85946 272176 86002 272232
rect 87142 269728 87198 269784
rect 84750 269456 84806 269512
rect 77666 269184 77722 269240
rect 91834 272312 91890 272368
rect 90638 269592 90694 269648
rect 97722 272720 97778 272776
rect 100114 272584 100170 272640
rect 98918 272448 98974 272504
rect 101310 270000 101366 270056
rect 96618 269864 96674 269920
rect 107198 272992 107254 273048
rect 106002 272856 106058 272912
rect 108394 270272 108450 270328
rect 103702 270136 103758 270192
rect 111982 273128 112038 273184
rect 115478 271632 115534 271688
rect 122562 271496 122618 271552
rect 121366 270408 121422 270464
rect 128542 268912 128598 268968
rect 127346 268776 127402 268832
rect 142710 268640 142766 268696
rect 153290 268504 153346 268560
rect 184938 268368 184994 268424
rect 194138 271768 194194 271824
rect 194506 271788 194562 271824
rect 194506 271768 194508 271788
rect 194508 271768 194560 271788
rect 194560 271768 194562 271788
rect 193678 269048 193734 269104
rect 196346 271904 196402 271960
rect 196806 269184 196862 269240
rect 199106 272040 199162 272096
rect 199934 272176 199990 272232
rect 199014 269456 199070 269512
rect 197726 269320 197782 269376
rect 200394 269728 200450 269784
rect 201314 272720 201370 272776
rect 202142 272312 202198 272368
rect 201682 269592 201738 269648
rect 203430 272992 203486 273048
rect 203062 268368 203118 268424
rect 203430 268096 203486 268152
rect 204810 272448 204866 272504
rect 204350 269864 204406 269920
rect 205730 272584 205786 272640
rect 205270 270000 205326 270056
rect 207478 272856 207534 272912
rect 207018 270136 207074 270192
rect 208490 271768 208546 271824
rect 207938 270272 207994 270328
rect 209226 273128 209282 273184
rect 208398 268096 208454 268152
rect 210606 271632 210662 271688
rect 213274 271496 213330 271552
rect 213734 270408 213790 270464
rect 215482 268776 215538 268832
rect 216402 268912 216458 268968
rect 221738 268640 221794 268696
rect 225786 268504 225842 268560
rect 353942 268232 353998 268288
rect 356610 268368 356666 268424
rect 358910 268640 358966 268696
rect 359370 268504 359426 268560
rect 362038 268776 362094 268832
rect 363326 271360 363382 271416
rect 364246 268912 364302 268968
rect 365534 271632 365590 271688
rect 365994 271496 366050 271552
rect 366914 270408 366970 270464
rect 368662 273128 368718 273184
rect 369582 270272 369638 270328
rect 371238 272992 371294 273048
rect 371330 272856 371386 272912
rect 372250 270136 372306 270192
rect 373998 272720 374054 272776
rect 378046 270000 378102 270056
rect 379334 272584 379390 272640
rect 383382 269864 383438 269920
rect 385130 266056 385186 266112
rect 386970 267552 387026 267608
rect 386510 266192 386566 266248
rect 388258 275848 388314 275904
rect 387798 267688 387854 267744
rect 389638 267416 389694 267472
rect 391294 275712 391350 275768
rect 390466 267280 390522 267336
rect 391386 269728 391442 269784
rect 392766 272448 392822 272504
rect 391846 267144 391902 267200
rect 393134 267008 393190 267064
rect 393594 275576 393650 275632
rect 394514 266872 394570 266928
rect 396262 275440 396318 275496
rect 395802 266736 395858 266792
rect 397182 266600 397238 266656
rect 398930 275304 398986 275360
rect 398102 272312 398158 272368
rect 398470 266464 398526 266520
rect 399850 266328 399906 266384
rect 401690 275168 401746 275224
rect 402702 274896 402758 274952
rect 402058 269592 402114 269648
rect 403438 272176 403494 272232
rect 404266 275032 404322 275088
rect 405370 274760 405426 274816
rect 404726 269456 404782 269512
rect 405462 265920 405518 265976
rect 406934 274624 406990 274680
rect 408222 274488 408278 274544
rect 407394 269320 407450 269376
rect 408314 265784 408370 265840
rect 408774 272040 408830 272096
rect 410890 271904 410946 271960
rect 409602 269184 409658 269240
rect 410062 269048 410118 269104
rect 411074 271768 411130 271824
rect 465906 265920 465962 265976
rect 459466 265784 459522 265840
rect 494978 268232 495034 268288
rect 502062 268368 502118 268424
rect 507950 268640 508006 268696
rect 509146 268504 509202 268560
rect 516230 268776 516286 268832
rect 519818 271360 519874 271416
rect 522210 268912 522266 268968
rect 525706 271632 525762 271688
rect 526902 271496 526958 271552
rect 529294 270408 529350 270464
rect 533986 273128 534042 273184
rect 536378 270272 536434 270328
rect 539874 272992 539930 273048
rect 541070 272856 541126 272912
rect 543462 270136 543518 270192
rect 548154 272720 548210 272776
rect 558826 270000 558882 270056
rect 562414 272584 562470 272640
rect 572994 269864 573050 269920
rect 586058 275848 586114 275904
rect 584862 267688 584918 267744
rect 582470 267552 582526 267608
rect 589554 267416 589610 267472
rect 593142 275712 593198 275768
rect 594338 269728 594394 269784
rect 591946 267280 592002 267336
rect 595442 267144 595498 267200
rect 597834 272448 597890 272504
rect 600226 275576 600282 275632
rect 599030 267008 599086 267064
rect 602526 266872 602582 266928
rect 607310 275440 607366 275496
rect 606114 266736 606170 266792
rect 612002 272312 612058 272368
rect 609702 266600 609758 266656
rect 614394 275304 614450 275360
rect 613198 266464 613254 266520
rect 621478 275168 621534 275224
rect 623870 274896 623926 274952
rect 628562 275032 628618 275088
rect 626170 272176 626226 272232
rect 622674 269592 622730 269648
rect 630954 274760 631010 274816
rect 635646 274624 635702 274680
rect 629758 269456 629814 269512
rect 638038 274488 638094 274544
rect 640430 272040 640486 272096
rect 636842 269320 636898 269376
rect 642730 269184 642786 269240
rect 645122 271904 645178 271960
rect 646318 271768 646374 271824
rect 643926 269048 643982 269104
rect 616786 266328 616842 266384
rect 581274 266192 581330 266248
rect 577778 266056 577834 266112
rect 418066 262656 418122 262712
rect 417790 260208 417846 260264
rect 184938 259936 184994 259992
rect 418342 257896 418398 257952
rect 416778 255448 416834 255504
rect 416778 253136 416834 253192
rect 184938 251912 184994 251968
rect 416778 250688 416834 250744
rect 418066 248240 418122 248296
rect 184938 244024 184994 244080
rect 106186 236952 106242 237008
rect 89626 236816 89682 236872
rect 81346 236408 81402 236464
rect 73066 236272 73122 236328
rect 62026 235864 62082 235920
rect 61106 222128 61162 222184
rect 63406 224984 63462 225040
rect 66166 222264 66222 222320
rect 70398 225120 70454 225176
rect 67822 222400 67878 222456
rect 72882 222672 72938 222728
rect 75826 236136 75882 236192
rect 74446 222536 74502 222592
rect 78586 236000 78642 236056
rect 77114 225256 77170 225312
rect 80426 225392 80482 225448
rect 79598 222808 79654 222864
rect 83830 225528 83886 225584
rect 88890 225800 88946 225856
rect 97906 236680 97962 236736
rect 95146 236544 95202 236600
rect 92202 225664 92258 225720
rect 96434 222944 96490 223000
rect 102046 226072 102102 226128
rect 98918 225936 98974 225992
rect 104806 223080 104862 223136
rect 111614 223216 111670 223272
rect 121366 223352 121422 223408
rect 153106 237088 153162 237144
rect 193402 224848 193458 224904
rect 194414 236272 194470 236328
rect 194782 235864 194838 235920
rect 196254 224984 196310 225040
rect 196162 222264 196218 222320
rect 196990 236816 197046 236872
rect 197634 236136 197690 236192
rect 196530 222128 196586 222184
rect 200486 236408 200542 236464
rect 199106 225120 199162 225176
rect 198738 222400 198794 222456
rect 201682 222672 201738 222728
rect 202970 236000 203026 236056
rect 202050 225256 202106 225312
rect 201866 222536 201922 222592
rect 203430 225392 203486 225448
rect 204350 222808 204406 222864
rect 204810 225528 204866 225584
rect 205822 236680 205878 236736
rect 206190 236544 206246 236600
rect 207570 236952 207626 237008
rect 206650 225800 206706 225856
rect 208030 225664 208086 225720
rect 210054 237088 210110 237144
rect 210882 225936 210938 225992
rect 211250 222944 211306 223000
rect 212814 226072 212870 226128
rect 214470 223080 214526 223136
rect 217690 235864 217746 235920
rect 217322 223216 217378 223272
rect 221554 223352 221610 223408
rect 226246 236000 226302 236056
rect 229006 236136 229062 236192
rect 234526 236272 234582 236328
rect 238758 236544 238814 236600
rect 240046 236408 240102 236464
rect 249890 236952 249946 237008
rect 249706 236680 249762 236736
rect 250166 237224 250222 237280
rect 252558 236816 252614 236872
rect 262862 235864 262918 235920
rect 265714 237224 265770 237280
rect 266082 236000 266138 236056
rect 267094 236136 267150 236192
rect 268566 236952 268622 237008
rect 268198 236544 268254 236600
rect 269946 236680 270002 236736
rect 268934 236272 268990 236328
rect 271418 236816 271474 236872
rect 271786 236408 271842 236464
rect 328090 222808 328146 222864
rect 330758 222672 330814 222728
rect 331034 223080 331090 223136
rect 331126 222944 331182 223000
rect 330942 222536 330998 222592
rect 333610 222400 333666 222456
rect 333702 222264 333758 222320
rect 336186 221992 336242 222048
rect 339314 223488 339370 223544
rect 341614 222128 341670 222184
rect 360934 226072 360990 226128
rect 364062 225936 364118 225992
rect 363694 225664 363750 225720
rect 366546 228792 366602 228848
rect 368018 228656 368074 228712
rect 367006 225800 367062 225856
rect 366362 225528 366418 225584
rect 369122 225392 369178 225448
rect 369766 228384 369822 228440
rect 371238 228520 371294 228576
rect 370870 228112 370926 228168
rect 369398 227976 369454 228032
rect 371974 225256 372030 225312
rect 369214 225120 369270 225176
rect 372618 228248 372674 228304
rect 374090 227840 374146 227896
rect 373722 227704 373778 227760
rect 372250 227568 372306 227624
rect 372066 224984 372122 225040
rect 375838 237088 375894 237144
rect 374734 224848 374790 224904
rect 374642 223352 374698 223408
rect 374182 222808 374238 222864
rect 375378 222672 375434 222728
rect 378322 236952 378378 237008
rect 378690 236816 378746 236872
rect 377586 223216 377642 223272
rect 376758 223080 376814 223136
rect 377954 223080 378010 223136
rect 377586 222944 377642 223000
rect 381174 236680 381230 236736
rect 381542 236408 381598 236464
rect 380714 222944 380770 223000
rect 380438 222808 380494 222864
rect 381082 222536 381138 222592
rect 383658 236544 383714 236600
rect 385866 236272 385922 236328
rect 382922 222536 382978 222592
rect 384302 222400 384358 222456
rect 387982 236136 388038 236192
rect 386234 222672 386290 222728
rect 387706 222264 387762 222320
rect 389086 236000 389142 236056
rect 388994 222400 389050 222456
rect 390190 221992 390246 222048
rect 391202 235864 391258 235920
rect 391846 222264 391902 222320
rect 396906 223488 396962 223544
rect 400402 222128 400458 222184
rect 411166 222128 411222 222184
rect 418434 245928 418490 245984
rect 418158 243480 418214 243536
rect 418526 241168 418582 241224
rect 486422 237088 486478 237144
rect 451554 226072 451610 226128
rect 454958 225936 455014 225992
rect 456614 225664 456670 225720
rect 460018 225800 460074 225856
rect 463698 225528 463754 225584
rect 465078 228792 465134 228848
rect 466734 225392 466790 225448
rect 468390 228656 468446 228712
rect 469218 228384 469274 228440
rect 470138 225120 470194 225176
rect 472622 228520 472678 228576
rect 471978 227976 472034 228032
rect 473450 225256 473506 225312
rect 476026 228248 476082 228304
rect 475106 228112 475162 228168
rect 476854 224984 476910 225040
rect 479338 227840 479394 227896
rect 478510 227568 478566 227624
rect 480258 224848 480314 224904
rect 481914 227704 481970 227760
rect 483846 223352 483902 223408
rect 492310 236952 492366 237008
rect 489458 223216 489514 223272
rect 488630 223080 488686 223136
rect 488630 221176 488686 221232
rect 492586 236816 492642 236872
rect 497002 236680 497058 236736
rect 494058 222808 494114 222864
rect 494058 221040 494114 221096
rect 492678 220904 492734 220960
rect 495346 222944 495402 223000
rect 496450 221040 496506 221096
rect 502706 236544 502762 236600
rect 499946 236408 500002 236464
rect 502614 222536 502670 222592
rect 502614 221448 502670 221504
rect 507858 236272 507914 236328
rect 507122 222672 507178 222728
rect 507122 221312 507178 221368
rect 513746 236136 513802 236192
rect 510618 222400 510674 222456
rect 510618 221584 510674 221640
rect 517426 236000 517482 236056
rect 512458 221584 512514 221640
rect 522946 235864 523002 235920
rect 517426 222264 517482 222320
rect 517886 222264 517942 222320
rect 519726 222400 519782 222456
rect 522946 221856 523002 221912
rect 528466 221992 528522 222048
rect 528650 222264 528706 222320
rect 527914 221720 527970 221776
rect 528466 221720 528522 221776
rect 528650 221720 528706 221776
rect 569314 222128 569370 222184
rect 569866 222128 569922 222184
rect 572626 222536 572682 222592
rect 574374 222536 574430 222592
rect 573546 222128 573602 222184
rect 579710 216144 579766 216200
rect 582286 214648 582342 214704
rect 580262 213152 580318 213208
rect 581642 211656 581698 211712
rect 580538 210160 580594 210216
rect 581458 208664 581514 208720
rect 582286 207068 582288 207088
rect 582288 207068 582340 207088
rect 582340 207068 582342 207088
rect 582286 207032 582342 207068
rect 582286 205536 582342 205592
rect 599766 209480 599822 209536
rect 628010 221992 628066 222048
rect 627090 221856 627146 221912
rect 626170 221720 626226 221776
rect 625250 221584 625306 221640
rect 623410 221448 623466 221504
rect 621478 221176 621534 221232
rect 624330 221312 624386 221368
rect 637394 221040 637450 221096
rect 636934 220904 636990 220960
rect 654690 922664 654746 922720
rect 654874 909472 654930 909528
rect 654690 896144 654746 896200
rect 655150 882816 655206 882872
rect 655242 856296 655298 856352
rect 654874 842968 654930 843024
rect 655058 816448 655114 816504
rect 655058 789928 655114 789984
rect 654690 763272 654746 763328
rect 654690 750080 654746 750136
rect 654138 736752 654194 736808
rect 654874 696904 654930 696960
rect 654138 683576 654194 683632
rect 654874 643728 654930 643784
rect 654138 630536 654194 630592
rect 654598 617208 654654 617264
rect 654322 603880 654378 603936
rect 654506 577360 654562 577416
rect 654322 564032 654378 564088
rect 655058 550840 655114 550896
rect 654690 537512 654746 537568
rect 654138 524184 654194 524240
rect 654782 510992 654838 511048
rect 655058 484336 655114 484392
rect 654874 471144 654930 471200
rect 654138 457816 654194 457872
rect 654874 431296 654930 431352
rect 655058 417968 655114 418024
rect 654874 404640 654930 404696
rect 654138 391448 654194 391504
rect 654874 351600 654930 351656
rect 654322 338272 654378 338328
rect 654322 324944 654378 325000
rect 654138 311752 654194 311808
rect 655518 975840 655574 975896
rect 655702 962512 655758 962568
rect 655794 949320 655850 949376
rect 655610 936128 655666 936184
rect 656806 869644 656862 869680
rect 656806 869624 656808 869644
rect 656808 869624 656860 869644
rect 656860 869624 656862 869644
rect 655518 829776 655574 829832
rect 656162 803276 656218 803312
rect 656162 803256 656164 803276
rect 656164 803256 656216 803276
rect 656216 803256 656218 803276
rect 655518 776600 655574 776656
rect 655518 723424 655574 723480
rect 655978 710232 656034 710288
rect 655518 670384 655574 670440
rect 656806 657076 656862 657112
rect 656806 657056 656808 657076
rect 656808 657056 656860 657076
rect 656860 657056 656862 657076
rect 656806 590708 656862 590744
rect 656806 590688 656808 590708
rect 656808 590688 656860 590708
rect 656860 590688 656862 590708
rect 656806 497684 656862 497720
rect 656806 497664 656808 497684
rect 656808 497664 656860 497684
rect 656860 497664 656862 497684
rect 656806 444508 656862 444544
rect 656806 444488 656808 444508
rect 656808 444488 656860 444508
rect 656860 444488 656862 444508
rect 656806 378156 656808 378176
rect 656808 378156 656860 378176
rect 656860 378156 656862 378176
rect 656806 378120 656862 378156
rect 656806 364792 656862 364848
rect 656806 298444 656862 298480
rect 656806 298424 656808 298444
rect 656808 298424 656860 298444
rect 656860 298424 656862 298444
rect 655702 285232 655758 285288
rect 658186 262384 658242 262440
rect 599950 208528 600006 208584
rect 599858 207440 599914 207496
rect 600042 206488 600098 206544
rect 599122 205400 599178 205456
rect 600962 204448 601018 204504
rect 581826 204040 581882 204096
rect 581090 202544 581146 202600
rect 601146 203360 601202 203416
rect 599950 202408 600006 202464
rect 599030 201320 599086 201376
rect 581090 201048 581146 201104
rect 599950 200368 600006 200424
rect 582286 199552 582342 199608
rect 599950 199280 600006 199336
rect 599122 198328 599178 198384
rect 581274 197920 581330 197976
rect 599306 197240 599362 197296
rect 580814 196424 580870 196480
rect 599950 196288 600006 196344
rect 599950 195200 600006 195256
rect 582286 194928 582342 194984
rect 599122 194248 599178 194304
rect 582194 193432 582250 193488
rect 599858 193160 599914 193216
rect 582286 191936 582342 191992
rect 599950 192208 600006 192264
rect 599858 191120 599914 191176
rect 581274 190440 581330 190496
rect 600962 190168 601018 190224
rect 579710 188808 579766 188864
rect 601606 189080 601662 189136
rect 601514 188128 601570 188184
rect 582286 187312 582342 187368
rect 599950 187040 600006 187096
rect 582194 185816 582250 185872
rect 599858 185000 599914 185056
rect 580906 184320 580962 184376
rect 599766 184048 599822 184104
rect 580262 182824 580318 182880
rect 580538 181328 580594 181384
rect 581826 179696 581882 179752
rect 600042 186088 600098 186144
rect 599950 182960 600006 183016
rect 599858 182008 599914 182064
rect 599674 178880 599730 178936
rect 581090 178200 581146 178256
rect 598938 176840 598994 176896
rect 580722 176704 580778 176760
rect 579710 172216 579766 172272
rect 580078 169088 580134 169144
rect 580170 166096 580226 166152
rect 579894 161472 579950 161528
rect 579710 158480 579766 158536
rect 580906 170584 580962 170640
rect 581458 175208 581514 175264
rect 582286 173748 582288 173768
rect 582288 173748 582340 173768
rect 582340 173748 582342 173768
rect 582286 173712 582342 173748
rect 581090 167592 581146 167648
rect 580814 164600 580870 164656
rect 580262 155488 580318 155544
rect 580078 152360 580134 152416
rect 579710 122032 579766 122088
rect 580722 143248 580778 143304
rect 580630 138760 580686 138816
rect 579802 119040 579858 119096
rect 579894 112920 579950 112976
rect 580078 108432 580134 108488
rect 581090 147872 581146 147928
rect 581826 163104 581882 163160
rect 581550 150864 581606 150920
rect 581642 149368 581698 149424
rect 581182 144880 581238 144936
rect 580998 141752 581054 141808
rect 580906 137264 580962 137320
rect 580814 134136 580870 134192
rect 580170 106800 580226 106856
rect 579986 105304 580042 105360
rect 580262 103808 580318 103864
rect 580446 100816 580502 100872
rect 580538 99320 580594 99376
rect 580354 97688 580410 97744
rect 580722 96192 580778 96248
rect 580998 111424 581054 111480
rect 581274 123528 581330 123584
rect 581458 125024 581514 125080
rect 581918 156984 581974 157040
rect 581734 146376 581790 146432
rect 581642 126656 581698 126712
rect 599766 177928 599822 177984
rect 600134 180920 600190 180976
rect 600042 179968 600098 180024
rect 599950 174800 600006 174856
rect 600226 175888 600282 175944
rect 599858 172760 599914 172816
rect 599950 171808 600006 171864
rect 598938 170720 598994 170776
rect 599950 169768 600006 169824
rect 599490 168680 599546 168736
rect 601422 173848 601478 173904
rect 599858 167728 599914 167784
rect 600042 166640 600098 166696
rect 582194 159976 582250 160032
rect 582010 140256 582066 140312
rect 599950 165688 600006 165744
rect 599858 164600 599914 164656
rect 599950 163648 600006 163704
rect 600042 162560 600098 162616
rect 599858 161608 599914 161664
rect 599950 160520 600006 160576
rect 600042 159568 600098 159624
rect 599858 158480 599914 158536
rect 599950 157548 600006 157584
rect 599950 157528 599952 157548
rect 599952 157528 600004 157548
rect 600004 157528 600006 157548
rect 599858 156440 599914 156496
rect 599950 155488 600006 155544
rect 600042 154400 600098 154456
rect 582286 153992 582342 154048
rect 599858 153448 599914 153504
rect 599950 152360 600006 152416
rect 582102 135768 582158 135824
rect 598938 151408 598994 151464
rect 599858 150320 599914 150376
rect 599950 149368 600006 149424
rect 599858 148280 599914 148336
rect 599950 147328 600006 147384
rect 582194 132640 582250 132696
rect 581918 131144 581974 131200
rect 581826 129648 581882 129704
rect 599582 146240 599638 146296
rect 599950 145288 600006 145344
rect 599674 144200 599730 144256
rect 599858 143248 599914 143304
rect 599306 141208 599362 141264
rect 599950 142160 600006 142216
rect 600042 140120 600098 140176
rect 599858 139168 599914 139224
rect 599950 138116 599952 138136
rect 599952 138116 600004 138136
rect 600004 138116 600006 138136
rect 599950 138080 600006 138116
rect 599858 137128 599914 137184
rect 599950 136040 600006 136096
rect 599858 135088 599914 135144
rect 599306 133048 599362 133104
rect 599950 134000 600006 134056
rect 598938 131960 598994 132016
rect 599858 131008 599914 131064
rect 599950 129920 600006 129976
rect 599858 128968 599914 129024
rect 582286 128152 582342 128208
rect 581734 120536 581790 120592
rect 581550 117544 581606 117600
rect 581182 114416 581238 114472
rect 581090 109928 581146 109984
rect 580906 102312 580962 102368
rect 580814 93200 580870 93256
rect 580630 91704 580686 91760
rect 194414 42200 194470 42256
rect 187606 41792 187662 41848
rect 209778 41248 209834 41304
rect 212446 41248 212502 41304
rect 218058 41248 218114 41304
rect 230478 10648 230534 10704
rect 230846 16632 230902 16688
rect 230754 13640 230810 13696
rect 415490 41928 415546 41984
rect 307298 41792 307354 41848
rect 362038 41792 362094 41848
rect 470322 41792 470378 41848
rect 518530 42064 518586 42120
rect 521658 42064 521714 42120
rect 524050 41928 524106 41984
rect 529662 41928 529718 41984
rect 535458 41928 535514 41984
rect 579618 82628 579620 82648
rect 579620 82628 579672 82648
rect 579672 82628 579674 82648
rect 579618 82592 579674 82628
rect 580722 65864 580778 65920
rect 580814 64368 580870 64424
rect 579618 59744 579674 59800
rect 579618 58248 579674 58304
rect 581366 115912 581422 115968
rect 581274 77968 581330 78024
rect 581366 74976 581422 75032
rect 581642 81096 581698 81152
rect 582010 90208 582066 90264
rect 599950 127880 600006 127936
rect 600042 126928 600098 126984
rect 599858 125840 599914 125896
rect 599950 124888 600006 124944
rect 598938 123800 598994 123856
rect 599858 122848 599914 122904
rect 582194 94696 582250 94752
rect 599950 121760 600006 121816
rect 600042 120808 600098 120864
rect 599858 119720 599914 119776
rect 582286 88576 582342 88632
rect 582102 87080 582158 87136
rect 581918 85584 581974 85640
rect 581826 84088 581882 84144
rect 581734 79464 581790 79520
rect 581550 76472 581606 76528
rect 581458 71984 581514 72040
rect 581182 70352 581238 70408
rect 581090 67360 581146 67416
rect 582010 62872 582066 62928
rect 581918 56752 581974 56808
rect 599950 118788 600006 118824
rect 599950 118768 599952 118788
rect 599952 118768 600004 118788
rect 600004 118768 600006 118788
rect 599858 117680 599914 117736
rect 599950 116728 600006 116784
rect 599858 115640 599914 115696
rect 599950 114688 600006 114744
rect 599950 112648 600006 112704
rect 599766 111560 599822 111616
rect 600226 110608 600282 110664
rect 599950 109520 600006 109576
rect 599950 107480 600006 107536
rect 599950 100408 600006 100464
rect 582286 68856 582342 68912
rect 582194 61240 582250 61296
rect 582102 55256 582158 55312
rect 580906 53760 580962 53816
rect 600318 108568 600374 108624
rect 600410 106528 600466 106584
rect 600594 105440 600650 105496
rect 600502 103400 600558 103456
rect 600686 104488 600742 104544
rect 600870 102448 600926 102504
rect 600778 101360 600834 101416
rect 622490 87896 622546 87952
rect 622306 86944 622362 87000
rect 621938 84088 621994 84144
rect 623226 88848 623282 88904
rect 623778 90616 623834 90672
rect 628286 95920 628342 95976
rect 640522 95684 640524 95704
rect 640524 95684 640576 95704
rect 640576 95684 640578 95704
rect 640522 95648 640578 95684
rect 627918 94424 627974 94480
rect 627274 93472 627330 93528
rect 626446 92520 626502 92576
rect 625894 91568 625950 91624
rect 623962 89664 624018 89720
rect 623410 85992 623466 86048
rect 623318 85040 623374 85096
rect 623134 83136 623190 83192
rect 622306 82184 622362 82240
rect 622490 81368 622546 81424
rect 641258 43560 641314 43616
rect 641166 42916 641168 42936
rect 641168 42916 641220 42936
rect 641220 42916 641222 42936
rect 641166 42880 641222 42916
rect 641258 42200 641314 42256
rect 594706 41792 594762 41848
rect 590750 41656 590806 41712
rect 565818 41520 565874 41576
rect 642730 92656 642786 92712
rect 645950 89664 646006 89720
rect 646042 87080 646098 87136
rect 653218 92520 653274 92576
rect 655334 93336 655390 93392
rect 654046 91432 654102 91488
rect 653494 90616 653550 90672
rect 656990 90344 657046 90400
rect 662234 95512 662290 95568
rect 657358 94696 657414 94752
rect 663246 93744 663302 93800
rect 663338 93064 663394 93120
rect 663430 92248 663486 92304
rect 663246 91024 663302 91080
rect 663522 89528 663578 89584
rect 663706 90344 663762 90400
rect 662142 88712 662198 88768
rect 646134 84632 646190 84688
rect 645858 82184 645914 82240
rect 666742 183776 666798 183832
rect 666742 180376 666798 180432
rect 666742 178744 666798 178800
rect 669134 983320 669190 983376
rect 668766 667256 668822 667312
rect 668674 621560 668730 621616
rect 666742 175344 666798 175400
rect 666742 173576 666798 173632
rect 666742 170176 666798 170232
rect 666742 168544 666798 168600
rect 666742 165144 666798 165200
rect 666742 163512 666798 163568
rect 666742 160112 666798 160168
rect 666742 158344 666798 158400
rect 666742 154944 666798 155000
rect 666742 153312 666798 153368
rect 666742 149912 666798 149968
rect 666650 148144 666706 148200
rect 666650 144880 666706 144936
rect 666650 143112 666706 143168
rect 666650 139712 666706 139768
rect 666650 132912 666706 132968
rect 672722 985496 672778 985552
rect 669686 983184 669742 983240
rect 670238 983048 670294 983104
rect 670054 982912 670110 982968
rect 669778 759192 669834 759248
rect 672538 985360 672594 985416
rect 671066 209208 671122 209264
rect 671066 205808 671122 205864
rect 670974 204176 671030 204232
rect 670974 200776 671030 200832
rect 670882 199008 670938 199064
rect 670882 195608 670938 195664
rect 670790 193976 670846 194032
rect 670790 190576 670846 190632
rect 670698 188944 670754 189000
rect 670698 185544 670754 185600
rect 670698 138080 670754 138136
rect 670698 134680 670754 134736
rect 666650 129512 666706 129568
rect 666650 127880 666706 127936
rect 666650 124480 666706 124536
rect 666650 122848 666706 122904
rect 666650 119448 666706 119504
rect 670790 104080 670846 104136
rect 671802 173576 671858 173632
rect 672078 183776 672134 183832
rect 672170 178744 672226 178800
rect 671434 112648 671490 112704
rect 671158 107480 671214 107536
rect 672354 168544 672410 168600
rect 672170 116048 672226 116104
rect 672078 114280 672134 114336
rect 675666 938712 675722 938768
rect 676310 939664 676366 939720
rect 676126 939256 676182 939312
rect 676218 938868 676274 938904
rect 676218 938848 676220 938868
rect 676220 938848 676272 938868
rect 676272 938848 676274 938868
rect 678978 937624 679034 937680
rect 676218 936400 676274 936456
rect 676034 935856 676090 935912
rect 675942 935468 675998 935504
rect 675942 935448 675944 935468
rect 675944 935448 675996 935468
rect 675996 935448 675998 935468
rect 675758 934632 675814 934688
rect 676034 935040 676090 935096
rect 675942 934224 675998 934280
rect 676126 933952 676182 934008
rect 676034 933408 676090 933464
rect 676034 933000 676090 933056
rect 675942 932184 675998 932240
rect 676126 932764 676128 932784
rect 676128 932764 676180 932784
rect 676180 932764 676182 932784
rect 676126 932728 676182 932764
rect 676034 931776 676090 931832
rect 676034 931368 676090 931424
rect 675942 930960 675998 931016
rect 676126 930688 676182 930744
rect 676034 930144 676090 930200
rect 678978 929464 679034 929520
rect 678978 929056 679034 929112
rect 684498 929056 684554 929112
rect 684498 928648 684554 928704
rect 675758 877240 675814 877296
rect 675666 876560 675722 876616
rect 675390 875880 675446 875936
rect 675482 873976 675538 874032
rect 673458 760280 673514 760336
rect 673458 759192 673514 759248
rect 675758 872208 675814 872264
rect 674286 797680 674342 797736
rect 674194 791968 674250 792024
rect 674378 777416 674434 777472
rect 675390 787752 675446 787808
rect 675390 787344 675446 787400
rect 675390 786800 675446 786856
rect 675390 784080 675446 784136
rect 675482 783808 675538 783864
rect 674194 770208 674250 770264
rect 673642 699760 673698 699816
rect 672446 163512 672502 163568
rect 675574 753752 675630 753808
rect 675482 744096 675538 744152
rect 679070 772656 679126 772712
rect 678978 761232 679034 761288
rect 676218 760824 676274 760880
rect 676126 760416 676182 760472
rect 676310 759600 676366 759656
rect 676034 759092 676036 759112
rect 676036 759092 676088 759112
rect 676088 759092 676090 759112
rect 676034 759056 676090 759092
rect 679070 759600 679126 759656
rect 678978 758376 679034 758432
rect 676126 757968 676182 758024
rect 676034 756608 676090 756664
rect 676310 757560 676366 757616
rect 676218 757152 676274 757208
rect 676126 755520 676182 755576
rect 676034 754976 676090 755032
rect 676034 754160 676090 754216
rect 676034 753344 676090 753400
rect 676034 752936 676090 752992
rect 679254 751032 679310 751088
rect 678978 750624 679034 750680
rect 679254 750624 679310 750680
rect 678978 750216 679034 750272
rect 675666 743960 675722 744016
rect 675758 742872 675814 742928
rect 675758 742464 675814 742520
rect 675482 741648 675538 741704
rect 675390 739744 675446 739800
rect 675390 739064 675446 739120
rect 675666 738520 675722 738576
rect 675758 737976 675814 738032
rect 676034 716524 676036 716544
rect 676036 716524 676088 716544
rect 676088 716524 676090 716544
rect 676034 716488 676090 716524
rect 676034 716116 676036 716136
rect 676036 716116 676088 716136
rect 676088 716116 676090 716136
rect 676034 716080 676090 716116
rect 676034 715708 676036 715728
rect 676036 715708 676088 715728
rect 676088 715708 676090 715728
rect 676034 715672 676090 715708
rect 676034 715284 676090 715320
rect 676034 715264 676036 715284
rect 676036 715264 676088 715284
rect 676088 715264 676090 715284
rect 676034 714892 676036 714912
rect 676036 714892 676088 714912
rect 676088 714892 676090 714912
rect 676034 714856 676090 714892
rect 678978 714448 679034 714504
rect 674010 699624 674066 699680
rect 672538 158344 672594 158400
rect 672630 153312 672686 153368
rect 674378 608912 674434 608968
rect 676034 714060 676090 714096
rect 676034 714040 676036 714060
rect 676036 714040 676088 714060
rect 676088 714040 676090 714060
rect 676034 713652 676090 713688
rect 676034 713632 676036 713652
rect 676036 713632 676088 713652
rect 676088 713632 676090 713652
rect 676034 713244 676090 713280
rect 676034 713224 676036 713244
rect 676036 713224 676088 713244
rect 676088 713224 676090 713244
rect 676034 712852 676036 712872
rect 676036 712852 676088 712872
rect 676088 712852 676090 712872
rect 676034 712816 676090 712852
rect 676034 712444 676036 712464
rect 676036 712444 676088 712464
rect 676088 712444 676090 712464
rect 676034 712408 676090 712444
rect 675850 711592 675906 711648
rect 675850 710504 675906 710560
rect 676034 710776 676090 710832
rect 676586 710538 676642 710594
rect 675942 710368 675998 710424
rect 676034 709960 676090 710016
rect 676034 708328 676090 708384
rect 676034 707920 676090 707976
rect 676034 707512 676090 707568
rect 675850 707104 675906 707160
rect 676034 706696 676090 706752
rect 675942 706288 675998 706344
rect 676034 705880 676090 705936
rect 675942 705492 675998 705528
rect 675942 705472 675944 705492
rect 675944 705472 675996 705492
rect 675996 705472 675998 705492
rect 676034 705064 676090 705120
rect 675666 699488 675722 699544
rect 675482 698128 675538 698184
rect 675390 697312 675446 697368
rect 675390 696632 675446 696688
rect 675390 694728 675446 694784
rect 675482 694320 675538 694376
rect 675390 693504 675446 693560
rect 675758 692960 675814 693016
rect 675758 690104 675814 690160
rect 676218 671064 676274 671120
rect 676034 670964 676036 670984
rect 676036 670964 676088 670984
rect 676088 670964 676090 670984
rect 676034 670928 676090 670964
rect 676034 670556 676036 670576
rect 676036 670556 676088 670576
rect 676088 670556 676090 670576
rect 676034 670520 676090 670556
rect 676218 670284 676220 670304
rect 676220 670284 676272 670304
rect 676272 670284 676274 670304
rect 676218 670248 676274 670284
rect 676034 669704 676090 669760
rect 678978 669432 679034 669488
rect 676034 668888 676090 668944
rect 675942 668092 675998 668128
rect 675942 668072 675944 668092
rect 675944 668072 675996 668092
rect 675996 668072 675998 668092
rect 676218 668652 676220 668672
rect 676220 668652 676272 668672
rect 676272 668652 676274 668672
rect 676218 668616 676274 668652
rect 675942 667700 675944 667720
rect 675944 667700 675996 667720
rect 675996 667700 675998 667720
rect 675942 667664 675998 667700
rect 676126 666576 676182 666632
rect 676034 665216 676090 665272
rect 676126 664944 676182 665000
rect 676034 663176 676090 663232
rect 678978 660864 679034 660920
rect 678978 660456 679034 660512
rect 684498 660456 684554 660512
rect 684498 660048 684554 660104
rect 675390 652840 675446 652896
rect 675482 652160 675538 652216
rect 675390 651616 675446 651672
rect 675390 648896 675446 648952
rect 675758 648624 675814 648680
rect 675482 608776 675538 608832
rect 678978 626048 679034 626104
rect 676126 625640 676182 625696
rect 676034 625096 676090 625152
rect 676310 625232 676366 625288
rect 676218 624416 676274 624472
rect 676034 623908 676036 623928
rect 676036 623908 676088 623928
rect 676088 623908 676090 623928
rect 676034 623872 676090 623908
rect 679070 624416 679126 624472
rect 679162 623600 679218 623656
rect 678978 623192 679034 623248
rect 676218 621968 676274 622024
rect 676034 621424 676090 621480
rect 676126 620336 676182 620392
rect 676034 619792 676090 619848
rect 676034 618196 676036 618216
rect 676036 618196 676088 618216
rect 676088 618196 676090 618216
rect 676034 618160 676090 618196
rect 676218 617924 676220 617944
rect 676220 617924 676272 617944
rect 676272 617924 676274 617944
rect 676218 617888 676274 617924
rect 676218 616700 676220 616720
rect 676220 616700 676272 616720
rect 676272 616700 676274 616720
rect 676218 616664 676274 616700
rect 679254 615848 679310 615904
rect 678978 615440 679034 615496
rect 679254 615440 679310 615496
rect 678978 615032 679034 615088
rect 675666 607552 675722 607608
rect 675758 607280 675814 607336
rect 675390 606464 675446 606520
rect 675390 604696 675446 604752
rect 675482 604288 675538 604344
rect 675482 603472 675538 603528
rect 675758 602928 675814 602984
rect 675390 574504 675446 574560
rect 676126 580896 676182 580952
rect 676310 580488 676366 580544
rect 676218 580100 676274 580136
rect 676218 580080 676220 580100
rect 676220 580080 676272 580100
rect 676272 580080 676274 580100
rect 676034 579808 676090 579864
rect 676218 579284 676274 579320
rect 676218 579264 676220 579284
rect 676220 579264 676272 579284
rect 676272 579264 676274 579284
rect 678978 579264 679034 579320
rect 676218 578468 676274 578504
rect 676218 578448 676220 578468
rect 676220 578448 676272 578468
rect 676272 578448 676274 578468
rect 676218 577652 676274 577688
rect 676218 577632 676220 577652
rect 676220 577632 676272 577652
rect 676272 577632 676274 577652
rect 676218 577224 676274 577280
rect 676034 576972 676090 577008
rect 676034 576952 676036 576972
rect 676036 576952 676088 576972
rect 676088 576952 676090 576972
rect 676034 576136 676090 576192
rect 675574 575320 675630 575376
rect 676034 574912 676090 574968
rect 676034 572872 676090 572928
rect 676034 572464 676090 572520
rect 676034 572056 676090 572112
rect 678978 570696 679034 570752
rect 678978 570288 679034 570344
rect 684498 570288 684554 570344
rect 684498 569880 684554 569936
rect 675482 564440 675538 564496
rect 675482 562400 675538 562456
rect 675758 561992 675814 562048
rect 675482 561176 675538 561232
rect 675390 558728 675446 558784
rect 675758 558320 675814 558376
rect 675758 557504 675814 557560
rect 676218 535880 676274 535936
rect 676034 535676 676090 535732
rect 678978 535064 679034 535120
rect 676034 534896 676036 534916
rect 676036 534896 676088 534916
rect 676088 534896 676090 534916
rect 676034 534860 676090 534896
rect 676126 534248 676182 534304
rect 676034 533264 676036 533284
rect 676036 533264 676088 533284
rect 676088 533264 676090 533284
rect 676034 533228 676090 533264
rect 675942 532820 675998 532876
rect 679070 534248 679126 534304
rect 679070 533432 679126 533488
rect 675758 532004 675814 532060
rect 675666 488824 675722 488880
rect 675206 488044 675208 488064
rect 675208 488044 675260 488064
rect 675260 488044 675262 488064
rect 675206 488008 675262 488044
rect 676218 532636 676274 532672
rect 676218 532616 676220 532636
rect 676220 532616 676272 532636
rect 676272 532616 676274 532636
rect 676034 531188 676090 531244
rect 676034 529964 676090 530020
rect 676034 529556 676090 529612
rect 676034 527924 676090 527980
rect 676034 527516 676090 527572
rect 676034 526292 676090 526348
rect 678978 525680 679034 525736
rect 678978 525272 679034 525328
rect 684590 525272 684646 525328
rect 684590 524864 684646 524920
rect 676034 492088 676090 492144
rect 675942 491680 675998 491736
rect 676034 491272 676090 491328
rect 675850 490864 675906 490920
rect 675942 490456 675998 490512
rect 675850 489640 675906 489696
rect 675758 488416 675814 488472
rect 672814 278432 672870 278488
rect 672722 148144 672778 148200
rect 672354 117680 672410 117736
rect 672262 109248 672318 109304
rect 676034 490048 676090 490104
rect 676034 489232 676090 489288
rect 676034 488008 676090 488064
rect 676034 487192 676090 487248
rect 675942 486376 675998 486432
rect 676034 485968 676090 486024
rect 676034 485560 676090 485616
rect 676034 483928 676090 483984
rect 676034 483520 676090 483576
rect 675942 482704 675998 482760
rect 676034 482296 676090 482352
rect 676034 481888 676090 481944
rect 675942 481480 675998 481536
rect 676034 481108 676036 481128
rect 676036 481108 676088 481128
rect 676088 481108 676090 481128
rect 676034 481072 676090 481108
rect 675942 480664 675998 480720
rect 675942 403436 675998 403472
rect 675942 403416 675944 403436
rect 675944 403416 675996 403436
rect 675996 403416 675998 403436
rect 675942 403008 675998 403064
rect 675850 401784 675906 401840
rect 675666 401376 675722 401432
rect 675574 400968 675630 401024
rect 675298 396888 675354 396944
rect 675758 400560 675814 400616
rect 676218 403688 676274 403744
rect 676126 402872 676182 402928
rect 676126 402056 676182 402112
rect 676034 400152 676090 400208
rect 676034 399744 676090 399800
rect 676034 399336 676090 399392
rect 675850 398520 675906 398576
rect 676126 398792 676182 398848
rect 676034 398112 676090 398168
rect 675942 397704 675998 397760
rect 676034 397296 676090 397352
rect 676034 396480 676090 396536
rect 675942 395664 675998 395720
rect 675942 395256 675998 395312
rect 676126 395936 676182 395992
rect 676034 394848 676090 394904
rect 676034 394440 676090 394496
rect 676034 394032 676090 394088
rect 678978 393488 679034 393544
rect 678978 393080 679034 393136
rect 684498 393080 684554 393136
rect 684498 392672 684554 392728
rect 674746 357448 674802 357504
rect 672998 343576 673054 343632
rect 672906 143112 672962 143168
rect 673182 343576 673238 343632
rect 675574 357060 675630 357096
rect 675574 357040 675576 357060
rect 675576 357040 675628 357060
rect 675628 357040 675630 357060
rect 675666 356632 675722 356688
rect 675850 358672 675906 358728
rect 675942 358264 675998 358320
rect 676034 357856 676090 357912
rect 676034 356224 676090 356280
rect 675758 355816 675814 355872
rect 676034 355428 676090 355464
rect 676034 355408 676036 355428
rect 676036 355408 676088 355428
rect 676088 355408 676090 355428
rect 675298 355000 675354 355056
rect 676034 354612 676090 354648
rect 676034 354592 676036 354612
rect 676036 354592 676088 354612
rect 676088 354592 676090 354612
rect 676034 354184 676090 354240
rect 676034 353368 676090 353424
rect 676034 352960 676090 353016
rect 675942 352552 675998 352608
rect 675298 351736 675354 351792
rect 676034 351328 676090 351384
rect 675942 350920 675998 350976
rect 676034 350104 676090 350160
rect 676034 349696 676090 349752
rect 675942 349288 675998 349344
rect 675850 348880 675906 348936
rect 675758 348472 675814 348528
rect 675666 348064 675722 348120
rect 675758 347656 675814 347712
rect 675666 347248 675722 347304
rect 675666 330520 675722 330576
rect 675758 328344 675814 328400
rect 675758 326848 675814 326904
rect 676218 313520 676274 313576
rect 676034 313284 676036 313304
rect 676036 313284 676088 313304
rect 676088 313284 676090 313304
rect 676034 313248 676090 313284
rect 676034 312876 676036 312896
rect 676036 312876 676088 312896
rect 676088 312876 676090 312896
rect 676034 312840 676090 312876
rect 676034 312468 676036 312488
rect 676036 312468 676088 312488
rect 676088 312468 676090 312488
rect 676034 312432 676090 312468
rect 676034 312060 676036 312080
rect 676036 312060 676088 312080
rect 676088 312060 676090 312080
rect 676034 312024 676090 312060
rect 676034 311652 676036 311672
rect 676036 311652 676088 311672
rect 676088 311652 676090 311672
rect 676034 311616 676090 311652
rect 676034 311208 676090 311264
rect 672998 138080 673054 138136
rect 676034 310836 676036 310856
rect 676036 310836 676088 310856
rect 676088 310836 676090 310856
rect 676034 310800 676090 310836
rect 676034 310428 676036 310448
rect 676036 310428 676088 310448
rect 676088 310428 676090 310448
rect 676034 310392 676090 310428
rect 676034 310020 676036 310040
rect 676036 310020 676088 310040
rect 676088 310020 676090 310040
rect 676034 309984 676090 310020
rect 676034 309612 676036 309632
rect 676036 309612 676088 309632
rect 676088 309612 676090 309632
rect 676034 309576 676090 309612
rect 676034 309188 676090 309224
rect 676034 309168 676036 309188
rect 676036 309168 676088 309188
rect 676088 309168 676090 309188
rect 676034 308760 676090 308816
rect 675758 308352 675814 308408
rect 676034 307944 676090 308000
rect 675942 307128 675998 307184
rect 676126 307400 676182 307456
rect 676034 306720 676090 306776
rect 676034 305904 676090 305960
rect 676126 305360 676182 305416
rect 676126 304952 676182 305008
rect 676034 304680 676090 304736
rect 675942 303864 675998 303920
rect 676126 304136 676182 304192
rect 679070 303320 679126 303376
rect 679070 302912 679126 302968
rect 684498 302912 684554 302968
rect 684498 302504 684554 302560
rect 675758 292168 675814 292224
rect 676126 268504 676182 268560
rect 676034 267824 676090 267880
rect 676218 268116 676274 268152
rect 676218 268096 676220 268116
rect 676220 268096 676272 268116
rect 676272 268096 676274 268116
rect 675942 267452 675944 267472
rect 675944 267452 675996 267472
rect 675996 267452 675998 267472
rect 675942 267416 675998 267452
rect 675758 267008 675814 267064
rect 675666 265376 675722 265432
rect 675574 260480 675630 260536
rect 675574 260072 675630 260128
rect 676034 266600 676090 266656
rect 676034 266192 676090 266248
rect 676218 266092 676220 266112
rect 676220 266092 676272 266112
rect 676272 266092 676274 266112
rect 676218 266056 676274 266092
rect 676218 264832 676274 264888
rect 676034 264152 676090 264208
rect 675850 263336 675906 263392
rect 676126 263608 676182 263664
rect 676034 262928 676090 262984
rect 675942 262520 675998 262576
rect 676034 262112 676090 262168
rect 676034 261704 676090 261760
rect 675942 260888 675998 260944
rect 676126 261160 676182 261216
rect 676126 259548 676182 259584
rect 676126 259528 676128 259548
rect 676128 259528 676180 259548
rect 676180 259528 676182 259548
rect 676034 259256 676090 259312
rect 676126 258712 676182 258768
rect 678978 258304 679034 258360
rect 678978 257896 679034 257952
rect 684498 257896 684554 257952
rect 684498 257488 684554 257544
rect 673090 132912 673146 132968
rect 672814 127880 672870 127936
rect 675574 221856 675630 221912
rect 704002 224304 704058 224360
rect 704462 224168 704518 224224
rect 708510 224168 708566 224224
rect 708970 224304 709026 224360
rect 676034 223488 676090 223544
rect 675850 223080 675906 223136
rect 675758 222264 675814 222320
rect 675758 221448 675814 221504
rect 675758 221040 675814 221096
rect 675942 222672 675998 222728
rect 675666 220632 675722 220688
rect 675390 212492 675446 212528
rect 675390 212472 675392 212492
rect 675392 212472 675444 212492
rect 675444 212472 675446 212492
rect 675666 216960 675722 217016
rect 675942 220224 675998 220280
rect 676034 219408 676090 219464
rect 676034 219000 676090 219056
rect 675942 218592 675998 218648
rect 676034 218184 676090 218240
rect 676034 217776 676090 217832
rect 675942 217368 675998 217424
rect 675758 216552 675814 216608
rect 676034 216144 676090 216200
rect 675942 215736 675998 215792
rect 675850 215328 675906 215384
rect 676034 214920 676090 214976
rect 676034 214512 676090 214568
rect 675942 214104 675998 214160
rect 675942 213696 675998 213752
rect 675850 212880 675906 212936
rect 675850 212064 675906 212120
rect 675758 178472 675814 178528
rect 703910 179288 703966 179344
rect 709062 179288 709118 179344
rect 675942 178064 675998 178120
rect 675850 177248 675906 177304
rect 676034 177656 676090 177712
rect 675942 176876 675944 176896
rect 675944 176876 675996 176896
rect 675996 176876 675998 176896
rect 675942 176840 675998 176876
rect 676034 176432 676090 176488
rect 675942 176044 675998 176080
rect 675942 176024 675944 176044
rect 675944 176024 675996 176044
rect 675996 176024 675998 176044
rect 676034 175616 676090 175672
rect 675942 175244 675944 175264
rect 675944 175244 675996 175264
rect 675996 175244 675998 175264
rect 675942 175208 675998 175244
rect 676034 174800 676090 174856
rect 676034 174428 676036 174448
rect 676036 174428 676088 174448
rect 676088 174428 676090 174448
rect 676034 174392 676090 174428
rect 676034 173984 676090 174040
rect 675758 173168 675814 173224
rect 676034 172760 676090 172816
rect 675942 172352 675998 172408
rect 676034 171536 676090 171592
rect 675942 171164 675944 171184
rect 675944 171164 675996 171184
rect 675996 171164 675998 171184
rect 675942 171128 675998 171164
rect 676034 170720 676090 170776
rect 675942 170312 675998 170368
rect 675942 169904 675998 169960
rect 676034 169496 676090 169552
rect 675942 169088 675998 169144
rect 675850 168680 675906 168736
rect 676034 168292 676090 168328
rect 676034 168272 676036 168292
rect 676036 168272 676088 168292
rect 676088 168272 676090 168292
rect 676034 167884 676090 167920
rect 676034 167864 676036 167884
rect 676036 167864 676088 167884
rect 676088 167864 676090 167884
rect 676034 167476 676090 167512
rect 676034 167456 676036 167476
rect 676036 167456 676088 167476
rect 676088 167456 676090 167476
rect 675758 148416 675814 148472
rect 675758 146240 675814 146296
rect 703818 134136 703874 134192
rect 709062 134136 709118 134192
rect 676126 133048 676182 133104
rect 676034 132912 676090 132968
rect 676218 132640 676274 132696
rect 676218 132268 676220 132288
rect 676220 132268 676272 132288
rect 676272 132268 676274 132288
rect 676218 132232 676274 132268
rect 676034 131708 676090 131744
rect 676034 131688 676036 131708
rect 676036 131688 676088 131708
rect 676088 131688 676090 131708
rect 676218 131452 676220 131472
rect 676220 131452 676272 131472
rect 676272 131452 676274 131472
rect 676218 131416 676274 131452
rect 676034 130892 676090 130928
rect 676034 130872 676036 130892
rect 676036 130872 676088 130892
rect 676088 130872 676090 130892
rect 676218 130636 676220 130656
rect 676220 130636 676272 130656
rect 676272 130636 676274 130656
rect 676218 130600 676274 130636
rect 676034 130076 676090 130112
rect 676034 130056 676036 130076
rect 676036 130056 676088 130076
rect 676088 130056 676090 130076
rect 676034 129684 676036 129704
rect 676036 129684 676088 129704
rect 676088 129684 676090 129704
rect 676034 129648 676090 129684
rect 676218 129412 676220 129432
rect 676220 129412 676272 129432
rect 676272 129412 676274 129432
rect 676218 129376 676274 129412
rect 676034 128832 676090 128888
rect 675758 128016 675814 128072
rect 673182 122848 673238 122904
rect 672906 110880 672962 110936
rect 672446 105848 672502 105904
rect 676034 127608 676090 127664
rect 675942 127200 675998 127256
rect 676034 126384 676090 126440
rect 675942 125976 675998 126032
rect 675850 125160 675906 125216
rect 675850 124752 675906 124808
rect 675942 124344 675998 124400
rect 676126 125296 676182 125352
rect 676034 123936 676090 123992
rect 675942 123528 675998 123584
rect 676034 123140 676090 123176
rect 676034 123120 676036 123140
rect 676036 123120 676088 123140
rect 676088 123120 676090 123140
rect 676034 122732 676090 122768
rect 676034 122712 676036 122732
rect 676036 122712 676088 122732
rect 676088 122712 676090 122732
rect 676034 122324 676090 122360
rect 676034 122304 676036 122324
rect 676036 122304 676088 122324
rect 676088 122304 676090 122324
rect 675758 103264 675814 103320
rect 671986 102448 672042 102504
rect 675758 101360 675814 101416
rect 670882 100816 670938 100872
rect 646318 45056 646374 45112
rect 642638 41248 642694 41304
rect 231030 15136 231086 15192
rect 230938 12144 230994 12200
rect 230662 9152 230718 9208
rect 230570 7656 230626 7712
rect 230386 6160 230442 6216
<< metal3 >>
rect 425973 1006090 426039 1006093
rect 425776 1006088 426039 1006090
rect 425776 1006032 425978 1006088
rect 426034 1006032 426039 1006088
rect 425776 1006030 426039 1006032
rect 425973 1006027 426039 1006030
rect 424317 1005954 424383 1005957
rect 424120 1005952 424383 1005954
rect 424120 1005896 424322 1005952
rect 424378 1005896 424383 1005952
rect 424120 1005894 424383 1005896
rect 424317 1005891 424383 1005894
rect 423857 1005818 423923 1005821
rect 423752 1005816 423923 1005818
rect 423752 1005760 423862 1005816
rect 423918 1005760 423923 1005816
rect 423752 1005758 423923 1005760
rect 423857 1005755 423923 1005758
rect 356053 1005682 356119 1005685
rect 504541 1005682 504607 1005685
rect 505001 1005682 505067 1005685
rect 355948 1005680 356119 1005682
rect 355948 1005624 356058 1005680
rect 356114 1005624 356119 1005680
rect 355948 1005622 356119 1005624
rect 504436 1005680 504607 1005682
rect 504436 1005624 504546 1005680
rect 504602 1005624 504607 1005680
rect 504436 1005622 504607 1005624
rect 504804 1005680 505067 1005682
rect 504804 1005624 505006 1005680
rect 505062 1005624 505067 1005680
rect 504804 1005622 505067 1005624
rect 356053 1005619 356119 1005622
rect 504541 1005619 504607 1005622
rect 505001 1005619 505067 1005622
rect 356881 1005546 356947 1005549
rect 502977 1005546 503043 1005549
rect 505369 1005546 505435 1005549
rect 356684 1005544 356947 1005546
rect 356684 1005488 356886 1005544
rect 356942 1005488 356947 1005544
rect 356684 1005486 356947 1005488
rect 502780 1005544 503043 1005546
rect 502780 1005488 502982 1005544
rect 503038 1005488 503043 1005544
rect 502780 1005486 503043 1005488
rect 505172 1005544 505435 1005546
rect 505172 1005488 505374 1005544
rect 505430 1005488 505435 1005544
rect 505172 1005486 505435 1005488
rect 356881 1005483 356947 1005486
rect 502977 1005483 503043 1005486
rect 505369 1005483 505435 1005486
rect 160277 1005410 160343 1005413
rect 209221 1005410 209287 1005413
rect 356513 1005410 356579 1005413
rect 361021 1005410 361087 1005413
rect 425145 1005410 425211 1005413
rect 428365 1005410 428431 1005413
rect 505829 1005410 505895 1005413
rect 160277 1005408 160540 1005410
rect 160277 1005352 160282 1005408
rect 160338 1005352 160540 1005408
rect 160277 1005350 160540 1005352
rect 209024 1005408 209287 1005410
rect 209024 1005352 209226 1005408
rect 209282 1005352 209287 1005408
rect 209024 1005350 209287 1005352
rect 356316 1005408 356579 1005410
rect 356316 1005352 356518 1005408
rect 356574 1005352 356579 1005408
rect 356316 1005350 356579 1005352
rect 360824 1005408 361087 1005410
rect 360824 1005352 361026 1005408
rect 361082 1005352 361087 1005408
rect 360824 1005350 361087 1005352
rect 424948 1005408 425211 1005410
rect 424948 1005352 425150 1005408
rect 425206 1005352 425211 1005408
rect 424948 1005350 425211 1005352
rect 428260 1005408 428431 1005410
rect 428260 1005352 428370 1005408
rect 428426 1005352 428431 1005408
rect 428260 1005350 428431 1005352
rect 505632 1005408 505895 1005410
rect 505632 1005352 505834 1005408
rect 505890 1005352 505895 1005408
rect 505632 1005350 505895 1005352
rect 160277 1005347 160343 1005350
rect 209221 1005347 209287 1005350
rect 356513 1005347 356579 1005350
rect 361021 1005347 361087 1005350
rect 425145 1005347 425211 1005350
rect 428365 1005347 428431 1005350
rect 505829 1005347 505895 1005350
rect 106457 1005274 106523 1005277
rect 106260 1005272 106523 1005274
rect 106260 1005216 106462 1005272
rect 106518 1005216 106523 1005272
rect 106260 1005214 106523 1005216
rect 106457 1005211 106523 1005214
rect 109309 1005274 109375 1005277
rect 259821 1005274 259887 1005277
rect 260189 1005274 260255 1005277
rect 360193 1005274 360259 1005277
rect 109309 1005272 109480 1005274
rect 109309 1005216 109314 1005272
rect 109370 1005216 109480 1005272
rect 109309 1005214 109480 1005216
rect 259624 1005272 259887 1005274
rect 259624 1005216 259826 1005272
rect 259882 1005216 259887 1005272
rect 259624 1005214 259887 1005216
rect 260084 1005272 260255 1005274
rect 260084 1005216 260194 1005272
rect 260250 1005216 260255 1005272
rect 260084 1005214 260255 1005216
rect 359996 1005272 360259 1005274
rect 359996 1005216 360198 1005272
rect 360254 1005216 360259 1005272
rect 359996 1005214 360259 1005216
rect 109309 1005211 109375 1005214
rect 259821 1005211 259887 1005214
rect 260189 1005211 260255 1005214
rect 360193 1005211 360259 1005214
rect 105629 1005138 105695 1005141
rect 201493 1005138 201559 1005141
rect 202321 1005138 202387 1005141
rect 105432 1005136 105695 1005138
rect 105432 1005080 105634 1005136
rect 105690 1005080 105695 1005136
rect 105432 1005078 105695 1005080
rect 201296 1005136 201559 1005138
rect 201296 1005080 201498 1005136
rect 201554 1005080 201559 1005136
rect 201296 1005078 201559 1005080
rect 202124 1005136 202387 1005138
rect 202124 1005080 202326 1005136
rect 202382 1005080 202387 1005136
rect 202124 1005078 202387 1005080
rect 105629 1005075 105695 1005078
rect 201493 1005075 201559 1005078
rect 202321 1005075 202387 1005078
rect 209589 1005138 209655 1005141
rect 210877 1005138 210943 1005141
rect 261017 1005138 261083 1005141
rect 263041 1005138 263107 1005141
rect 209589 1005136 209852 1005138
rect 209589 1005080 209594 1005136
rect 209650 1005080 209852 1005136
rect 209589 1005078 209852 1005080
rect 210680 1005136 210943 1005138
rect 210680 1005080 210882 1005136
rect 210938 1005080 210943 1005136
rect 210680 1005078 210943 1005080
rect 260820 1005136 261083 1005138
rect 260820 1005080 261022 1005136
rect 261078 1005080 261083 1005136
rect 260820 1005078 261083 1005080
rect 262844 1005136 263107 1005138
rect 262844 1005080 263046 1005136
rect 263102 1005080 263107 1005136
rect 262844 1005078 263107 1005080
rect 209589 1005075 209655 1005078
rect 210877 1005075 210943 1005078
rect 261017 1005075 261083 1005078
rect 263041 1005075 263107 1005078
rect 264329 1005138 264395 1005141
rect 269205 1005138 269271 1005141
rect 427537 1005138 427603 1005141
rect 428825 1005138 428891 1005141
rect 502517 1005138 502583 1005141
rect 264329 1005136 269271 1005138
rect 264329 1005080 264334 1005136
rect 264390 1005080 269210 1005136
rect 269266 1005080 269271 1005136
rect 264329 1005078 269271 1005080
rect 427340 1005136 427603 1005138
rect 427340 1005080 427542 1005136
rect 427598 1005080 427603 1005136
rect 427340 1005078 427603 1005080
rect 428628 1005136 428891 1005138
rect 428628 1005080 428830 1005136
rect 428886 1005080 428891 1005136
rect 428628 1005078 428891 1005080
rect 502412 1005136 502583 1005138
rect 502412 1005080 502522 1005136
rect 502578 1005080 502583 1005136
rect 502412 1005078 502583 1005080
rect 264329 1005075 264395 1005078
rect 269205 1005075 269271 1005078
rect 427537 1005075 427603 1005078
rect 428825 1005075 428891 1005078
rect 502517 1005075 502583 1005078
rect 150893 1005002 150959 1005005
rect 157793 1005002 157859 1005005
rect 208393 1005002 208459 1005005
rect 252829 1005002 252895 1005005
rect 150696 1005000 150959 1005002
rect 150696 1004972 150898 1005000
rect 150666 1004944 150898 1004972
rect 150954 1004944 150959 1005000
rect 150666 1004942 150959 1004944
rect 157596 1005000 157859 1005002
rect 157596 1004944 157798 1005000
rect 157854 1004944 157859 1005000
rect 157596 1004942 157859 1004944
rect 208196 1005000 208459 1005002
rect 208196 1004944 208398 1005000
rect 208454 1004944 208459 1005000
rect 208196 1004942 208459 1004944
rect 252724 1005000 252895 1005002
rect 252724 1004944 252834 1005000
rect 252890 1004944 252895 1005000
rect 252724 1004942 252895 1004944
rect 108021 1004866 108087 1004869
rect 107916 1004864 108087 1004866
rect 107916 1004808 108026 1004864
rect 108082 1004808 108087 1004864
rect 107916 1004806 108087 1004808
rect 108021 1004803 108087 1004806
rect 109677 1004866 109743 1004869
rect 114645 1004866 114711 1004869
rect 109677 1004864 114711 1004866
rect 109677 1004808 109682 1004864
rect 109738 1004808 114650 1004864
rect 114706 1004808 114711 1004864
rect 109677 1004806 114711 1004808
rect 109677 1004803 109743 1004806
rect 114645 1004803 114711 1004806
rect 98269 1004730 98335 1004733
rect 98072 1004728 98335 1004730
rect 98072 1004672 98274 1004728
rect 98330 1004672 98335 1004728
rect 98072 1004670 98335 1004672
rect 98269 1004667 98335 1004670
rect 98637 1004730 98703 1004733
rect 99465 1004730 99531 1004733
rect 98637 1004728 98900 1004730
rect 98637 1004672 98642 1004728
rect 98698 1004672 98900 1004728
rect 99268 1004728 99531 1004730
rect 99268 1004700 99470 1004728
rect 98637 1004670 98900 1004672
rect 99238 1004672 99470 1004700
rect 99526 1004672 99531 1004728
rect 99238 1004670 99531 1004672
rect 98637 1004667 98703 1004670
rect 87822 996372 87828 996436
rect 87892 996434 87898 996436
rect 96521 996434 96587 996437
rect 87892 996432 96587 996434
rect 87892 996376 96526 996432
rect 96582 996376 96587 996432
rect 87892 996374 96587 996376
rect 87892 996372 87898 996374
rect 96521 996371 96587 996374
rect 96429 995890 96495 995893
rect 82770 995888 96495 995890
rect 82770 995832 96434 995888
rect 96490 995832 96495 995888
rect 82770 995830 96495 995832
rect 98502 995890 98562 996132
rect 99238 995890 99298 1004670
rect 99465 1004667 99531 1004670
rect 108849 1004730 108915 1004733
rect 149697 1004730 149763 1004733
rect 108849 1004728 109112 1004730
rect 108849 1004672 108854 1004728
rect 108910 1004672 109112 1004728
rect 108849 1004670 109112 1004672
rect 149500 1004728 149763 1004730
rect 149500 1004672 149702 1004728
rect 149758 1004672 149763 1004728
rect 149500 1004670 149763 1004672
rect 108849 1004667 108915 1004670
rect 149697 1004667 149763 1004670
rect 150065 1004730 150131 1004733
rect 150065 1004728 150328 1004730
rect 150065 1004672 150070 1004728
rect 150126 1004672 150328 1004728
rect 150065 1004670 150328 1004672
rect 150065 1004667 150131 1004670
rect 102777 999834 102843 999837
rect 104341 999834 104407 999837
rect 102777 999832 102948 999834
rect 102777 999776 102782 999832
rect 102838 999776 102948 999832
rect 102777 999774 102948 999776
rect 104341 999832 104604 999834
rect 104341 999776 104346 999832
rect 104402 999776 104604 999832
rect 104341 999774 104604 999776
rect 102777 999771 102843 999774
rect 104341 999771 104407 999774
rect 102317 999698 102383 999701
rect 102317 999696 102580 999698
rect 102317 999640 102322 999696
rect 102378 999640 102580 999696
rect 102317 999638 102580 999640
rect 102317 999635 102383 999638
rect 101949 999562 102015 999565
rect 101949 999560 102212 999562
rect 101949 999504 101954 999560
rect 102010 999504 102212 999560
rect 101949 999502 102212 999504
rect 101949 999499 102015 999502
rect 103145 999426 103211 999429
rect 103145 999424 103408 999426
rect 103145 999368 103150 999424
rect 103206 999368 103408 999424
rect 103145 999366 103408 999368
rect 103145 999363 103211 999366
rect 107653 997250 107719 997253
rect 107456 997248 107719 997250
rect 107456 997192 107658 997248
rect 107714 997192 107719 997248
rect 107456 997190 107719 997192
rect 107653 997187 107719 997190
rect 115933 997250 115999 997253
rect 144269 997250 144335 997253
rect 115933 997248 144335 997250
rect 115933 997192 115938 997248
rect 115994 997192 144274 997248
rect 144330 997192 144335 997248
rect 115933 997190 144335 997192
rect 115933 997187 115999 997190
rect 144269 997187 144335 997190
rect 101121 996434 101187 996437
rect 148869 996434 148935 996437
rect 101121 996432 101292 996434
rect 101121 996376 101126 996432
rect 101182 996376 101292 996432
rect 101121 996374 101292 996376
rect 142846 996432 148935 996434
rect 142846 996376 148874 996432
rect 148930 996376 148935 996432
rect 142846 996374 148935 996376
rect 101121 996371 101187 996374
rect 100293 996162 100359 996165
rect 100753 996162 100819 996165
rect 101489 996162 101555 996165
rect 108481 996162 108547 996165
rect 108849 996162 108915 996165
rect 100293 996160 100556 996162
rect 98502 995830 99298 995890
rect 81617 995482 81683 995485
rect 82770 995482 82830 995830
rect 96429 995827 96495 995830
rect 86585 995754 86651 995757
rect 99698 995754 99758 996132
rect 86585 995752 99758 995754
rect 86585 995696 86590 995752
rect 86646 995696 99758 995752
rect 86585 995694 99758 995696
rect 86585 995691 86651 995694
rect 87781 995620 87847 995621
rect 87781 995618 87828 995620
rect 87736 995616 87828 995618
rect 87736 995560 87786 995616
rect 87736 995558 87828 995560
rect 87781 995556 87828 995558
rect 87892 995556 87898 995620
rect 100066 995618 100126 996132
rect 100293 996104 100298 996160
rect 100354 996104 100556 996160
rect 100293 996102 100556 996104
rect 100753 996160 100924 996162
rect 100753 996104 100758 996160
rect 100814 996104 100924 996160
rect 100753 996102 100924 996104
rect 101489 996160 101752 996162
rect 101489 996104 101494 996160
rect 101550 996104 101752 996160
rect 108284 996160 108547 996162
rect 101489 996102 101752 996104
rect 100293 996099 100359 996102
rect 100753 996099 100819 996102
rect 101489 996099 101555 996102
rect 92614 995558 100126 995618
rect 100201 995618 100267 995621
rect 103746 995618 103806 996132
rect 104206 995621 104266 996132
rect 100201 995616 103806 995618
rect 100201 995560 100206 995616
rect 100262 995560 103806 995616
rect 100201 995558 103806 995560
rect 104157 995616 104266 995621
rect 104157 995560 104162 995616
rect 104218 995560 104266 995616
rect 104157 995558 104266 995560
rect 104341 995618 104407 995621
rect 104942 995618 105002 996132
rect 104341 995616 105002 995618
rect 104341 995560 104346 995616
rect 104402 995560 105002 995616
rect 104341 995558 105002 995560
rect 105862 995618 105922 996132
rect 106598 995754 106658 996132
rect 107058 995890 107118 996132
rect 108284 996104 108486 996160
rect 108542 996104 108547 996160
rect 108284 996102 108547 996104
rect 108652 996160 108915 996162
rect 108652 996104 108854 996160
rect 108910 996104 108915 996160
rect 108652 996102 108915 996104
rect 108481 996099 108547 996102
rect 108849 996099 108915 996102
rect 110413 995890 110479 995893
rect 107058 995888 110479 995890
rect 107058 995832 110418 995888
rect 110474 995832 110479 995888
rect 107058 995830 110479 995832
rect 110413 995827 110479 995830
rect 142846 995757 142906 996374
rect 148869 996371 148935 996374
rect 149838 995890 149898 996132
rect 150666 995890 150726 1004942
rect 150893 1004939 150959 1004942
rect 157793 1004939 157859 1004942
rect 208393 1004939 208459 1004942
rect 252829 1004939 252895 1004942
rect 253289 1005002 253355 1005005
rect 260649 1005002 260715 1005005
rect 262673 1005002 262739 1005005
rect 253289 1005000 253460 1005002
rect 253289 1004944 253294 1005000
rect 253350 1004944 253460 1005000
rect 253289 1004942 253460 1004944
rect 260452 1005000 260715 1005002
rect 260452 1004944 260654 1005000
rect 260710 1004944 260715 1005000
rect 260452 1004942 260715 1004944
rect 262476 1005000 262739 1005002
rect 262476 1004944 262678 1005000
rect 262734 1004944 262739 1005000
rect 262476 1004942 262739 1004944
rect 253289 1004939 253355 1004942
rect 260649 1004939 260715 1004942
rect 262673 1004939 262739 1004942
rect 264329 1005002 264395 1005005
rect 267825 1005002 267891 1005005
rect 264329 1005000 267891 1005002
rect 264329 1004944 264334 1005000
rect 264390 1004944 267830 1005000
rect 267886 1004944 267891 1005000
rect 264329 1004942 267891 1004944
rect 264329 1004939 264395 1004942
rect 267825 1004939 267891 1004942
rect 350257 1005002 350323 1005005
rect 353661 1005002 353727 1005005
rect 358169 1005002 358235 1005005
rect 425513 1005002 425579 1005005
rect 426801 1005002 426867 1005005
rect 504173 1005002 504239 1005005
rect 350257 1005000 353727 1005002
rect 350257 1004944 350262 1005000
rect 350318 1004944 353666 1005000
rect 353722 1004944 353727 1005000
rect 350257 1004942 353727 1004944
rect 357972 1005000 358235 1005002
rect 357972 1004944 358174 1005000
rect 358230 1004944 358235 1005000
rect 357972 1004942 358235 1004944
rect 425316 1005000 425579 1005002
rect 425316 1004944 425518 1005000
rect 425574 1004944 425579 1005000
rect 425316 1004942 425579 1004944
rect 426604 1005000 426867 1005002
rect 426604 1004944 426806 1005000
rect 426862 1004944 426867 1005000
rect 426604 1004942 426867 1004944
rect 503976 1005000 504239 1005002
rect 503976 1004944 504178 1005000
rect 504234 1004944 504239 1005000
rect 503976 1004942 504239 1004944
rect 350257 1004939 350323 1004942
rect 353661 1004939 353727 1004942
rect 358169 1004939 358235 1004942
rect 425513 1004939 425579 1004942
rect 426801 1004939 426867 1004942
rect 504173 1004939 504239 1004942
rect 546309 1005002 546375 1005005
rect 549437 1005002 549503 1005005
rect 552749 1005002 552815 1005005
rect 546309 1005000 549503 1005002
rect 546309 1004944 546314 1005000
rect 546370 1004944 549442 1005000
rect 549498 1004944 549503 1005000
rect 546309 1004942 549503 1004944
rect 552552 1005000 552815 1005002
rect 552552 1004944 552754 1005000
rect 552810 1004944 552815 1005000
rect 552552 1004942 552815 1004944
rect 546309 1004939 546375 1004942
rect 549437 1004939 549503 1004942
rect 552749 1004939 552815 1004942
rect 156965 1004866 157031 1004869
rect 261845 1004866 261911 1004869
rect 269021 1004866 269087 1004869
rect 423489 1004866 423555 1004869
rect 427169 1004866 427235 1004869
rect 553117 1004866 553183 1004869
rect 156860 1004864 157031 1004866
rect 156860 1004808 156970 1004864
rect 157026 1004808 157031 1004864
rect 156860 1004806 157031 1004808
rect 261648 1004864 261911 1004866
rect 261648 1004808 261850 1004864
rect 261906 1004808 261911 1004864
rect 261648 1004806 261911 1004808
rect 263764 1004864 269087 1004866
rect 263764 1004808 269026 1004864
rect 269082 1004808 269087 1004864
rect 263764 1004806 269087 1004808
rect 423292 1004864 423555 1004866
rect 423292 1004808 423494 1004864
rect 423550 1004808 423555 1004864
rect 423292 1004806 423555 1004808
rect 426972 1004864 427235 1004866
rect 426972 1004808 427174 1004864
rect 427230 1004808 427235 1004864
rect 426972 1004806 427235 1004808
rect 552920 1004864 553183 1004866
rect 552920 1004808 553122 1004864
rect 553178 1004808 553183 1004864
rect 552920 1004806 553183 1004808
rect 156965 1004803 157031 1004806
rect 261845 1004803 261911 1004806
rect 269021 1004803 269087 1004806
rect 423489 1004803 423555 1004806
rect 427169 1004803 427235 1004806
rect 553117 1004803 553183 1004806
rect 154941 1004730 155007 1004733
rect 159449 1004730 159515 1004733
rect 154941 1004728 155204 1004730
rect 154941 1004672 154946 1004728
rect 155002 1004672 155204 1004728
rect 154941 1004670 155204 1004672
rect 159252 1004728 159515 1004730
rect 159252 1004672 159454 1004728
rect 159510 1004672 159515 1004728
rect 159252 1004670 159515 1004672
rect 154941 1004667 155007 1004670
rect 159449 1004667 159515 1004670
rect 160645 1004730 160711 1004733
rect 205173 1004730 205239 1004733
rect 205909 1004730 205975 1004733
rect 206369 1004730 206435 1004733
rect 218053 1004730 218119 1004733
rect 252461 1004730 252527 1004733
rect 160645 1004728 160908 1004730
rect 160645 1004672 160650 1004728
rect 160706 1004672 160908 1004728
rect 160645 1004670 160908 1004672
rect 205173 1004728 205344 1004730
rect 205173 1004672 205178 1004728
rect 205234 1004672 205344 1004728
rect 205173 1004670 205344 1004672
rect 205909 1004728 206172 1004730
rect 205909 1004672 205914 1004728
rect 205970 1004672 206172 1004728
rect 205909 1004670 206172 1004672
rect 206369 1004728 206540 1004730
rect 206369 1004672 206374 1004728
rect 206430 1004672 206540 1004728
rect 206369 1004670 206540 1004672
rect 212336 1004728 218119 1004730
rect 212336 1004672 218058 1004728
rect 218114 1004672 218119 1004728
rect 212336 1004670 218119 1004672
rect 252264 1004728 252527 1004730
rect 252264 1004672 252466 1004728
rect 252522 1004672 252527 1004728
rect 252264 1004670 252527 1004672
rect 160645 1004667 160711 1004670
rect 205173 1004667 205239 1004670
rect 205909 1004667 205975 1004670
rect 206369 1004667 206435 1004670
rect 218053 1004667 218119 1004670
rect 252461 1004667 252527 1004670
rect 252829 1004730 252895 1004733
rect 261477 1004730 261543 1004733
rect 262213 1004730 262279 1004733
rect 263501 1004730 263567 1004733
rect 252829 1004728 253092 1004730
rect 252829 1004672 252834 1004728
rect 252890 1004672 253092 1004728
rect 252829 1004670 253092 1004672
rect 261280 1004728 261543 1004730
rect 261280 1004672 261482 1004728
rect 261538 1004672 261543 1004728
rect 261280 1004670 261543 1004672
rect 262108 1004728 262279 1004730
rect 262108 1004672 262218 1004728
rect 262274 1004672 262279 1004728
rect 262108 1004670 262279 1004672
rect 263304 1004728 263567 1004730
rect 263304 1004672 263506 1004728
rect 263562 1004672 263567 1004728
rect 263304 1004670 263567 1004672
rect 252829 1004667 252895 1004670
rect 261477 1004667 261543 1004670
rect 262213 1004667 262279 1004670
rect 263501 1004667 263567 1004670
rect 263869 1004730 263935 1004733
rect 267733 1004730 267799 1004733
rect 304073 1004730 304139 1004733
rect 263869 1004728 267799 1004730
rect 263869 1004672 263874 1004728
rect 263930 1004672 267738 1004728
rect 267794 1004672 267799 1004728
rect 263869 1004670 267799 1004672
rect 303876 1004728 304139 1004730
rect 303876 1004672 304078 1004728
rect 304134 1004672 304139 1004728
rect 303876 1004670 304139 1004672
rect 263869 1004667 263935 1004670
rect 267733 1004667 267799 1004670
rect 304073 1004667 304139 1004670
rect 304441 1004730 304507 1004733
rect 315113 1004730 315179 1004733
rect 321461 1004730 321527 1004733
rect 354489 1004730 354555 1004733
rect 304441 1004728 304704 1004730
rect 304441 1004672 304446 1004728
rect 304502 1004672 304704 1004728
rect 304441 1004670 304704 1004672
rect 314916 1004728 315179 1004730
rect 314916 1004672 315118 1004728
rect 315174 1004672 315179 1004728
rect 314916 1004670 315179 1004672
rect 315284 1004728 321527 1004730
rect 315284 1004672 321466 1004728
rect 321522 1004672 321527 1004728
rect 315284 1004670 321527 1004672
rect 354292 1004728 354555 1004730
rect 354292 1004672 354494 1004728
rect 354550 1004672 354555 1004728
rect 354292 1004670 354555 1004672
rect 304441 1004667 304507 1004670
rect 315113 1004667 315179 1004670
rect 321461 1004667 321527 1004670
rect 354489 1004667 354555 1004670
rect 354857 1004730 354923 1004733
rect 358537 1004730 358603 1004733
rect 359733 1004730 359799 1004733
rect 422293 1004730 422359 1004733
rect 354857 1004728 355120 1004730
rect 354857 1004672 354862 1004728
rect 354918 1004672 355120 1004728
rect 354857 1004670 355120 1004672
rect 358340 1004728 358603 1004730
rect 358340 1004672 358542 1004728
rect 358598 1004672 358603 1004728
rect 358340 1004670 358603 1004672
rect 359628 1004728 359799 1004730
rect 359628 1004672 359738 1004728
rect 359794 1004672 359799 1004728
rect 359628 1004670 359799 1004672
rect 422096 1004728 422359 1004730
rect 422096 1004672 422298 1004728
rect 422354 1004672 422359 1004728
rect 422096 1004670 422359 1004672
rect 354857 1004667 354923 1004670
rect 358537 1004667 358603 1004670
rect 359733 1004667 359799 1004670
rect 422293 1004667 422359 1004670
rect 422661 1004730 422727 1004733
rect 424685 1004730 424751 1004733
rect 499297 1004730 499363 1004733
rect 422661 1004728 422924 1004730
rect 422661 1004672 422666 1004728
rect 422722 1004672 422924 1004728
rect 422661 1004670 422924 1004672
rect 424580 1004728 424751 1004730
rect 424580 1004672 424690 1004728
rect 424746 1004672 424751 1004728
rect 424580 1004670 424751 1004672
rect 499100 1004728 499363 1004730
rect 499100 1004672 499302 1004728
rect 499358 1004672 499363 1004728
rect 499100 1004670 499363 1004672
rect 422661 1004667 422727 1004670
rect 424685 1004667 424751 1004670
rect 499297 1004667 499363 1004670
rect 499665 1004730 499731 1004733
rect 501689 1004730 501755 1004733
rect 502149 1004730 502215 1004733
rect 550265 1004730 550331 1004733
rect 499665 1004728 499928 1004730
rect 499665 1004672 499670 1004728
rect 499726 1004672 499928 1004728
rect 499665 1004670 499928 1004672
rect 501492 1004728 501755 1004730
rect 501492 1004672 501694 1004728
rect 501750 1004672 501755 1004728
rect 501492 1004670 501755 1004672
rect 501952 1004728 502215 1004730
rect 501952 1004672 502154 1004728
rect 502210 1004672 502215 1004728
rect 501952 1004670 502215 1004672
rect 550068 1004728 550331 1004730
rect 550068 1004672 550270 1004728
rect 550326 1004672 550331 1004728
rect 550068 1004670 550331 1004672
rect 499665 1004667 499731 1004670
rect 501689 1004667 501755 1004670
rect 502149 1004667 502215 1004670
rect 550265 1004667 550331 1004670
rect 550633 1004730 550699 1004733
rect 551921 1004730 551987 1004733
rect 554313 1004730 554379 1004733
rect 561305 1004730 561371 1004733
rect 567285 1004730 567351 1004733
rect 550633 1004728 550896 1004730
rect 550633 1004672 550638 1004728
rect 550694 1004672 550896 1004728
rect 550633 1004670 550896 1004672
rect 551724 1004728 551987 1004730
rect 551724 1004672 551926 1004728
rect 551982 1004672 551987 1004728
rect 551724 1004670 551987 1004672
rect 554116 1004728 554379 1004730
rect 554116 1004672 554318 1004728
rect 554374 1004672 554379 1004728
rect 554116 1004670 554379 1004672
rect 561108 1004728 561371 1004730
rect 561108 1004672 561310 1004728
rect 561366 1004672 561371 1004728
rect 561108 1004670 561371 1004672
rect 561476 1004728 567351 1004730
rect 561476 1004672 567290 1004728
rect 567346 1004672 567351 1004728
rect 561476 1004670 567351 1004672
rect 550633 1004667 550699 1004670
rect 551921 1004667 551987 1004670
rect 554313 1004667 554379 1004670
rect 561305 1004667 561371 1004670
rect 567285 1004667 567351 1004670
rect 553945 1003914 554011 1003917
rect 553748 1003912 554011 1003914
rect 553748 1003856 553950 1003912
rect 554006 1003856 554011 1003912
rect 553748 1003854 554011 1003856
rect 553945 1003851 554011 1003854
rect 555509 1003370 555575 1003373
rect 555404 1003368 555575 1003370
rect 555404 1003312 555514 1003368
rect 555570 1003312 555575 1003368
rect 555404 1003310 555575 1003312
rect 555509 1003307 555575 1003310
rect 554773 1003234 554839 1003237
rect 554576 1003232 554839 1003234
rect 554576 1003176 554778 1003232
rect 554834 1003176 554839 1003232
rect 554576 1003174 554839 1003176
rect 554773 1003171 554839 1003174
rect 360561 1000786 360627 1000789
rect 360364 1000784 360627 1000786
rect 360364 1000728 360566 1000784
rect 360622 1000728 360627 1000784
rect 360364 1000726 360627 1000728
rect 360561 1000723 360627 1000726
rect 361389 1000650 361455 1000653
rect 427997 1000650 428063 1000653
rect 361192 1000648 361455 1000650
rect 361192 1000592 361394 1000648
rect 361450 1000592 361455 1000648
rect 361192 1000590 361455 1000592
rect 427800 1000648 428063 1000650
rect 427800 1000592 428002 1000648
rect 428058 1000592 428063 1000648
rect 427800 1000590 428063 1000592
rect 361389 1000587 361455 1000590
rect 427997 1000587 428063 1000590
rect 358905 1000514 358971 1000517
rect 426341 1000514 426407 1000517
rect 358800 1000512 358971 1000514
rect 358800 1000456 358910 1000512
rect 358966 1000456 358971 1000512
rect 358800 1000454 358971 1000456
rect 426144 1000512 426407 1000514
rect 426144 1000456 426346 1000512
rect 426402 1000456 426407 1000512
rect 426144 1000454 426407 1000456
rect 358905 1000451 358971 1000454
rect 426341 1000451 426407 1000454
rect 258625 999970 258691 999973
rect 503345 999970 503411 999973
rect 258625 999968 258796 999970
rect 258625 999912 258630 999968
rect 258686 999912 258796 999968
rect 258625 999910 258796 999912
rect 503148 999968 503411 999970
rect 503148 999912 503350 999968
rect 503406 999912 503411 999968
rect 503148 999910 503411 999912
rect 258625 999907 258691 999910
rect 503345 999907 503411 999910
rect 516041 999970 516107 999973
rect 524045 999970 524111 999973
rect 516041 999968 524111 999970
rect 516041 999912 516046 999968
rect 516102 999912 524050 999968
rect 524106 999912 524111 999968
rect 516041 999910 524111 999912
rect 516041 999907 516107 999910
rect 524045 999907 524111 999910
rect 256969 999834 257035 999837
rect 257337 999834 257403 999837
rect 311433 999834 311499 999837
rect 312169 999834 312235 999837
rect 430849 999834 430915 999837
rect 508681 999834 508747 999837
rect 560845 999834 560911 999837
rect 256969 999832 257140 999834
rect 256969 999776 256974 999832
rect 257030 999776 257140 999832
rect 256969 999774 257140 999776
rect 257337 999832 257600 999834
rect 257337 999776 257342 999832
rect 257398 999776 257600 999832
rect 257337 999774 257600 999776
rect 311236 999832 311499 999834
rect 311236 999776 311438 999832
rect 311494 999776 311499 999832
rect 311236 999774 311499 999776
rect 312064 999832 312235 999834
rect 312064 999776 312174 999832
rect 312230 999776 312235 999832
rect 312064 999774 312235 999776
rect 430652 999832 430915 999834
rect 430652 999776 430854 999832
rect 430910 999776 430915 999832
rect 430652 999774 430915 999776
rect 508484 999832 508747 999834
rect 508484 999776 508686 999832
rect 508742 999776 508747 999832
rect 508484 999774 508747 999776
rect 560740 999832 560911 999834
rect 560740 999776 560850 999832
rect 560906 999776 560911 999832
rect 560740 999774 560911 999776
rect 256969 999771 257035 999774
rect 257337 999771 257403 999774
rect 311433 999771 311499 999774
rect 312169 999771 312235 999774
rect 430849 999771 430915 999774
rect 508681 999771 508747 999774
rect 560845 999771 560911 999774
rect 205541 999698 205607 999701
rect 257797 999698 257863 999701
rect 310145 999698 310211 999701
rect 313825 999698 313891 999701
rect 429193 999698 429259 999701
rect 431677 999698 431743 999701
rect 506197 999698 506263 999701
rect 507025 999698 507091 999701
rect 560477 999698 560543 999701
rect 205541 999696 205804 999698
rect 205541 999640 205546 999696
rect 205602 999640 205804 999696
rect 205541 999638 205804 999640
rect 257797 999696 257968 999698
rect 257797 999640 257802 999696
rect 257858 999640 257968 999696
rect 257797 999638 257968 999640
rect 309948 999696 310211 999698
rect 309948 999640 310150 999696
rect 310206 999640 310211 999696
rect 309948 999638 310211 999640
rect 313628 999696 313891 999698
rect 313628 999640 313830 999696
rect 313886 999640 313891 999696
rect 313628 999638 313891 999640
rect 428996 999696 429259 999698
rect 428996 999640 429198 999696
rect 429254 999640 429259 999696
rect 428996 999638 429259 999640
rect 431480 999696 431743 999698
rect 431480 999640 431682 999696
rect 431738 999640 431743 999696
rect 431480 999638 431743 999640
rect 506000 999696 506263 999698
rect 506000 999640 506202 999696
rect 506258 999640 506263 999696
rect 506000 999638 506263 999640
rect 506828 999696 507091 999698
rect 506828 999640 507030 999696
rect 507086 999640 507091 999696
rect 506828 999638 507091 999640
rect 560280 999696 560543 999698
rect 560280 999640 560482 999696
rect 560538 999640 560543 999696
rect 560280 999638 560543 999640
rect 205541 999635 205607 999638
rect 257797 999635 257863 999638
rect 310145 999635 310211 999638
rect 313825 999635 313891 999638
rect 429193 999635 429259 999638
rect 431677 999635 431743 999638
rect 506197 999635 506263 999638
rect 507025 999635 507091 999638
rect 560477 999635 560543 999638
rect 155769 999562 155835 999565
rect 159081 999562 159147 999565
rect 155572 999560 155835 999562
rect 155572 999504 155774 999560
rect 155830 999504 155835 999560
rect 155572 999502 155835 999504
rect 158884 999560 159147 999562
rect 158884 999504 159086 999560
rect 159142 999504 159147 999560
rect 158884 999502 159147 999504
rect 155769 999499 155835 999502
rect 159081 999499 159147 999502
rect 203517 999562 203583 999565
rect 203885 999562 203951 999565
rect 312997 999562 313063 999565
rect 314653 999562 314719 999565
rect 430021 999562 430087 999565
rect 431217 999562 431283 999565
rect 507853 999562 507919 999565
rect 508221 999562 508287 999565
rect 203517 999560 203780 999562
rect 203517 999504 203522 999560
rect 203578 999504 203780 999560
rect 203517 999502 203780 999504
rect 203885 999560 204148 999562
rect 203885 999504 203890 999560
rect 203946 999504 204148 999560
rect 203885 999502 204148 999504
rect 312892 999560 313063 999562
rect 312892 999504 313002 999560
rect 313058 999504 313063 999560
rect 312892 999502 313063 999504
rect 314548 999560 314719 999562
rect 314548 999504 314658 999560
rect 314714 999504 314719 999560
rect 314548 999502 314719 999504
rect 429824 999560 430087 999562
rect 429824 999504 430026 999560
rect 430082 999504 430087 999560
rect 429824 999502 430087 999504
rect 431020 999560 431283 999562
rect 431020 999504 431222 999560
rect 431278 999504 431283 999560
rect 431020 999502 431283 999504
rect 507656 999560 507919 999562
rect 507656 999504 507858 999560
rect 507914 999504 507919 999560
rect 507656 999502 507919 999504
rect 508116 999560 508287 999562
rect 508116 999504 508226 999560
rect 508282 999504 508287 999560
rect 508116 999502 508287 999504
rect 203517 999499 203583 999502
rect 203885 999499 203951 999502
rect 312997 999499 313063 999502
rect 314653 999499 314719 999502
rect 430021 999499 430087 999502
rect 431217 999499 431283 999502
rect 507853 999499 507919 999502
rect 508221 999499 508287 999502
rect 202321 999426 202387 999429
rect 204713 999426 204779 999429
rect 309777 999426 309843 999429
rect 312629 999426 312695 999429
rect 429653 999426 429719 999429
rect 432505 999426 432571 999429
rect 500493 999426 500559 999429
rect 506565 999426 506631 999429
rect 509049 999426 509115 999429
rect 202321 999424 202492 999426
rect 202321 999368 202326 999424
rect 202382 999368 202492 999424
rect 202321 999366 202492 999368
rect 204713 999424 204976 999426
rect 204713 999368 204718 999424
rect 204774 999368 204976 999424
rect 204713 999366 204976 999368
rect 309580 999424 309843 999426
rect 309580 999368 309782 999424
rect 309838 999368 309843 999424
rect 309580 999366 309843 999368
rect 312432 999424 312695 999426
rect 312432 999368 312634 999424
rect 312690 999368 312695 999424
rect 312432 999366 312695 999368
rect 429456 999424 429719 999426
rect 429456 999368 429658 999424
rect 429714 999368 429719 999424
rect 429456 999366 429719 999368
rect 432308 999424 432571 999426
rect 432308 999368 432510 999424
rect 432566 999368 432571 999424
rect 432308 999366 432571 999368
rect 500296 999424 500559 999426
rect 500296 999368 500498 999424
rect 500554 999368 500559 999424
rect 500296 999366 500559 999368
rect 506460 999424 506631 999426
rect 506460 999368 506570 999424
rect 506626 999368 506631 999424
rect 506460 999366 506631 999368
rect 508852 999424 509115 999426
rect 508852 999368 509054 999424
rect 509110 999368 509115 999424
rect 508852 999366 509115 999368
rect 202321 999363 202387 999366
rect 204713 999363 204779 999366
rect 309777 999363 309843 999366
rect 312629 999363 312695 999366
rect 429653 999363 429719 999366
rect 432505 999363 432571 999366
rect 500493 999363 500559 999366
rect 506565 999363 506631 999366
rect 509049 999363 509115 999366
rect 202689 999290 202755 999293
rect 204345 999290 204411 999293
rect 256509 999290 256575 999293
rect 310973 999290 311039 999293
rect 311801 999290 311867 999293
rect 357341 999290 357407 999293
rect 432045 999290 432111 999293
rect 432873 999290 432939 999293
rect 500861 999290 500927 999293
rect 507393 999290 507459 999293
rect 509509 999290 509575 999293
rect 202689 999288 202952 999290
rect 202689 999232 202694 999288
rect 202750 999232 202952 999288
rect 202689 999230 202952 999232
rect 204345 999288 204516 999290
rect 204345 999232 204350 999288
rect 204406 999232 204516 999288
rect 204345 999230 204516 999232
rect 256509 999288 256772 999290
rect 256509 999232 256514 999288
rect 256570 999232 256772 999288
rect 256509 999230 256772 999232
rect 310868 999288 311039 999290
rect 310868 999232 310978 999288
rect 311034 999232 311039 999288
rect 310868 999230 311039 999232
rect 311604 999288 311867 999290
rect 311604 999232 311806 999288
rect 311862 999232 311867 999288
rect 311604 999230 311867 999232
rect 357144 999288 357407 999290
rect 357144 999232 357346 999288
rect 357402 999232 357407 999288
rect 357144 999230 357407 999232
rect 431940 999288 432111 999290
rect 431940 999232 432050 999288
rect 432106 999232 432111 999288
rect 431940 999230 432111 999232
rect 432676 999288 432939 999290
rect 432676 999232 432878 999288
rect 432934 999232 432939 999288
rect 432676 999230 432939 999232
rect 500756 999288 500927 999290
rect 500756 999232 500866 999288
rect 500922 999232 500927 999288
rect 500756 999230 500927 999232
rect 507196 999288 507459 999290
rect 507196 999232 507398 999288
rect 507454 999232 507459 999288
rect 507196 999230 507459 999232
rect 509312 999288 509575 999290
rect 509312 999232 509514 999288
rect 509570 999232 509575 999288
rect 509312 999230 509575 999232
rect 202689 999227 202755 999230
rect 204345 999227 204411 999230
rect 256509 999227 256575 999230
rect 310973 999227 311039 999230
rect 311801 999227 311867 999230
rect 357341 999227 357407 999230
rect 432045 999227 432111 999230
rect 432873 999227 432939 999230
rect 500861 999227 500927 999230
rect 507393 999227 507459 999230
rect 509509 999227 509575 999230
rect 158253 999154 158319 999157
rect 203057 999154 203123 999157
rect 258533 999154 258599 999157
rect 314285 999154 314351 999157
rect 357709 999154 357775 999157
rect 430389 999154 430455 999157
rect 437749 999154 437815 999157
rect 509877 999154 509943 999157
rect 515029 999154 515095 999157
rect 158253 999152 158516 999154
rect 158253 999096 158258 999152
rect 158314 999096 158516 999152
rect 158253 999094 158516 999096
rect 203057 999152 203320 999154
rect 203057 999096 203062 999152
rect 203118 999096 203320 999152
rect 203057 999094 203320 999096
rect 258428 999152 258599 999154
rect 258428 999096 258538 999152
rect 258594 999096 258599 999152
rect 258428 999094 258599 999096
rect 314088 999152 314351 999154
rect 314088 999096 314290 999152
rect 314346 999096 314351 999152
rect 314088 999094 314351 999096
rect 357604 999152 357775 999154
rect 357604 999096 357714 999152
rect 357770 999096 357775 999152
rect 357604 999094 357775 999096
rect 430284 999152 430455 999154
rect 430284 999096 430394 999152
rect 430450 999096 430455 999152
rect 430284 999094 430455 999096
rect 433136 999152 437815 999154
rect 433136 999096 437754 999152
rect 437810 999096 437815 999152
rect 433136 999094 437815 999096
rect 509680 999152 509943 999154
rect 509680 999096 509882 999152
rect 509938 999096 509943 999152
rect 509680 999094 509943 999096
rect 510140 999152 515095 999154
rect 510140 999096 515034 999152
rect 515090 999096 515095 999152
rect 510140 999094 515095 999096
rect 158253 999091 158319 999094
rect 203057 999091 203123 999094
rect 258533 999091 258599 999094
rect 314285 999091 314351 999094
rect 357709 999091 357775 999094
rect 430389 999091 430455 999094
rect 437749 999091 437815 999094
rect 509877 999091 509943 999094
rect 515029 999091 515095 999094
rect 519077 999154 519143 999157
rect 523769 999154 523835 999157
rect 552289 999154 552355 999157
rect 519077 999152 523835 999154
rect 519077 999096 519082 999152
rect 519138 999096 523774 999152
rect 523830 999096 523835 999152
rect 519077 999094 523835 999096
rect 552092 999152 552355 999154
rect 552092 999096 552294 999152
rect 552350 999096 552355 999152
rect 552092 999094 552355 999096
rect 519077 999091 519143 999094
rect 523769 999091 523835 999094
rect 552289 999091 552355 999094
rect 156137 997794 156203 997797
rect 501321 997794 501387 997797
rect 553485 997794 553551 997797
rect 156137 997792 156400 997794
rect 156137 997736 156142 997792
rect 156198 997736 156400 997792
rect 156137 997734 156400 997736
rect 501124 997792 501387 997794
rect 501124 997736 501326 997792
rect 501382 997736 501387 997792
rect 501124 997734 501387 997736
rect 553380 997792 553551 997794
rect 553380 997736 553490 997792
rect 553546 997736 553551 997792
rect 553380 997734 553551 997736
rect 156137 997731 156203 997734
rect 501321 997731 501387 997734
rect 553485 997731 553551 997734
rect 556337 997658 556403 997661
rect 556232 997656 556403 997658
rect 556232 997600 556342 997656
rect 556398 997600 556403 997656
rect 556232 997598 556403 997600
rect 556337 997595 556403 997598
rect 557165 997522 557231 997525
rect 557060 997520 557231 997522
rect 557060 997464 557170 997520
rect 557226 997464 557231 997520
rect 557060 997462 557231 997464
rect 557165 997459 557231 997462
rect 187734 997188 187740 997252
rect 187804 997250 187810 997252
rect 195145 997250 195211 997253
rect 210417 997250 210483 997253
rect 187804 997248 195211 997250
rect 187804 997192 195150 997248
rect 195206 997192 195211 997248
rect 187804 997190 195211 997192
rect 210220 997248 210483 997250
rect 210220 997192 210422 997248
rect 210478 997192 210483 997248
rect 210220 997190 210483 997192
rect 187804 997188 187810 997190
rect 195145 997187 195211 997190
rect 210417 997187 210483 997190
rect 215293 997250 215359 997253
rect 246573 997250 246639 997253
rect 215293 997248 246639 997250
rect 215293 997192 215298 997248
rect 215354 997192 246578 997248
rect 246634 997192 246639 997248
rect 215293 997190 246639 997192
rect 215293 997187 215359 997190
rect 246573 997187 246639 997190
rect 266261 997250 266327 997253
rect 298737 997250 298803 997253
rect 363413 997250 363479 997253
rect 266261 997248 298803 997250
rect 266261 997192 266266 997248
rect 266322 997192 298742 997248
rect 298798 997192 298803 997248
rect 266261 997190 298803 997192
rect 363308 997248 363479 997250
rect 363308 997192 363418 997248
rect 363474 997192 363479 997248
rect 363308 997190 363479 997192
rect 266261 997187 266327 997190
rect 298737 997187 298803 997190
rect 363413 997187 363479 997190
rect 367093 997250 367159 997253
rect 399937 997250 400003 997253
rect 367093 997248 400003 997250
rect 367093 997192 367098 997248
rect 367154 997192 399942 997248
rect 399998 997192 400003 997248
rect 367093 997190 400003 997192
rect 367093 997187 367159 997190
rect 399937 997187 400003 997190
rect 162853 997114 162919 997117
rect 195329 997114 195395 997117
rect 162853 997112 195395 997114
rect 162853 997056 162858 997112
rect 162914 997056 195334 997112
rect 195390 997056 195395 997112
rect 162853 997054 195395 997056
rect 162853 997051 162919 997054
rect 195329 997051 195395 997054
rect 438117 997114 438183 997117
rect 489453 997114 489519 997117
rect 438117 997112 489519 997114
rect 438117 997056 438122 997112
rect 438178 997056 489458 997112
rect 489514 997056 489519 997112
rect 438117 997054 489519 997056
rect 438117 997051 438183 997054
rect 489453 997051 489519 997054
rect 523769 996570 523835 996573
rect 523769 996568 532250 996570
rect 523769 996512 523774 996568
rect 523830 996512 532250 996568
rect 523769 996510 532250 996512
rect 523769 996507 523835 996510
rect 151721 996434 151787 996437
rect 154113 996434 154179 996437
rect 381721 996434 381787 996437
rect 461025 996434 461091 996437
rect 476430 996434 476436 996436
rect 151721 996432 151892 996434
rect 151721 996376 151726 996432
rect 151782 996376 151892 996432
rect 151721 996374 151892 996376
rect 154113 996432 154376 996434
rect 154113 996376 154118 996432
rect 154174 996376 154376 996432
rect 154113 996374 154376 996376
rect 381721 996432 388178 996434
rect 381721 996376 381726 996432
rect 381782 996376 388178 996432
rect 381721 996374 388178 996376
rect 151721 996371 151787 996374
rect 154113 996371 154179 996374
rect 381721 996371 381787 996374
rect 153745 996298 153811 996301
rect 308121 996298 308187 996301
rect 308949 996298 309015 996301
rect 365437 996298 365503 996301
rect 153745 996296 153916 996298
rect 153745 996240 153750 996296
rect 153806 996240 153916 996296
rect 153745 996238 153916 996240
rect 308121 996296 308384 996298
rect 308121 996240 308126 996296
rect 308182 996240 308384 996296
rect 308121 996238 308384 996240
rect 308949 996296 309212 996298
rect 308949 996240 308954 996296
rect 309010 996240 309212 996296
rect 308949 996238 309212 996240
rect 365332 996296 365503 996298
rect 365332 996240 365442 996296
rect 365498 996240 365503 996296
rect 365332 996238 365503 996240
rect 153745 996235 153811 996238
rect 308121 996235 308187 996238
rect 308949 996235 309015 996238
rect 365437 996235 365503 996238
rect 150893 996162 150959 996165
rect 151261 996162 151327 996165
rect 152549 996162 152615 996165
rect 152917 996162 152983 996165
rect 153377 996162 153443 996165
rect 154573 996162 154639 996165
rect 156965 996162 157031 996165
rect 157793 996162 157859 996165
rect 159449 996162 159515 996165
rect 208761 996162 208827 996165
rect 209589 996162 209655 996165
rect 211245 996162 211311 996165
rect 150893 996160 151156 996162
rect 150893 996104 150898 996160
rect 150954 996104 151156 996160
rect 150893 996102 151156 996104
rect 151261 996160 151524 996162
rect 151261 996104 151266 996160
rect 151322 996104 151524 996160
rect 152549 996160 152720 996162
rect 151261 996102 151524 996104
rect 150893 996099 150959 996102
rect 151261 996099 151327 996102
rect 149838 995830 150726 995890
rect 110781 995754 110847 995757
rect 106598 995752 110847 995754
rect 106598 995696 110786 995752
rect 110842 995696 110847 995752
rect 106598 995694 110847 995696
rect 110781 995691 110847 995694
rect 142797 995752 142906 995757
rect 142797 995696 142802 995752
rect 142858 995696 142906 995752
rect 142797 995694 142906 995696
rect 142797 995691 142863 995694
rect 110597 995618 110663 995621
rect 105862 995616 110663 995618
rect 105862 995560 110602 995616
rect 110658 995560 110663 995616
rect 105862 995558 110663 995560
rect 87781 995555 87847 995556
rect 81617 995480 82830 995482
rect 81617 995424 81622 995480
rect 81678 995424 82830 995480
rect 81617 995422 82830 995424
rect 85297 995482 85363 995485
rect 92614 995482 92674 995558
rect 100201 995555 100267 995558
rect 104157 995555 104223 995558
rect 104341 995555 104407 995558
rect 110597 995555 110663 995558
rect 137369 995618 137435 995621
rect 152322 995618 152382 996132
rect 152549 996104 152554 996160
rect 152610 996104 152720 996160
rect 152549 996102 152720 996104
rect 152917 996160 153180 996162
rect 152917 996104 152922 996160
rect 152978 996104 153180 996160
rect 152917 996102 153180 996104
rect 153377 996160 153548 996162
rect 153377 996104 153382 996160
rect 153438 996104 153548 996160
rect 153377 996102 153548 996104
rect 154573 996160 154836 996162
rect 154573 996104 154578 996160
rect 154634 996104 154836 996160
rect 156965 996160 157228 996162
rect 154573 996102 154836 996104
rect 152549 996099 152615 996102
rect 152917 996099 152983 996102
rect 153377 996099 153443 996102
rect 154573 996099 154639 996102
rect 137369 995616 152382 995618
rect 137369 995560 137374 995616
rect 137430 995560 152382 995616
rect 137369 995558 152382 995560
rect 137369 995555 137435 995558
rect 85297 995480 92674 995482
rect 85297 995424 85302 995480
rect 85358 995424 92674 995480
rect 85297 995422 92674 995424
rect 133689 995482 133755 995485
rect 141049 995482 141115 995485
rect 156002 995482 156062 996132
rect 156965 996104 156970 996160
rect 157026 996104 157228 996160
rect 156965 996102 157228 996104
rect 157793 996160 158056 996162
rect 157793 996104 157798 996160
rect 157854 996132 158056 996160
rect 159449 996160 159712 996162
rect 157854 996104 158086 996132
rect 157793 996102 158086 996104
rect 156965 996099 157031 996102
rect 157793 996099 157859 996102
rect 158026 995618 158086 996102
rect 159449 996104 159454 996160
rect 159510 996132 159712 996160
rect 208656 996160 208827 996162
rect 159510 996104 159742 996132
rect 159449 996102 159742 996104
rect 159449 996099 159515 996102
rect 159682 995754 159742 996102
rect 160050 995890 160110 996132
rect 168373 995890 168439 995893
rect 160050 995888 168439 995890
rect 160050 995832 168378 995888
rect 168434 995832 168439 995888
rect 160050 995830 168439 995832
rect 200806 995890 200866 996132
rect 201726 995890 201786 996132
rect 200806 995830 201786 995890
rect 206970 995893 207030 996132
rect 206970 995888 207079 995893
rect 206970 995832 207018 995888
rect 207074 995832 207079 995888
rect 206970 995830 207079 995832
rect 168373 995827 168439 995830
rect 207013 995827 207079 995830
rect 162945 995754 163011 995757
rect 159682 995752 163011 995754
rect 159682 995696 162950 995752
rect 163006 995696 163011 995752
rect 159682 995694 163011 995696
rect 162945 995691 163011 995694
rect 187601 995754 187667 995757
rect 187734 995754 187740 995756
rect 187601 995752 187740 995754
rect 187601 995696 187606 995752
rect 187662 995696 187740 995752
rect 187601 995694 187740 995696
rect 187601 995691 187667 995694
rect 187734 995692 187740 995694
rect 187804 995692 187810 995756
rect 162853 995618 162919 995621
rect 158026 995616 162919 995618
rect 158026 995560 162858 995616
rect 162914 995560 162919 995616
rect 158026 995558 162919 995560
rect 162853 995555 162919 995558
rect 192477 995618 192543 995621
rect 207430 995618 207490 996132
rect 207798 995621 207858 996132
rect 208656 996104 208766 996160
rect 208822 996104 208827 996160
rect 208656 996102 208827 996104
rect 209484 996160 209655 996162
rect 209484 996104 209594 996160
rect 209650 996104 209655 996160
rect 209484 996102 209655 996104
rect 211140 996160 211311 996162
rect 211140 996104 211250 996160
rect 211306 996104 211311 996160
rect 211613 996162 211679 996165
rect 253657 996162 253723 996165
rect 254117 996162 254183 996165
rect 254485 996162 254551 996165
rect 305269 996162 305335 996165
rect 305729 996162 305795 996165
rect 306465 996162 306531 996165
rect 306925 996162 306991 996165
rect 307293 996162 307359 996165
rect 307753 996162 307819 996165
rect 310145 996162 310211 996165
rect 362585 996162 362651 996165
rect 364241 996162 364307 996165
rect 364701 996162 364767 996165
rect 365069 996162 365135 996165
rect 371509 996162 371575 996165
rect 211613 996160 211876 996162
rect 211140 996102 211311 996104
rect 208761 996099 208827 996102
rect 209589 996099 209655 996102
rect 211245 996099 211311 996102
rect 211478 995890 211538 996132
rect 211613 996104 211618 996160
rect 211674 996104 211876 996160
rect 211613 996102 211876 996104
rect 253657 996160 253920 996162
rect 253657 996104 253662 996160
rect 253718 996104 253920 996160
rect 253657 996102 253920 996104
rect 254117 996160 254380 996162
rect 254117 996104 254122 996160
rect 254178 996104 254380 996160
rect 254117 996102 254380 996104
rect 254485 996160 254748 996162
rect 254485 996104 254490 996160
rect 254546 996104 254748 996160
rect 305269 996160 305532 996162
rect 254485 996102 254748 996104
rect 211613 996099 211679 996102
rect 253657 996099 253723 996102
rect 254117 996099 254183 996102
rect 254485 996099 254551 996102
rect 246941 996026 247007 996029
rect 237330 996024 247007 996026
rect 237330 995968 246946 996024
rect 247002 995968 247007 996024
rect 237330 995966 247007 995968
rect 216581 995890 216647 995893
rect 211478 995888 216647 995890
rect 211478 995832 216586 995888
rect 216642 995832 216647 995888
rect 211478 995830 216647 995832
rect 216581 995827 216647 995830
rect 234521 995754 234587 995757
rect 237330 995754 237390 995966
rect 246941 995963 247007 995966
rect 255086 995890 255146 996132
rect 240734 995830 255146 995890
rect 234521 995752 237390 995754
rect 234521 995696 234526 995752
rect 234582 995696 237390 995752
rect 234521 995694 237390 995696
rect 240041 995754 240107 995757
rect 240734 995754 240794 995830
rect 240041 995752 240794 995754
rect 240041 995696 240046 995752
rect 240102 995696 240794 995752
rect 240041 995694 240794 995696
rect 234521 995691 234587 995694
rect 240041 995691 240107 995694
rect 192477 995616 207490 995618
rect 192477 995560 192482 995616
rect 192538 995560 207490 995616
rect 192477 995558 207490 995560
rect 207749 995616 207858 995621
rect 207749 995560 207754 995616
rect 207810 995560 207858 995616
rect 207749 995558 207858 995560
rect 242065 995618 242131 995621
rect 255546 995618 255606 996132
rect 242065 995616 255606 995618
rect 242065 995560 242070 995616
rect 242126 995560 255606 995616
rect 242065 995558 255606 995560
rect 192477 995555 192543 995558
rect 207749 995555 207815 995558
rect 242065 995555 242131 995558
rect 133689 995480 140790 995482
rect 133689 995424 133694 995480
rect 133750 995424 140790 995480
rect 133689 995422 140790 995424
rect 81617 995419 81683 995422
rect 85297 995419 85363 995422
rect 133689 995419 133755 995422
rect 81985 995346 82051 995349
rect 96521 995346 96587 995349
rect 81985 995344 96587 995346
rect 81985 995288 81990 995344
rect 82046 995288 96526 995344
rect 96582 995288 96587 995344
rect 81985 995286 96587 995288
rect 140730 995346 140790 995422
rect 141049 995480 156062 995482
rect 141049 995424 141054 995480
rect 141110 995424 156062 995480
rect 141049 995422 156062 995424
rect 235901 995482 235967 995485
rect 255914 995482 255974 996132
rect 235901 995480 255974 995482
rect 235901 995424 235906 995480
rect 235962 995424 255974 995480
rect 235901 995422 255974 995424
rect 141049 995419 141115 995422
rect 235901 995419 235967 995422
rect 146201 995346 146267 995349
rect 140730 995344 146267 995346
rect 140730 995288 146206 995344
rect 146262 995288 146267 995344
rect 140730 995286 146267 995288
rect 81985 995283 82051 995286
rect 96521 995283 96587 995286
rect 146201 995283 146267 995286
rect 236223 995346 236289 995349
rect 254485 995346 254551 995349
rect 236223 995344 254551 995346
rect 236223 995288 236228 995344
rect 236284 995288 254490 995344
rect 254546 995288 254551 995344
rect 236223 995286 254551 995288
rect 236223 995283 236289 995286
rect 254485 995283 254551 995286
rect 80697 995210 80763 995213
rect 84469 995210 84535 995213
rect 99281 995210 99347 995213
rect 80697 995208 82830 995210
rect 80697 995152 80702 995208
rect 80758 995152 82830 995208
rect 80697 995150 82830 995152
rect 80697 995147 80763 995150
rect 82770 995074 82830 995150
rect 84469 995208 99347 995210
rect 84469 995152 84474 995208
rect 84530 995152 99286 995208
rect 99342 995152 99347 995208
rect 84469 995150 99347 995152
rect 84469 995147 84535 995150
rect 99281 995147 99347 995150
rect 234935 995210 235001 995213
rect 256374 995210 256434 996132
rect 234935 995208 256434 995210
rect 234935 995152 234940 995208
rect 234996 995152 256434 995208
rect 234935 995150 256434 995152
rect 234935 995147 235001 995150
rect 92749 995074 92815 995077
rect 82770 995072 92815 995074
rect 82770 995016 92754 995072
rect 92810 995016 92815 995072
rect 82770 995014 92815 995016
rect 92749 995011 92815 995014
rect 232221 994122 232287 994125
rect 253841 994122 253907 994125
rect 232221 994120 253907 994122
rect 232221 994064 232226 994120
rect 232282 994064 253846 994120
rect 253902 994064 253907 994120
rect 232221 994062 253907 994064
rect 232221 994059 232287 994062
rect 253841 994059 253907 994062
rect 232865 993986 232931 993989
rect 259134 993986 259194 996132
rect 300761 995890 300827 995893
rect 304214 995890 304274 996132
rect 305134 995890 305194 996132
rect 305269 996104 305274 996160
rect 305330 996104 305532 996160
rect 305269 996102 305532 996104
rect 305729 996160 305900 996162
rect 305729 996104 305734 996160
rect 305790 996104 305900 996160
rect 306465 996160 306728 996162
rect 305729 996102 305900 996104
rect 305269 996099 305335 996102
rect 305729 996099 305795 996102
rect 306330 995890 306390 996132
rect 306465 996104 306470 996160
rect 306526 996104 306728 996160
rect 306465 996102 306728 996104
rect 306925 996160 307188 996162
rect 306925 996104 306930 996160
rect 306986 996104 307188 996160
rect 306925 996102 307188 996104
rect 307293 996160 307556 996162
rect 307293 996104 307298 996160
rect 307354 996104 307556 996160
rect 307293 996102 307556 996104
rect 307753 996160 307924 996162
rect 307753 996104 307758 996160
rect 307814 996104 307924 996160
rect 310145 996160 310408 996162
rect 307753 996102 307924 996104
rect 306465 996099 306531 996102
rect 306925 996099 306991 996102
rect 307293 996099 307359 996102
rect 307753 996099 307819 996102
rect 292254 995830 300594 995890
rect 288065 995754 288131 995757
rect 292254 995754 292314 995830
rect 288065 995752 292314 995754
rect 288065 995696 288070 995752
rect 288126 995696 292314 995752
rect 288065 995694 292314 995696
rect 292481 995754 292547 995757
rect 300534 995754 300594 995830
rect 300761 995888 305194 995890
rect 300761 995832 300766 995888
rect 300822 995832 305194 995888
rect 300761 995830 305194 995832
rect 305318 995830 306390 995890
rect 300761 995827 300827 995830
rect 305318 995754 305378 995830
rect 292481 995752 300410 995754
rect 292481 995696 292486 995752
rect 292542 995696 300410 995752
rect 292481 995694 300410 995696
rect 300534 995694 305378 995754
rect 288065 995691 288131 995694
rect 292481 995691 292547 995694
rect 290641 995618 290707 995621
rect 300209 995618 300275 995621
rect 290641 995616 300275 995618
rect 290641 995560 290646 995616
rect 290702 995560 300214 995616
rect 300270 995560 300275 995616
rect 290641 995558 300275 995560
rect 300350 995618 300410 995694
rect 305269 995618 305335 995621
rect 300350 995616 305335 995618
rect 300350 995560 305274 995616
rect 305330 995560 305335 995616
rect 300350 995558 305335 995560
rect 290641 995555 290707 995558
rect 300209 995555 300275 995558
rect 305269 995555 305335 995558
rect 291101 995482 291167 995485
rect 297265 995482 297331 995485
rect 308722 995482 308782 996132
rect 310145 996104 310150 996160
rect 310206 996104 310408 996160
rect 362388 996160 362651 996162
rect 310145 996102 310408 996104
rect 310145 996099 310211 996102
rect 353661 995890 353727 995893
rect 354630 995890 354690 996132
rect 355458 995890 355518 996132
rect 353661 995888 355518 995890
rect 353661 995832 353666 995888
rect 353722 995832 355518 995888
rect 353661 995830 355518 995832
rect 353661 995827 353727 995830
rect 359138 995621 359198 996132
rect 359138 995616 359247 995621
rect 359138 995560 359186 995616
rect 359242 995560 359247 995616
rect 359138 995558 359247 995560
rect 361622 995618 361682 996132
rect 361990 995754 362050 996132
rect 362388 996104 362590 996160
rect 362646 996104 362651 996160
rect 364044 996160 364307 996162
rect 362388 996102 362651 996104
rect 362585 996099 362651 996102
rect 362818 995890 362878 996132
rect 364044 996104 364246 996160
rect 364302 996104 364307 996160
rect 364044 996102 364307 996104
rect 364504 996160 364767 996162
rect 364504 996104 364706 996160
rect 364762 996104 364767 996160
rect 364504 996102 364767 996104
rect 364872 996160 365135 996162
rect 364872 996104 365074 996160
rect 365130 996104 365135 996160
rect 364872 996102 365135 996104
rect 365700 996160 371575 996162
rect 365700 996104 371514 996160
rect 371570 996104 371575 996160
rect 365700 996102 371575 996104
rect 364241 996099 364307 996102
rect 364701 996099 364767 996102
rect 365069 996099 365135 996102
rect 371509 996099 371575 996102
rect 367093 995890 367159 995893
rect 362818 995888 367159 995890
rect 362818 995832 367098 995888
rect 367154 995832 367159 995888
rect 362818 995830 367159 995832
rect 367093 995827 367159 995830
rect 388118 995757 388178 996374
rect 461025 996432 476436 996434
rect 461025 996376 461030 996432
rect 461086 996376 476436 996432
rect 461025 996374 476436 996376
rect 461025 996371 461091 996374
rect 476430 996372 476436 996374
rect 476500 996372 476506 996436
rect 519537 996434 519603 996437
rect 526110 996434 526116 996436
rect 519537 996432 526116 996434
rect 519537 996376 519542 996432
rect 519598 996376 526116 996432
rect 519537 996374 526116 996376
rect 519537 996371 519603 996374
rect 526110 996372 526116 996374
rect 526180 996372 526186 996436
rect 421606 995890 421666 996132
rect 422526 995890 422586 996132
rect 421606 995830 422586 995890
rect 498702 995890 498762 996132
rect 499438 995890 499498 996132
rect 498702 995830 499498 995890
rect 367185 995754 367251 995757
rect 361990 995752 367251 995754
rect 361990 995696 367190 995752
rect 367246 995696 367251 995752
rect 361990 995694 367251 995696
rect 388118 995752 388227 995757
rect 388118 995696 388166 995752
rect 388222 995696 388227 995752
rect 388118 995694 388227 995696
rect 367185 995691 367251 995694
rect 388161 995691 388227 995694
rect 447133 995754 447199 995757
rect 481449 995754 481515 995757
rect 447133 995752 481515 995754
rect 447133 995696 447138 995752
rect 447194 995696 481454 995752
rect 481510 995696 481515 995752
rect 447133 995694 481515 995696
rect 447133 995691 447199 995694
rect 481449 995691 481515 995694
rect 503578 995621 503638 996132
rect 532190 995757 532250 996510
rect 558453 996162 558519 996165
rect 558256 996160 558519 996162
rect 549437 995890 549503 995893
rect 550406 995890 550466 996132
rect 551326 995890 551386 996132
rect 549437 995888 551386 995890
rect 549437 995832 549442 995888
rect 549498 995832 551386 995888
rect 549437 995830 551386 995832
rect 549437 995827 549503 995830
rect 523861 995754 523927 995757
rect 527909 995754 527975 995757
rect 523861 995752 527975 995754
rect 523861 995696 523866 995752
rect 523922 995696 527914 995752
rect 527970 995696 527975 995752
rect 523861 995694 527975 995696
rect 532190 995752 532299 995757
rect 532190 995696 532238 995752
rect 532294 995696 532299 995752
rect 532190 995694 532299 995696
rect 523861 995691 523927 995694
rect 527909 995691 527975 995694
rect 532233 995691 532299 995694
rect 555006 995621 555066 996132
rect 367461 995618 367527 995621
rect 361622 995616 367527 995618
rect 361622 995560 367466 995616
rect 367522 995560 367527 995616
rect 361622 995558 367527 995560
rect 359181 995555 359247 995558
rect 367461 995555 367527 995558
rect 471697 995618 471763 995621
rect 477677 995618 477743 995621
rect 471697 995616 477743 995618
rect 471697 995560 471702 995616
rect 471758 995560 477682 995616
rect 477738 995560 477743 995616
rect 471697 995558 477743 995560
rect 503578 995616 503687 995621
rect 503578 995560 503626 995616
rect 503682 995560 503687 995616
rect 503578 995558 503687 995560
rect 471697 995555 471763 995558
rect 477677 995555 477743 995558
rect 503621 995555 503687 995558
rect 521561 995618 521627 995621
rect 530117 995618 530183 995621
rect 521561 995616 530183 995618
rect 521561 995560 521566 995616
rect 521622 995560 530122 995616
rect 530178 995560 530183 995616
rect 521561 995558 530183 995560
rect 555006 995616 555115 995621
rect 555006 995560 555054 995616
rect 555110 995560 555115 995616
rect 555006 995558 555115 995560
rect 521561 995555 521627 995558
rect 530117 995555 530183 995558
rect 555049 995555 555115 995558
rect 476481 995484 476547 995485
rect 526161 995484 526227 995485
rect 291101 995480 295350 995482
rect 291101 995424 291106 995480
rect 291162 995424 295350 995480
rect 291101 995422 295350 995424
rect 291101 995419 291167 995422
rect 295290 995346 295350 995422
rect 297265 995480 308782 995482
rect 297265 995424 297270 995480
rect 297326 995424 308782 995480
rect 297265 995422 308782 995424
rect 297265 995419 297331 995422
rect 476430 995420 476436 995484
rect 476500 995482 476547 995484
rect 476500 995480 476592 995482
rect 476542 995424 476592 995480
rect 476500 995422 476592 995424
rect 476500 995420 476547 995422
rect 526110 995420 526116 995484
rect 526180 995482 526227 995484
rect 526180 995480 526272 995482
rect 526222 995424 526272 995480
rect 526180 995422 526272 995424
rect 526180 995420 526227 995422
rect 476481 995419 476547 995420
rect 526161 995419 526227 995420
rect 305729 995346 305795 995349
rect 295290 995344 305795 995346
rect 295290 995288 305734 995344
rect 305790 995288 305795 995344
rect 295290 995286 305795 995288
rect 305729 995283 305795 995286
rect 469397 995346 469463 995349
rect 481081 995346 481147 995349
rect 469397 995344 481147 995346
rect 469397 995288 469402 995344
rect 469458 995288 481086 995344
rect 481142 995288 481147 995344
rect 469397 995286 481147 995288
rect 469397 995283 469463 995286
rect 481081 995283 481147 995286
rect 521285 995346 521351 995349
rect 533981 995346 534047 995349
rect 537385 995346 537451 995349
rect 521285 995344 534047 995346
rect 521285 995288 521290 995344
rect 521346 995288 533986 995344
rect 534042 995288 534047 995344
rect 521285 995286 534047 995288
rect 521285 995283 521351 995286
rect 533981 995283 534047 995286
rect 535410 995344 537451 995346
rect 535410 995288 537390 995344
rect 537446 995288 537451 995344
rect 535410 995286 537451 995288
rect 555742 995346 555802 996132
rect 556570 995482 556630 996132
rect 557398 995618 557458 996132
rect 557766 995757 557826 996132
rect 558256 996104 558458 996160
rect 558514 996104 558519 996160
rect 559281 996162 559347 996165
rect 559281 996160 559452 996162
rect 558256 996102 558519 996104
rect 558453 996099 558519 996102
rect 558594 995757 558654 996132
rect 557717 995752 557826 995757
rect 557717 995696 557722 995752
rect 557778 995696 557826 995752
rect 557717 995694 557826 995696
rect 558545 995752 558654 995757
rect 558545 995696 558550 995752
rect 558606 995696 558654 995752
rect 558545 995694 558654 995696
rect 559054 995754 559114 996132
rect 559281 996104 559286 996160
rect 559342 996104 559452 996160
rect 559281 996102 559452 996104
rect 559281 996099 559347 996102
rect 559790 995890 559850 996132
rect 564709 995890 564775 995893
rect 559790 995888 564775 995890
rect 559790 995832 564714 995888
rect 564770 995832 564775 995888
rect 559790 995830 564775 995832
rect 564709 995827 564775 995830
rect 564341 995754 564407 995757
rect 559054 995752 564407 995754
rect 559054 995696 564346 995752
rect 564402 995696 564407 995752
rect 559054 995694 564407 995696
rect 557717 995691 557783 995694
rect 558545 995691 558611 995694
rect 564341 995691 564407 995694
rect 561673 995618 561739 995621
rect 557398 995616 561739 995618
rect 557398 995560 561678 995616
rect 561734 995560 561739 995616
rect 557398 995558 561739 995560
rect 561673 995555 561739 995558
rect 561489 995482 561555 995485
rect 556570 995480 561555 995482
rect 556570 995424 561494 995480
rect 561550 995424 561555 995480
rect 556570 995422 561555 995424
rect 561489 995419 561555 995422
rect 561305 995346 561371 995349
rect 555742 995344 561371 995346
rect 555742 995288 561310 995344
rect 561366 995288 561371 995344
rect 555742 995286 561371 995288
rect 521653 995210 521719 995213
rect 535410 995210 535470 995286
rect 537385 995283 537451 995286
rect 561305 995283 561371 995286
rect 521653 995208 535470 995210
rect 521653 995152 521658 995208
rect 521714 995152 535470 995208
rect 521653 995150 535470 995152
rect 638539 995210 638605 995213
rect 641161 995210 641227 995213
rect 638539 995208 641227 995210
rect 638539 995152 638544 995208
rect 638600 995152 641166 995208
rect 641222 995152 641227 995208
rect 638539 995150 641227 995152
rect 521653 995147 521719 995150
rect 638539 995147 638605 995150
rect 641161 995147 641227 995150
rect 568665 994258 568731 994261
rect 634813 994258 634879 994261
rect 568665 994256 634879 994258
rect 568665 994200 568670 994256
rect 568726 994200 634818 994256
rect 634874 994200 634879 994256
rect 568665 994198 634879 994200
rect 568665 994195 568731 994198
rect 634813 994195 634879 994198
rect 568573 994122 568639 994125
rect 637021 994122 637087 994125
rect 568573 994120 637087 994122
rect 568573 994064 568578 994120
rect 568634 994064 637026 994120
rect 637082 994064 637087 994120
rect 568573 994062 637087 994064
rect 568573 994059 568639 994062
rect 637021 994059 637087 994062
rect 232865 993984 259194 993986
rect 232865 993928 232870 993984
rect 232926 993928 259194 993984
rect 232865 993926 259194 993928
rect 570137 993986 570203 993989
rect 635181 993986 635247 993989
rect 570137 993984 635247 993986
rect 570137 993928 570142 993984
rect 570198 993928 635186 993984
rect 635242 993928 635247 993984
rect 570137 993926 635247 993928
rect 232865 993923 232931 993926
rect 570137 993923 570203 993926
rect 635181 993923 635247 993926
rect 80145 993850 80211 993853
rect 100201 993850 100267 993853
rect 80145 993848 100267 993850
rect 80145 993792 80150 993848
rect 80206 993792 100206 993848
rect 100262 993792 100267 993848
rect 80145 993790 100267 993792
rect 80145 993787 80211 993790
rect 100201 993787 100267 993790
rect 243261 993850 243327 993853
rect 316769 993850 316835 993853
rect 243261 993848 316835 993850
rect 243261 993792 243266 993848
rect 243322 993792 316774 993848
rect 316830 993792 316835 993848
rect 243261 993790 316835 993792
rect 243261 993787 243327 993790
rect 316769 993787 316835 993790
rect 378133 993850 378199 993853
rect 396993 993850 397059 993853
rect 378133 993848 397059 993850
rect 378133 993792 378138 993848
rect 378194 993792 396998 993848
rect 397054 993792 397059 993848
rect 378133 993790 397059 993792
rect 378133 993787 378199 993790
rect 396993 993787 397059 993790
rect 561305 993850 561371 993853
rect 629661 993850 629727 993853
rect 561305 993848 629727 993850
rect 561305 993792 561310 993848
rect 561366 993792 629666 993848
rect 629722 993792 629727 993848
rect 561305 993790 629727 993792
rect 561305 993787 561371 993790
rect 629661 993787 629727 993790
rect 78305 993714 78371 993717
rect 104341 993714 104407 993717
rect 78305 993712 104407 993714
rect 78305 993656 78310 993712
rect 78366 993656 104346 993712
rect 104402 993656 104407 993712
rect 78305 993654 104407 993656
rect 78305 993651 78371 993654
rect 104341 993651 104407 993654
rect 191833 993714 191899 993717
rect 248321 993714 248387 993717
rect 191833 993712 248387 993714
rect 191833 993656 191838 993712
rect 191894 993656 248326 993712
rect 248382 993656 248387 993712
rect 191833 993654 248387 993656
rect 191833 993651 191899 993654
rect 248321 993651 248387 993654
rect 294505 993714 294571 993717
rect 366173 993714 366239 993717
rect 294505 993712 366239 993714
rect 294505 993656 294510 993712
rect 294566 993656 366178 993712
rect 366234 993656 366239 993712
rect 294505 993654 366239 993656
rect 294505 993651 294571 993654
rect 366173 993651 366239 993654
rect 374453 993714 374519 993717
rect 395153 993714 395219 993717
rect 374453 993712 395219 993714
rect 374453 993656 374458 993712
rect 374514 993656 395158 993712
rect 395214 993656 395219 993712
rect 374453 993654 395219 993656
rect 374453 993651 374519 993654
rect 395153 993651 395219 993654
rect 447317 993714 447383 993717
rect 478597 993714 478663 993717
rect 447317 993712 478663 993714
rect 447317 993656 447322 993712
rect 447378 993656 478602 993712
rect 478658 993656 478663 993712
rect 447317 993654 478663 993656
rect 447317 993651 447383 993654
rect 478597 993651 478663 993654
rect 561489 993714 561555 993717
rect 638861 993714 638927 993717
rect 561489 993712 638927 993714
rect 561489 993656 561494 993712
rect 561550 993656 638866 993712
rect 638922 993656 638927 993712
rect 561489 993654 638927 993656
rect 561489 993651 561555 993654
rect 638861 993651 638927 993654
rect 564433 985826 564499 985829
rect 674782 985826 674788 985828
rect 564433 985824 674788 985826
rect 564433 985768 564438 985824
rect 564494 985768 674788 985824
rect 564433 985766 674788 985768
rect 564433 985763 564499 985766
rect 674782 985764 674788 985766
rect 674852 985764 674858 985828
rect 561673 985690 561739 985693
rect 674966 985690 674972 985692
rect 561673 985688 674972 985690
rect 561673 985632 561678 985688
rect 561734 985632 674972 985688
rect 561673 985630 674972 985632
rect 561673 985627 561739 985630
rect 674966 985628 674972 985630
rect 675036 985628 675042 985692
rect 44030 985492 44036 985556
rect 44100 985554 44106 985556
rect 672717 985554 672783 985557
rect 44100 985552 672783 985554
rect 44100 985496 672722 985552
rect 672778 985496 672783 985552
rect 44100 985494 672783 985496
rect 44100 985492 44106 985494
rect 672717 985491 672783 985494
rect 43478 985356 43484 985420
rect 43548 985418 43554 985420
rect 672533 985418 672599 985421
rect 43548 985416 672599 985418
rect 43548 985360 672538 985416
rect 672594 985360 672599 985416
rect 43548 985358 672599 985360
rect 43548 985356 43554 985358
rect 672533 985355 672599 985358
rect 43662 983316 43668 983380
rect 43732 983378 43738 983380
rect 669129 983378 669195 983381
rect 43732 983376 669195 983378
rect 43732 983320 669134 983376
rect 669190 983320 669195 983376
rect 43732 983318 669195 983320
rect 43732 983316 43738 983318
rect 669129 983315 669195 983318
rect 43294 983180 43300 983244
rect 43364 983242 43370 983244
rect 669681 983242 669747 983245
rect 43364 983240 669747 983242
rect 43364 983184 669686 983240
rect 669742 983184 669747 983240
rect 43364 983182 669747 983184
rect 43364 983180 43370 983182
rect 669681 983179 669747 983182
rect 43846 983044 43852 983108
rect 43916 983106 43922 983108
rect 670233 983106 670299 983109
rect 43916 983104 670299 983106
rect 43916 983048 670238 983104
rect 670294 983048 670299 983104
rect 43916 983046 670299 983048
rect 43916 983044 43922 983046
rect 670233 983043 670299 983046
rect 43110 982908 43116 982972
rect 43180 982970 43186 982972
rect 670049 982970 670115 982973
rect 43180 982968 670115 982970
rect 43180 982912 670054 982968
rect 670110 982912 670115 982968
rect 43180 982910 670115 982912
rect 43180 982908 43186 982910
rect 670049 982907 670115 982910
rect 58433 976034 58499 976037
rect 58433 976032 64492 976034
rect 58433 975976 58438 976032
rect 58494 975976 64492 976032
rect 58433 975974 64492 975976
rect 58433 975971 58499 975974
rect 655513 975898 655579 975901
rect 650164 975896 655579 975898
rect 650164 975840 655518 975896
rect 655574 975840 655579 975896
rect 650164 975838 655579 975840
rect 655513 975835 655579 975838
rect 41454 968764 41460 968828
rect 41524 968826 41530 968828
rect 41781 968826 41847 968829
rect 41524 968824 41847 968826
rect 41524 968768 41786 968824
rect 41842 968768 41847 968824
rect 41524 968766 41847 968768
rect 41524 968764 41530 968766
rect 41781 968763 41847 968766
rect 41638 965092 41644 965156
rect 41708 965154 41714 965156
rect 41781 965154 41847 965157
rect 41708 965152 41847 965154
rect 41708 965096 41786 965152
rect 41842 965096 41847 965152
rect 41708 965094 41847 965096
rect 41708 965092 41714 965094
rect 41781 965091 41847 965094
rect 41781 963388 41847 963389
rect 41781 963384 41828 963388
rect 41892 963386 41898 963388
rect 41781 963328 41786 963384
rect 41781 963324 41828 963328
rect 41892 963326 41938 963386
rect 41892 963324 41898 963326
rect 41781 963323 41847 963324
rect 57973 962978 58039 962981
rect 57973 962976 64492 962978
rect 57973 962920 57978 962976
rect 58034 962920 64492 962976
rect 57973 962918 64492 962920
rect 57973 962915 58039 962918
rect 655697 962570 655763 962573
rect 650164 962568 655763 962570
rect 650164 962512 655702 962568
rect 655758 962512 655763 962568
rect 650164 962510 655763 962512
rect 655697 962507 655763 962510
rect 58433 949922 58499 949925
rect 58433 949920 64492 949922
rect 58433 949864 58438 949920
rect 58494 949864 64492 949920
rect 58433 949862 64492 949864
rect 58433 949859 58499 949862
rect 35801 949514 35867 949517
rect 41822 949514 41828 949516
rect 35801 949512 41828 949514
rect 35801 949456 35806 949512
rect 35862 949456 41828 949512
rect 35801 949454 41828 949456
rect 35801 949451 35867 949454
rect 41822 949452 41828 949454
rect 41892 949452 41898 949516
rect 655789 949378 655855 949381
rect 650164 949376 655855 949378
rect 650164 949320 655794 949376
rect 655850 949320 655855 949376
rect 650164 949318 655855 949320
rect 655789 949315 655855 949318
rect 41505 943938 41571 943941
rect 41462 943936 41571 943938
rect 41462 943880 41510 943936
rect 41566 943880 41571 943936
rect 41462 943875 41571 943880
rect 41462 943500 41522 943875
rect 41781 943122 41847 943125
rect 41492 943120 41847 943122
rect 41492 943064 41786 943120
rect 41842 943064 41847 943120
rect 41492 943062 41847 943064
rect 41781 943059 41847 943062
rect 41781 942714 41847 942717
rect 41492 942712 41847 942714
rect 41492 942656 41786 942712
rect 41842 942656 41847 942712
rect 41492 942654 41847 942656
rect 41781 942651 41847 942654
rect 41873 942306 41939 942309
rect 41492 942304 41939 942306
rect 41492 942248 41878 942304
rect 41934 942248 41939 942304
rect 41492 942246 41939 942248
rect 41873 942243 41939 942246
rect 41965 941898 42031 941901
rect 41492 941896 42031 941898
rect 41492 941840 41970 941896
rect 42026 941840 42031 941896
rect 41492 941838 42031 941840
rect 41965 941835 42031 941838
rect 41781 941490 41847 941493
rect 41492 941488 41847 941490
rect 41492 941432 41786 941488
rect 41842 941432 41847 941488
rect 41492 941430 41847 941432
rect 41781 941427 41847 941430
rect 41873 941082 41939 941085
rect 41492 941080 41939 941082
rect 41492 941024 41878 941080
rect 41934 941024 41939 941080
rect 41492 941022 41939 941024
rect 41873 941019 41939 941022
rect 41492 940614 41752 940674
rect 41692 940541 41752 940614
rect 41689 940536 41755 940541
rect 41689 940480 41694 940536
rect 41750 940480 41755 940536
rect 41689 940475 41755 940480
rect 41965 940266 42031 940269
rect 41492 940264 42031 940266
rect 41492 940208 41970 940264
rect 42026 940208 42031 940264
rect 41492 940206 42031 940208
rect 41965 940203 42031 940206
rect 42977 939858 43043 939861
rect 41492 939856 43043 939858
rect 41492 939800 42982 939856
rect 43038 939800 43043 939856
rect 41492 939798 43043 939800
rect 42977 939795 43043 939798
rect 676262 939725 676322 939964
rect 676262 939720 676371 939725
rect 676262 939664 676310 939720
rect 676366 939664 676371 939720
rect 676262 939662 676371 939664
rect 676305 939659 676371 939662
rect 62297 939450 62363 939453
rect 41492 939448 62363 939450
rect 41492 939392 62302 939448
rect 62358 939392 62363 939448
rect 41492 939390 62363 939392
rect 62297 939387 62363 939390
rect 676121 939314 676187 939317
rect 676262 939314 676322 939556
rect 676121 939312 676322 939314
rect 676121 939256 676126 939312
rect 676182 939256 676322 939312
rect 676121 939254 676322 939256
rect 676121 939251 676187 939254
rect 42333 939042 42399 939045
rect 41492 939040 42399 939042
rect 41492 938984 42338 939040
rect 42394 938984 42399 939040
rect 41492 938982 42399 938984
rect 42333 938979 42399 938982
rect 676262 938909 676322 939148
rect 676213 938904 676322 938909
rect 676213 938848 676218 938904
rect 676274 938848 676322 938904
rect 676213 938846 676322 938848
rect 676213 938843 676279 938846
rect 675661 938770 675727 938773
rect 675661 938768 676292 938770
rect 675661 938712 675666 938768
rect 675722 938712 676292 938768
rect 675661 938710 676292 938712
rect 675661 938707 675727 938710
rect 42793 938634 42859 938637
rect 41492 938632 42859 938634
rect 41492 938576 42798 938632
rect 42854 938576 42859 938632
rect 41492 938574 42859 938576
rect 42793 938571 42859 938574
rect 41965 938498 42031 938501
rect 62481 938498 62547 938501
rect 41965 938496 62547 938498
rect 41965 938440 41970 938496
rect 42026 938440 62486 938496
rect 62542 938440 62547 938496
rect 41965 938438 62547 938440
rect 41965 938435 42031 938438
rect 62481 938435 62547 938438
rect 673862 938300 673868 938364
rect 673932 938362 673938 938364
rect 673932 938302 676292 938362
rect 673932 938300 673938 938302
rect 42241 938226 42307 938229
rect 41492 938224 42307 938226
rect 41492 938168 42246 938224
rect 42302 938168 42307 938224
rect 41492 938166 42307 938168
rect 42241 938163 42307 938166
rect 43253 937818 43319 937821
rect 41492 937816 43319 937818
rect 41492 937760 43258 937816
rect 43314 937760 43319 937816
rect 41492 937758 43319 937760
rect 43253 937755 43319 937758
rect 679022 937685 679082 937924
rect 678973 937680 679082 937685
rect 678973 937624 678978 937680
rect 679034 937624 679082 937680
rect 678973 937622 679082 937624
rect 678973 937619 679039 937622
rect 43069 937410 43135 937413
rect 41492 937408 43135 937410
rect 41492 937352 43074 937408
rect 43130 937352 43135 937408
rect 41492 937350 43135 937352
rect 43069 937347 43135 937350
rect 676814 937276 676874 937516
rect 676806 937212 676812 937276
rect 676876 937212 676882 937276
rect 674782 937076 674788 937140
rect 674852 937138 674858 937140
rect 674852 937078 676292 937138
rect 674852 937076 674858 937078
rect 41822 937002 41828 937004
rect 41492 936942 41828 937002
rect 41822 936940 41828 936942
rect 41892 936940 41898 937004
rect 58433 937002 58499 937005
rect 58433 937000 64492 937002
rect 58433 936944 58438 937000
rect 58494 936944 64492 937000
rect 58433 936942 64492 936944
rect 58433 936939 58499 936942
rect 41781 936594 41847 936597
rect 41492 936592 41847 936594
rect 41492 936536 41786 936592
rect 41842 936536 41847 936592
rect 41492 936534 41847 936536
rect 41781 936531 41847 936534
rect 676262 936461 676322 936700
rect 676213 936456 676322 936461
rect 676213 936400 676218 936456
rect 676274 936400 676322 936456
rect 676213 936398 676322 936400
rect 676213 936395 676279 936398
rect 674966 936260 674972 936324
rect 675036 936322 675042 936324
rect 675036 936262 676292 936322
rect 675036 936260 675042 936262
rect 43161 936186 43227 936189
rect 655605 936186 655671 936189
rect 41492 936184 43227 936186
rect 41492 936128 43166 936184
rect 43222 936128 43227 936184
rect 41492 936126 43227 936128
rect 650164 936184 655671 936186
rect 650164 936128 655610 936184
rect 655666 936128 655671 936184
rect 650164 936126 655671 936128
rect 43161 936123 43227 936126
rect 655605 936123 655671 936126
rect 676029 935914 676095 935917
rect 676029 935912 676292 935914
rect 676029 935856 676034 935912
rect 676090 935856 676292 935912
rect 676029 935854 676292 935856
rect 676029 935851 676095 935854
rect 43345 935778 43411 935781
rect 41492 935776 43411 935778
rect 41492 935720 43350 935776
rect 43406 935720 43411 935776
rect 41492 935718 43411 935720
rect 43345 935715 43411 935718
rect 675937 935506 676003 935509
rect 675937 935504 676292 935506
rect 675937 935448 675942 935504
rect 675998 935448 676292 935504
rect 675937 935446 676292 935448
rect 675937 935443 676003 935446
rect 42006 935370 42012 935372
rect 41492 935310 42012 935370
rect 42006 935308 42012 935310
rect 42076 935308 42082 935372
rect 676029 935098 676095 935101
rect 676029 935096 676292 935098
rect 676029 935040 676034 935096
rect 676090 935040 676292 935096
rect 676029 935038 676292 935040
rect 676029 935035 676095 935038
rect 35801 934962 35867 934965
rect 35788 934960 35867 934962
rect 35788 934904 35806 934960
rect 35862 934904 35867 934960
rect 35788 934902 35867 934904
rect 35801 934899 35867 934902
rect 675753 934690 675819 934693
rect 675753 934688 676292 934690
rect 675753 934632 675758 934688
rect 675814 934632 676292 934688
rect 675753 934630 676292 934632
rect 675753 934627 675819 934630
rect 35709 934554 35775 934557
rect 35709 934552 35788 934554
rect 35709 934496 35714 934552
rect 35770 934496 35788 934552
rect 35709 934494 35788 934496
rect 35709 934491 35775 934494
rect 675937 934282 676003 934285
rect 675937 934280 676292 934282
rect 675937 934224 675942 934280
rect 675998 934224 676292 934280
rect 675937 934222 676292 934224
rect 675937 934219 676003 934222
rect 35617 934146 35683 934149
rect 35604 934144 35683 934146
rect 35604 934088 35622 934144
rect 35678 934088 35683 934144
rect 35604 934086 35683 934088
rect 35617 934083 35683 934086
rect 676121 934010 676187 934013
rect 676121 934008 676322 934010
rect 676121 933952 676126 934008
rect 676182 933952 676322 934008
rect 676121 933950 676322 933952
rect 676121 933947 676187 933950
rect 676262 933844 676322 933950
rect 42885 933738 42951 933741
rect 41492 933736 42951 933738
rect 41492 933680 42890 933736
rect 42946 933680 42951 933736
rect 41492 933678 42951 933680
rect 42885 933675 42951 933678
rect 676029 933466 676095 933469
rect 676029 933464 676292 933466
rect 676029 933408 676034 933464
rect 676090 933408 676292 933464
rect 676029 933406 676292 933408
rect 676029 933403 676095 933406
rect 41781 933330 41847 933333
rect 41492 933328 41847 933330
rect 41492 933272 41786 933328
rect 41842 933272 41847 933328
rect 41492 933270 41847 933272
rect 41781 933267 41847 933270
rect 676029 933058 676095 933061
rect 676029 933056 676292 933058
rect 676029 933000 676034 933056
rect 676090 933000 676292 933056
rect 676029 932998 676292 933000
rect 676029 932995 676095 932998
rect 21958 932850 23490 932910
rect 23430 932076 23490 932850
rect 676121 932786 676187 932789
rect 676121 932784 676322 932786
rect 676121 932728 676126 932784
rect 676182 932728 676322 932784
rect 676121 932726 676322 932728
rect 676121 932723 676187 932726
rect 676262 932620 676322 932726
rect 41781 932514 41847 932517
rect 41492 932512 41847 932514
rect 41492 932456 41786 932512
rect 41842 932456 41847 932512
rect 41492 932454 41847 932456
rect 41781 932451 41847 932454
rect 675937 932242 676003 932245
rect 675937 932240 676292 932242
rect 675937 932184 675942 932240
rect 675998 932184 676292 932240
rect 675937 932182 676292 932184
rect 675937 932179 676003 932182
rect 676029 931834 676095 931837
rect 676029 931832 676292 931834
rect 676029 931776 676034 931832
rect 676090 931776 676292 931832
rect 676029 931774 676292 931776
rect 676029 931771 676095 931774
rect 676029 931426 676095 931429
rect 676029 931424 676292 931426
rect 676029 931368 676034 931424
rect 676090 931368 676292 931424
rect 676029 931366 676292 931368
rect 676029 931363 676095 931366
rect 675937 931018 676003 931021
rect 675937 931016 676292 931018
rect 675937 930960 675942 931016
rect 675998 930960 676292 931016
rect 675937 930958 676292 930960
rect 675937 930955 676003 930958
rect 676121 930746 676187 930749
rect 676121 930744 676322 930746
rect 676121 930688 676126 930744
rect 676182 930688 676322 930744
rect 676121 930686 676322 930688
rect 676121 930683 676187 930686
rect 676262 930580 676322 930686
rect 676029 930202 676095 930205
rect 676029 930200 676292 930202
rect 676029 930144 676034 930200
rect 676090 930144 676292 930200
rect 676029 930142 676292 930144
rect 676029 930139 676095 930142
rect 679022 929525 679082 929764
rect 678973 929520 679082 929525
rect 678973 929464 678978 929520
rect 679034 929464 679082 929520
rect 678973 929462 679082 929464
rect 678973 929459 679039 929462
rect 684542 929117 684602 929356
rect 678973 929114 679039 929117
rect 678973 929112 679082 929114
rect 678973 929056 678978 929112
rect 679034 929056 679082 929112
rect 678973 929051 679082 929056
rect 684493 929112 684602 929117
rect 684493 929056 684498 929112
rect 684554 929056 684602 929112
rect 684493 929054 684602 929056
rect 684493 929051 684559 929054
rect 679022 928948 679082 929051
rect 684493 928706 684559 928709
rect 684493 928704 684602 928706
rect 684493 928648 684498 928704
rect 684554 928648 684602 928704
rect 684493 928643 684602 928648
rect 684542 928540 684602 928643
rect 43110 927148 43116 927212
rect 43180 927210 43186 927212
rect 43989 927210 44055 927213
rect 43180 927208 44055 927210
rect 43180 927152 43994 927208
rect 44050 927152 44055 927208
rect 43180 927150 44055 927152
rect 43180 927148 43186 927150
rect 43989 927147 44055 927150
rect 58433 923810 58499 923813
rect 58433 923808 64492 923810
rect 58433 923752 58438 923808
rect 58494 923752 64492 923808
rect 58433 923750 64492 923752
rect 58433 923747 58499 923750
rect 654685 922722 654751 922725
rect 650164 922720 654751 922722
rect 650164 922664 654690 922720
rect 654746 922664 654751 922720
rect 650164 922662 654751 922664
rect 654685 922659 654751 922662
rect 41505 922042 41571 922045
rect 42558 922042 42564 922044
rect 41505 922040 42564 922042
rect 41505 921984 41510 922040
rect 41566 921984 42564 922040
rect 41505 921982 42564 921984
rect 41505 921979 41571 921982
rect 42558 921980 42564 921982
rect 42628 921980 42634 922044
rect 42793 922042 42859 922045
rect 43478 922042 43484 922044
rect 42793 922040 43484 922042
rect 42793 921984 42798 922040
rect 42854 921984 43484 922040
rect 42793 921982 43484 921984
rect 42793 921979 42859 921982
rect 43478 921980 43484 921982
rect 43548 921980 43554 922044
rect 58065 910754 58131 910757
rect 58065 910752 64492 910754
rect 58065 910696 58070 910752
rect 58126 910696 64492 910752
rect 58065 910694 64492 910696
rect 58065 910691 58131 910694
rect 654869 909530 654935 909533
rect 650164 909528 654935 909530
rect 650164 909472 654874 909528
rect 654930 909472 654935 909528
rect 650164 909470 654935 909472
rect 654869 909467 654935 909470
rect 58525 897834 58591 897837
rect 58525 897832 64492 897834
rect 58525 897776 58530 897832
rect 58586 897776 64492 897832
rect 58525 897774 64492 897776
rect 58525 897771 58591 897774
rect 654685 896202 654751 896205
rect 650164 896200 654751 896202
rect 650164 896144 654690 896200
rect 654746 896144 654751 896200
rect 650164 896142 654751 896144
rect 654685 896139 654751 896142
rect 58433 884778 58499 884781
rect 58433 884776 64492 884778
rect 58433 884720 58438 884776
rect 58494 884720 64492 884776
rect 58433 884718 64492 884720
rect 58433 884715 58499 884718
rect 655145 882874 655211 882877
rect 650164 882872 655211 882874
rect 650164 882816 655150 882872
rect 655206 882816 655211 882872
rect 650164 882814 655211 882816
rect 655145 882811 655211 882814
rect 675753 877298 675819 877301
rect 676070 877298 676076 877300
rect 675753 877296 676076 877298
rect 675753 877240 675758 877296
rect 675814 877240 676076 877296
rect 675753 877238 676076 877240
rect 675753 877235 675819 877238
rect 676070 877236 676076 877238
rect 676140 877236 676146 877300
rect 675661 876620 675727 876621
rect 675661 876616 675708 876620
rect 675772 876618 675778 876620
rect 675661 876560 675666 876616
rect 675661 876556 675708 876560
rect 675772 876558 675818 876618
rect 675772 876556 675778 876558
rect 675661 876555 675727 876556
rect 675385 875940 675451 875941
rect 675334 875938 675340 875940
rect 675294 875878 675340 875938
rect 675404 875936 675451 875940
rect 675446 875880 675451 875936
rect 675334 875876 675340 875878
rect 675404 875876 675451 875880
rect 675385 875875 675451 875876
rect 675477 874036 675543 874037
rect 675477 874032 675524 874036
rect 675588 874034 675594 874036
rect 675477 873976 675482 874032
rect 675477 873972 675524 873976
rect 675588 873974 675634 874034
rect 675588 873972 675594 873974
rect 675477 873971 675543 873972
rect 675753 872266 675819 872269
rect 675886 872266 675892 872268
rect 675753 872264 675892 872266
rect 675753 872208 675758 872264
rect 675814 872208 675892 872264
rect 675753 872206 675892 872208
rect 675753 872203 675819 872206
rect 675886 872204 675892 872206
rect 675956 872204 675962 872268
rect 58433 871722 58499 871725
rect 58433 871720 64492 871722
rect 58433 871664 58438 871720
rect 58494 871664 64492 871720
rect 58433 871662 64492 871664
rect 58433 871659 58499 871662
rect 656801 869682 656867 869685
rect 650164 869680 656867 869682
rect 650164 869624 656806 869680
rect 656862 869624 656867 869680
rect 650164 869622 656867 869624
rect 656801 869619 656867 869622
rect 58433 858666 58499 858669
rect 58433 858664 64492 858666
rect 58433 858608 58438 858664
rect 58494 858608 64492 858664
rect 58433 858606 64492 858608
rect 58433 858603 58499 858606
rect 655237 856354 655303 856357
rect 650164 856352 655303 856354
rect 650164 856296 655242 856352
rect 655298 856296 655303 856352
rect 650164 856294 655303 856296
rect 655237 856291 655303 856294
rect 58433 845610 58499 845613
rect 58433 845608 64492 845610
rect 58433 845552 58438 845608
rect 58494 845552 64492 845608
rect 58433 845550 64492 845552
rect 58433 845547 58499 845550
rect 654869 843026 654935 843029
rect 650164 843024 654935 843026
rect 650164 842968 654874 843024
rect 654930 842968 654935 843024
rect 650164 842966 654935 842968
rect 654869 842963 654935 842966
rect 57973 832554 58039 832557
rect 57973 832552 64492 832554
rect 57973 832496 57978 832552
rect 58034 832496 64492 832552
rect 57973 832494 64492 832496
rect 57973 832491 58039 832494
rect 655513 829834 655579 829837
rect 650164 829832 655579 829834
rect 650164 829776 655518 829832
rect 655574 829776 655579 829832
rect 650164 829774 655579 829776
rect 655513 829771 655579 829774
rect 59169 819498 59235 819501
rect 59169 819496 64492 819498
rect 59169 819440 59174 819496
rect 59230 819440 64492 819496
rect 59169 819438 64492 819440
rect 59169 819435 59235 819438
rect 41781 817730 41847 817733
rect 41492 817728 41847 817730
rect 41492 817672 41786 817728
rect 41842 817672 41847 817728
rect 41492 817670 41847 817672
rect 41781 817667 41847 817670
rect 41781 817322 41847 817325
rect 41492 817320 41847 817322
rect 41492 817264 41786 817320
rect 41842 817264 41847 817320
rect 41492 817262 41847 817264
rect 41781 817259 41847 817262
rect 53833 816914 53899 816917
rect 41492 816912 53899 816914
rect 41492 816856 53838 816912
rect 53894 816856 53899 816912
rect 41492 816854 53899 816856
rect 53833 816851 53899 816854
rect 41965 816506 42031 816509
rect 655053 816506 655119 816509
rect 41492 816504 42031 816506
rect 41492 816448 41970 816504
rect 42026 816448 42031 816504
rect 41492 816446 42031 816448
rect 650164 816504 655119 816506
rect 650164 816448 655058 816504
rect 655114 816448 655119 816504
rect 650164 816446 655119 816448
rect 41965 816443 42031 816446
rect 655053 816443 655119 816446
rect 42701 816098 42767 816101
rect 41492 816096 42767 816098
rect 41492 816040 42706 816096
rect 42762 816040 42767 816096
rect 41492 816038 42767 816040
rect 42701 816035 42767 816038
rect 41689 815824 41755 815829
rect 41689 815768 41694 815824
rect 41750 815768 41755 815824
rect 41689 815763 41755 815768
rect 41692 815690 41752 815763
rect 41492 815630 41752 815690
rect 43529 815282 43595 815285
rect 41492 815280 43595 815282
rect 41492 815224 43534 815280
rect 43590 815224 43595 815280
rect 41492 815222 43595 815224
rect 43529 815219 43595 815222
rect 43437 814874 43503 814877
rect 41492 814872 43503 814874
rect 41492 814816 43442 814872
rect 43498 814816 43503 814872
rect 41492 814814 43503 814816
rect 43437 814811 43503 814814
rect 41094 814299 41154 814436
rect 41094 814294 41203 814299
rect 41094 814238 41142 814294
rect 41198 814238 41203 814294
rect 41094 814236 41203 814238
rect 41137 814233 41203 814236
rect 41822 814132 41828 814196
rect 41892 814194 41898 814196
rect 41965 814194 42031 814197
rect 62849 814194 62915 814197
rect 41892 814192 62915 814194
rect 41892 814136 41970 814192
rect 42026 814136 62854 814192
rect 62910 814136 62915 814192
rect 41892 814134 62915 814136
rect 41892 814132 41898 814134
rect 41965 814131 42031 814134
rect 62849 814131 62915 814134
rect 41873 814058 41939 814061
rect 42333 814058 42399 814061
rect 41492 814056 42399 814058
rect 41492 814000 41878 814056
rect 41934 814000 42338 814056
rect 42394 814000 42399 814056
rect 41492 813998 42399 814000
rect 41873 813995 41939 813998
rect 42333 813995 42399 813998
rect 41781 813650 41847 813653
rect 41492 813648 41847 813650
rect 41492 813592 41786 813648
rect 41842 813592 41847 813648
rect 41492 813590 41847 813592
rect 41781 813587 41847 813590
rect 43345 813242 43411 813245
rect 41492 813240 43411 813242
rect 41492 813184 43350 813240
rect 43406 813184 43411 813240
rect 41492 813182 43411 813184
rect 43345 813179 43411 813182
rect 42885 812834 42951 812837
rect 41492 812832 42951 812834
rect 41492 812776 42890 812832
rect 42946 812776 42951 812832
rect 41492 812774 42951 812776
rect 42885 812771 42951 812774
rect 42977 812426 43043 812429
rect 41492 812424 43043 812426
rect 41492 812368 42982 812424
rect 43038 812368 43043 812424
rect 41492 812366 43043 812368
rect 42977 812363 43043 812366
rect 43069 812018 43135 812021
rect 41492 812016 43135 812018
rect 41492 811960 43074 812016
rect 43130 811960 43135 812016
rect 41492 811958 43135 811960
rect 43069 811955 43135 811958
rect 41781 811610 41847 811613
rect 41492 811608 41847 811610
rect 41492 811552 41786 811608
rect 41842 811552 41847 811608
rect 41492 811550 41847 811552
rect 41781 811547 41847 811550
rect 41965 811202 42031 811205
rect 41492 811200 42031 811202
rect 41492 811144 41970 811200
rect 42026 811144 42031 811200
rect 41492 811142 42031 811144
rect 41965 811139 42031 811142
rect 43805 810794 43871 810797
rect 41492 810792 43871 810794
rect 41492 810736 43810 810792
rect 43866 810736 43871 810792
rect 41492 810734 43871 810736
rect 43805 810731 43871 810734
rect 44081 810386 44147 810389
rect 41492 810384 44147 810386
rect 41492 810328 44086 810384
rect 44142 810328 44147 810384
rect 41492 810326 44147 810328
rect 44081 810323 44147 810326
rect 43897 809978 43963 809981
rect 41492 809976 43963 809978
rect 41492 809920 43902 809976
rect 43958 809920 43963 809976
rect 41492 809918 43963 809920
rect 43897 809915 43963 809918
rect 42609 809570 42675 809573
rect 41492 809568 42675 809570
rect 41492 809512 42614 809568
rect 42670 809512 42675 809568
rect 41492 809510 42675 809512
rect 42609 809507 42675 809510
rect 43253 809162 43319 809165
rect 41492 809160 43319 809162
rect 41492 809104 43258 809160
rect 43314 809104 43319 809160
rect 41492 809102 43319 809104
rect 43253 809099 43319 809102
rect 43621 808754 43687 808757
rect 41492 808752 43687 808754
rect 41492 808696 43626 808752
rect 43682 808696 43687 808752
rect 41492 808694 43687 808696
rect 43621 808691 43687 808694
rect 41781 808346 41847 808349
rect 41492 808344 41847 808346
rect 41492 808288 41786 808344
rect 41842 808288 41847 808344
rect 41492 808286 41847 808288
rect 41781 808283 41847 808286
rect 41873 807938 41939 807941
rect 41492 807936 41939 807938
rect 41492 807880 41878 807936
rect 41934 807880 41939 807936
rect 41492 807878 41939 807880
rect 41873 807875 41939 807878
rect 41781 807530 41847 807533
rect 41492 807528 41847 807530
rect 41492 807472 41786 807528
rect 41842 807472 41847 807528
rect 41492 807470 41847 807472
rect 41781 807467 41847 807470
rect 22694 806276 22754 807092
rect 41781 806714 41847 806717
rect 41492 806712 41847 806714
rect 41492 806656 41786 806712
rect 41842 806656 41847 806712
rect 41492 806654 41847 806656
rect 41781 806651 41847 806654
rect 58433 806578 58499 806581
rect 58433 806576 64492 806578
rect 58433 806520 58438 806576
rect 58494 806520 64492 806576
rect 58433 806518 64492 806520
rect 58433 806515 58499 806518
rect 656157 803314 656223 803317
rect 650164 803312 656223 803314
rect 650164 803256 656162 803312
rect 656218 803256 656223 803312
rect 650164 803254 656223 803256
rect 656157 803251 656223 803254
rect 674281 797738 674347 797741
rect 676254 797738 676260 797740
rect 674281 797736 676260 797738
rect 674281 797680 674286 797736
rect 674342 797680 676260 797736
rect 674281 797678 676260 797680
rect 674281 797675 674347 797678
rect 676254 797676 676260 797678
rect 676324 797676 676330 797740
rect 58065 793522 58131 793525
rect 58065 793520 64492 793522
rect 58065 793464 58070 793520
rect 58126 793464 64492 793520
rect 58065 793462 64492 793464
rect 58065 793459 58131 793462
rect 674189 792026 674255 792029
rect 676438 792026 676444 792028
rect 674189 792024 676444 792026
rect 674189 791968 674194 792024
rect 674250 791968 676444 792024
rect 674189 791966 676444 791968
rect 674189 791963 674255 791966
rect 676438 791964 676444 791966
rect 676508 791964 676514 792028
rect 655053 789986 655119 789989
rect 650164 789984 655119 789986
rect 650164 789928 655058 789984
rect 655114 789928 655119 789984
rect 650164 789926 655119 789928
rect 655053 789923 655119 789926
rect 674966 787748 674972 787812
rect 675036 787810 675042 787812
rect 675385 787810 675451 787813
rect 675036 787808 675451 787810
rect 675036 787752 675390 787808
rect 675446 787752 675451 787808
rect 675036 787750 675451 787752
rect 675036 787748 675042 787750
rect 675385 787747 675451 787750
rect 674598 787340 674604 787404
rect 674668 787402 674674 787404
rect 675385 787402 675451 787405
rect 674668 787400 675451 787402
rect 674668 787344 675390 787400
rect 675446 787344 675451 787400
rect 674668 787342 675451 787344
rect 674668 787340 674674 787342
rect 675385 787339 675451 787342
rect 675150 786796 675156 786860
rect 675220 786858 675226 786860
rect 675385 786858 675451 786861
rect 675220 786856 675451 786858
rect 675220 786800 675390 786856
rect 675446 786800 675451 786856
rect 675220 786798 675451 786800
rect 675220 786796 675226 786798
rect 675385 786795 675451 786798
rect 674782 784076 674788 784140
rect 674852 784138 674858 784140
rect 675385 784138 675451 784141
rect 674852 784136 675451 784138
rect 674852 784080 675390 784136
rect 675446 784080 675451 784136
rect 674852 784078 675451 784080
rect 674852 784076 674858 784078
rect 675385 784075 675451 784078
rect 674414 783804 674420 783868
rect 674484 783866 674490 783868
rect 675477 783866 675543 783869
rect 674484 783864 675543 783866
rect 674484 783808 675482 783864
rect 675538 783808 675543 783864
rect 674484 783806 675543 783808
rect 674484 783804 674490 783806
rect 675477 783803 675543 783806
rect 58433 780466 58499 780469
rect 58433 780464 64492 780466
rect 58433 780408 58438 780464
rect 58494 780408 64492 780464
rect 58433 780406 64492 780408
rect 58433 780403 58499 780406
rect 674230 777412 674236 777476
rect 674300 777474 674306 777476
rect 674373 777474 674439 777477
rect 674300 777472 674439 777474
rect 674300 777416 674378 777472
rect 674434 777416 674439 777472
rect 674300 777414 674439 777416
rect 674300 777412 674306 777414
rect 674373 777411 674439 777414
rect 655513 776658 655579 776661
rect 650164 776656 655579 776658
rect 650164 776600 655518 776656
rect 655574 776600 655579 776656
rect 650164 776598 655579 776600
rect 655513 776595 655579 776598
rect 41505 774754 41571 774757
rect 41462 774752 41571 774754
rect 41462 774696 41510 774752
rect 41566 774696 41571 774752
rect 41462 774691 41571 774696
rect 41462 774452 41522 774691
rect 41781 774074 41847 774077
rect 41492 774072 41847 774074
rect 41492 774016 41786 774072
rect 41842 774016 41847 774072
rect 41492 774014 41847 774016
rect 41781 774011 41847 774014
rect 41505 773938 41571 773941
rect 41462 773936 41571 773938
rect 41462 773880 41510 773936
rect 41566 773880 41571 773936
rect 41462 773875 41571 773880
rect 41462 773636 41522 773875
rect 41505 773530 41571 773533
rect 41462 773528 41571 773530
rect 41462 773472 41510 773528
rect 41566 773472 41571 773528
rect 41462 773467 41571 773472
rect 41462 773228 41522 773467
rect 39982 773060 39988 773124
rect 40052 773060 40058 773124
rect 39990 772820 40050 773060
rect 676806 772652 676812 772716
rect 676876 772714 676882 772716
rect 679065 772714 679131 772717
rect 676876 772712 679131 772714
rect 676876 772656 679070 772712
rect 679126 772656 679131 772712
rect 676876 772654 679131 772656
rect 676876 772652 676882 772654
rect 679065 772651 679131 772654
rect 43437 772442 43503 772445
rect 41492 772440 43503 772442
rect 41492 772384 43442 772440
rect 43498 772384 43503 772440
rect 41492 772382 43503 772384
rect 43437 772379 43503 772382
rect 42149 772034 42215 772037
rect 41492 772032 42215 772034
rect 41492 771976 42154 772032
rect 42210 771976 42215 772032
rect 41492 771974 42215 771976
rect 42149 771971 42215 771974
rect 39990 771492 40050 771596
rect 39982 771428 39988 771492
rect 40052 771428 40058 771492
rect 42885 771218 42951 771221
rect 41492 771216 42951 771218
rect 41492 771160 42890 771216
rect 42946 771160 42951 771216
rect 41492 771158 42951 771160
rect 42885 771155 42951 771158
rect 42425 770810 42491 770813
rect 41492 770808 42491 770810
rect 41492 770752 42430 770808
rect 42486 770752 42491 770808
rect 41492 770750 42491 770752
rect 42425 770747 42491 770750
rect 43529 770402 43595 770405
rect 41492 770400 43595 770402
rect 41492 770344 43534 770400
rect 43590 770344 43595 770400
rect 41492 770342 43595 770344
rect 43529 770339 43595 770342
rect 674189 770268 674255 770269
rect 674189 770266 674236 770268
rect 674144 770264 674236 770266
rect 674144 770208 674194 770264
rect 674144 770206 674236 770208
rect 674189 770204 674236 770206
rect 674300 770204 674306 770268
rect 674189 770203 674255 770204
rect 42701 769994 42767 769997
rect 41492 769992 42767 769994
rect 41492 769936 42706 769992
rect 42762 769936 42767 769992
rect 41492 769934 42767 769936
rect 42701 769931 42767 769934
rect 43069 769586 43135 769589
rect 41492 769584 43135 769586
rect 41492 769528 43074 769584
rect 43130 769528 43135 769584
rect 41492 769526 43135 769528
rect 43069 769523 43135 769526
rect 43713 769178 43779 769181
rect 41492 769176 43779 769178
rect 41492 769120 43718 769176
rect 43774 769120 43779 769176
rect 41492 769118 43779 769120
rect 43713 769115 43779 769118
rect 44081 768770 44147 768773
rect 41492 768768 44147 768770
rect 41492 768712 44086 768768
rect 44142 768712 44147 768768
rect 41492 768710 44147 768712
rect 44081 768707 44147 768710
rect 43161 768362 43227 768365
rect 41492 768360 43227 768362
rect 41492 768304 43166 768360
rect 43222 768304 43227 768360
rect 41492 768302 43227 768304
rect 43161 768299 43227 768302
rect 41873 767954 41939 767957
rect 41492 767952 41939 767954
rect 41492 767896 41878 767952
rect 41934 767896 41939 767952
rect 41492 767894 41939 767896
rect 41873 767891 41939 767894
rect 43253 767546 43319 767549
rect 41492 767544 43319 767546
rect 41492 767488 43258 767544
rect 43314 767488 43319 767544
rect 41492 767486 43319 767488
rect 43253 767483 43319 767486
rect 58433 767410 58499 767413
rect 58433 767408 64492 767410
rect 58433 767352 58438 767408
rect 58494 767352 64492 767408
rect 58433 767350 64492 767352
rect 58433 767347 58499 767350
rect 44081 767138 44147 767141
rect 41492 767136 44147 767138
rect 41492 767080 44086 767136
rect 44142 767080 44147 767136
rect 41492 767078 44147 767080
rect 44081 767075 44147 767078
rect 42057 766730 42123 766733
rect 41492 766728 42123 766730
rect 41492 766672 42062 766728
rect 42118 766672 42123 766728
rect 41492 766670 42123 766672
rect 42057 766667 42123 766670
rect 43161 766322 43227 766325
rect 41492 766320 43227 766322
rect 41492 766264 43166 766320
rect 43222 766264 43227 766320
rect 41492 766262 43227 766264
rect 43161 766259 43227 766262
rect 43529 765914 43595 765917
rect 41492 765912 43595 765914
rect 41492 765856 43534 765912
rect 43590 765856 43595 765912
rect 41492 765854 43595 765856
rect 43529 765851 43595 765854
rect 43989 765506 44055 765509
rect 41492 765504 44055 765506
rect 41492 765448 43994 765504
rect 44050 765448 44055 765504
rect 41492 765446 44055 765448
rect 43989 765443 44055 765446
rect 43437 765098 43503 765101
rect 41492 765096 43503 765098
rect 41492 765040 43442 765096
rect 43498 765040 43503 765096
rect 41492 765038 43503 765040
rect 43437 765035 43503 765038
rect 42885 764690 42951 764693
rect 41492 764688 42951 764690
rect 41492 764632 42890 764688
rect 42946 764632 42951 764688
rect 41492 764630 42951 764632
rect 42885 764627 42951 764630
rect 41462 764149 41522 764252
rect 41462 764144 41571 764149
rect 41462 764088 41510 764144
rect 41566 764088 41571 764144
rect 41462 764086 41571 764088
rect 41505 764083 41571 764086
rect 30422 763741 30482 763844
rect 30373 763736 30482 763741
rect 30373 763680 30378 763736
rect 30434 763680 30482 763736
rect 30373 763678 30482 763680
rect 30373 763675 30439 763678
rect 41462 763333 41522 763436
rect 30373 763330 30439 763333
rect 30373 763328 30482 763330
rect 30373 763272 30378 763328
rect 30434 763272 30482 763328
rect 30373 763267 30482 763272
rect 41462 763328 41571 763333
rect 654685 763330 654751 763333
rect 41462 763272 41510 763328
rect 41566 763272 41571 763328
rect 41462 763270 41571 763272
rect 650164 763328 654751 763330
rect 650164 763272 654690 763328
rect 654746 763272 654751 763328
rect 650164 763270 654751 763272
rect 41505 763267 41571 763270
rect 654685 763267 654751 763270
rect 30422 763028 30482 763267
rect 679022 761293 679082 761532
rect 678973 761288 679082 761293
rect 678973 761232 678978 761288
rect 679034 761232 679082 761288
rect 678973 761230 679082 761232
rect 678973 761227 679039 761230
rect 676262 760885 676322 761124
rect 676213 760880 676322 760885
rect 676213 760824 676218 760880
rect 676274 760824 676322 760880
rect 676213 760822 676322 760824
rect 676213 760819 676279 760822
rect 676121 760474 676187 760477
rect 676262 760474 676322 760716
rect 676121 760472 676322 760474
rect 676121 760416 676126 760472
rect 676182 760416 676322 760472
rect 676121 760414 676322 760416
rect 676121 760411 676187 760414
rect 673453 760338 673519 760341
rect 673862 760338 673868 760340
rect 673453 760336 673868 760338
rect 673453 760280 673458 760336
rect 673514 760280 673868 760336
rect 673453 760278 673868 760280
rect 673453 760275 673519 760278
rect 673862 760276 673868 760278
rect 673932 760338 673938 760340
rect 673932 760278 676292 760338
rect 673932 760276 673938 760278
rect 676262 759661 676322 759900
rect 676262 759656 676371 759661
rect 679065 759658 679131 759661
rect 676262 759600 676310 759656
rect 676366 759600 676371 759656
rect 676262 759598 676371 759600
rect 676305 759595 676371 759598
rect 679022 759656 679131 759658
rect 679022 759600 679070 759656
rect 679126 759600 679131 759656
rect 679022 759595 679131 759600
rect 679022 759492 679082 759595
rect 669773 759250 669839 759253
rect 673453 759250 673519 759253
rect 669773 759248 673519 759250
rect 669773 759192 669778 759248
rect 669834 759192 673458 759248
rect 673514 759192 673519 759248
rect 669773 759190 673519 759192
rect 669773 759187 669839 759190
rect 673453 759187 673519 759190
rect 676029 759114 676095 759117
rect 676029 759112 676292 759114
rect 676029 759056 676034 759112
rect 676090 759056 676292 759112
rect 676029 759054 676292 759056
rect 676029 759051 676095 759054
rect 679022 758437 679082 758676
rect 678973 758432 679082 758437
rect 678973 758376 678978 758432
rect 679034 758376 679082 758432
rect 678973 758374 679082 758376
rect 678973 758371 679039 758374
rect 676121 758026 676187 758029
rect 676262 758026 676322 758268
rect 676121 758024 676322 758026
rect 676121 757968 676126 758024
rect 676182 757968 676322 758024
rect 676121 757966 676322 757968
rect 676121 757963 676187 757966
rect 676262 757621 676322 757860
rect 676262 757616 676371 757621
rect 676262 757560 676310 757616
rect 676366 757560 676371 757616
rect 676262 757558 676371 757560
rect 676305 757555 676371 757558
rect 676262 757213 676322 757452
rect 676213 757208 676322 757213
rect 676213 757152 676218 757208
rect 676274 757152 676322 757208
rect 676213 757150 676322 757152
rect 676213 757147 676279 757150
rect 41965 757076 42031 757077
rect 41965 757072 42012 757076
rect 42076 757074 42082 757076
rect 41965 757016 41970 757072
rect 41965 757012 42012 757016
rect 42076 757014 42122 757074
rect 42076 757012 42082 757014
rect 675334 757012 675340 757076
rect 675404 757074 675410 757076
rect 675404 757014 676292 757074
rect 675404 757012 675410 757014
rect 41965 757011 42031 757012
rect 676029 756666 676095 756669
rect 676029 756664 676292 756666
rect 676029 756608 676034 756664
rect 676090 756608 676292 756664
rect 676029 756606 676292 756608
rect 676029 756603 676095 756606
rect 676070 756332 676076 756396
rect 676140 756394 676146 756396
rect 676140 756334 676322 756394
rect 676140 756332 676146 756334
rect 676262 756228 676322 756334
rect 675518 755788 675524 755852
rect 675588 755850 675594 755852
rect 675588 755790 676292 755850
rect 675588 755788 675594 755790
rect 676121 755578 676187 755581
rect 676121 755576 676322 755578
rect 676121 755520 676126 755576
rect 676182 755520 676322 755576
rect 676121 755518 676322 755520
rect 676121 755515 676187 755518
rect 676262 755412 676322 755518
rect 676029 755034 676095 755037
rect 676029 755032 676292 755034
rect 676029 754976 676034 755032
rect 676090 754976 676292 755032
rect 676029 754974 676292 754976
rect 676029 754971 676095 754974
rect 675702 754564 675708 754628
rect 675772 754626 675778 754628
rect 675772 754566 676292 754626
rect 675772 754564 675778 754566
rect 58341 754354 58407 754357
rect 58341 754352 64492 754354
rect 58341 754296 58346 754352
rect 58402 754296 64492 754352
rect 58341 754294 64492 754296
rect 58341 754291 58407 754294
rect 676029 754218 676095 754221
rect 676029 754216 676292 754218
rect 676029 754160 676034 754216
rect 676090 754160 676292 754216
rect 676029 754158 676292 754160
rect 676029 754155 676095 754158
rect 42057 754084 42123 754085
rect 42006 754020 42012 754084
rect 42076 754082 42123 754084
rect 42076 754080 42168 754082
rect 42118 754024 42168 754080
rect 42076 754022 42168 754024
rect 42076 754020 42123 754022
rect 42057 754019 42123 754020
rect 675569 753810 675635 753813
rect 675569 753808 676292 753810
rect 675569 753752 675574 753808
rect 675630 753752 676292 753808
rect 675569 753750 676292 753752
rect 675569 753747 675635 753750
rect 676029 753402 676095 753405
rect 676029 753400 676292 753402
rect 676029 753344 676034 753400
rect 676090 753344 676292 753400
rect 676029 753342 676292 753344
rect 676029 753339 676095 753342
rect 676029 752994 676095 752997
rect 676029 752992 676292 752994
rect 676029 752936 676034 752992
rect 676090 752936 676292 752992
rect 676029 752934 676292 752936
rect 676029 752931 676095 752934
rect 675886 752524 675892 752588
rect 675956 752586 675962 752588
rect 675956 752526 676292 752586
rect 675956 752524 675962 752526
rect 676438 752252 676444 752316
rect 676508 752252 676514 752316
rect 676446 752148 676506 752252
rect 676254 751844 676260 751908
rect 676324 751844 676330 751908
rect 676262 751740 676322 751844
rect 679206 751093 679266 751332
rect 679206 751088 679315 751093
rect 679206 751032 679254 751088
rect 679310 751032 679315 751088
rect 679206 751030 679315 751032
rect 679249 751027 679315 751030
rect 679022 750685 679082 750924
rect 678973 750680 679082 750685
rect 679249 750682 679315 750685
rect 678973 750624 678978 750680
rect 679034 750624 679082 750680
rect 678973 750622 679082 750624
rect 679206 750680 679315 750682
rect 679206 750624 679254 750680
rect 679310 750624 679315 750680
rect 678973 750619 679039 750622
rect 679206 750619 679315 750624
rect 679206 750516 679266 750619
rect 678973 750274 679039 750277
rect 678973 750272 679082 750274
rect 678973 750216 678978 750272
rect 679034 750216 679082 750272
rect 678973 750211 679082 750216
rect 654685 750138 654751 750141
rect 650164 750136 654751 750138
rect 650164 750080 654690 750136
rect 654746 750080 654751 750136
rect 679022 750108 679082 750211
rect 650164 750078 654751 750080
rect 654685 750075 654751 750078
rect 675477 744154 675543 744157
rect 676622 744154 676628 744156
rect 675477 744152 676628 744154
rect 675477 744096 675482 744152
rect 675538 744096 676628 744152
rect 675477 744094 676628 744096
rect 675477 744091 675543 744094
rect 676622 744092 676628 744094
rect 676692 744092 676698 744156
rect 675661 744018 675727 744021
rect 676254 744018 676260 744020
rect 675661 744016 676260 744018
rect 675661 743960 675666 744016
rect 675722 743960 676260 744016
rect 675661 743958 676260 743960
rect 675661 743955 675727 743958
rect 676254 743956 676260 743958
rect 676324 743956 676330 744020
rect 675753 742930 675819 742933
rect 675886 742930 675892 742932
rect 675753 742928 675892 742930
rect 675753 742872 675758 742928
rect 675814 742872 675892 742928
rect 675753 742870 675892 742872
rect 675753 742867 675819 742870
rect 675886 742868 675892 742870
rect 675956 742868 675962 742932
rect 675753 742522 675819 742525
rect 676070 742522 676076 742524
rect 675753 742520 676076 742522
rect 675753 742464 675758 742520
rect 675814 742464 676076 742520
rect 675753 742462 676076 742464
rect 675753 742459 675819 742462
rect 676070 742460 676076 742462
rect 676140 742460 676146 742524
rect 674230 741644 674236 741708
rect 674300 741706 674306 741708
rect 675477 741706 675543 741709
rect 674300 741704 675543 741706
rect 674300 741648 675482 741704
rect 675538 741648 675543 741704
rect 674300 741646 675543 741648
rect 674300 741644 674306 741646
rect 675477 741643 675543 741646
rect 58433 741298 58499 741301
rect 58433 741296 64492 741298
rect 58433 741240 58438 741296
rect 58494 741240 64492 741296
rect 58433 741238 64492 741240
rect 58433 741235 58499 741238
rect 675385 739804 675451 739805
rect 675334 739802 675340 739804
rect 675294 739742 675340 739802
rect 675404 739800 675451 739804
rect 675446 739744 675451 739800
rect 675334 739740 675340 739742
rect 675404 739740 675451 739744
rect 675385 739739 675451 739740
rect 673862 739060 673868 739124
rect 673932 739122 673938 739124
rect 675385 739122 675451 739125
rect 673932 739120 675451 739122
rect 673932 739064 675390 739120
rect 675446 739064 675451 739120
rect 673932 739062 675451 739064
rect 673932 739060 673938 739062
rect 675385 739059 675451 739062
rect 675661 738580 675727 738581
rect 675661 738576 675708 738580
rect 675772 738578 675778 738580
rect 675661 738520 675666 738576
rect 675661 738516 675708 738520
rect 675772 738518 675818 738578
rect 675772 738516 675778 738518
rect 675661 738515 675727 738516
rect 675753 738034 675819 738037
rect 676438 738034 676444 738036
rect 675753 738032 676444 738034
rect 675753 737976 675758 738032
rect 675814 737976 676444 738032
rect 675753 737974 676444 737976
rect 675753 737971 675819 737974
rect 676438 737972 676444 737974
rect 676508 737972 676514 738036
rect 654133 736810 654199 736813
rect 650164 736808 654199 736810
rect 650164 736752 654138 736808
rect 654194 736752 654199 736808
rect 650164 736750 654199 736752
rect 654133 736747 654199 736750
rect 41781 731370 41847 731373
rect 41492 731368 41847 731370
rect 41492 731312 41786 731368
rect 41842 731312 41847 731368
rect 41492 731310 41847 731312
rect 41781 731307 41847 731310
rect 39389 731098 39455 731101
rect 39982 731098 39988 731100
rect 39389 731096 39988 731098
rect 39389 731040 39394 731096
rect 39450 731040 39988 731096
rect 39389 731038 39988 731040
rect 39389 731035 39455 731038
rect 39982 731036 39988 731038
rect 40052 731036 40058 731100
rect 41505 731098 41571 731101
rect 41462 731096 41571 731098
rect 41462 731040 41510 731096
rect 41566 731040 41571 731096
rect 41462 731035 41571 731040
rect 41462 730932 41522 731035
rect 41505 730690 41571 730693
rect 41462 730688 41571 730690
rect 41462 730632 41510 730688
rect 41566 730632 41571 730688
rect 41462 730627 41571 730632
rect 41462 730524 41522 730627
rect 42793 730146 42859 730149
rect 44173 730146 44239 730149
rect 41492 730144 44239 730146
rect 41492 730088 42798 730144
rect 42854 730088 44178 730144
rect 44234 730088 44239 730144
rect 41492 730086 44239 730088
rect 42793 730083 42859 730086
rect 44173 730083 44239 730086
rect 39389 729874 39455 729877
rect 63217 729874 63283 729877
rect 39389 729872 63283 729874
rect 39389 729816 39394 729872
rect 39450 729816 63222 729872
rect 63278 729816 63283 729872
rect 39389 729814 63283 729816
rect 39389 729811 39455 729814
rect 63217 729811 63283 729814
rect 43345 729738 43411 729741
rect 41492 729736 43411 729738
rect 41492 729680 43350 729736
rect 43406 729680 43411 729736
rect 41492 729678 43411 729680
rect 43345 729675 43411 729678
rect 41505 729466 41571 729469
rect 41462 729464 41571 729466
rect 41462 729408 41510 729464
rect 41566 729408 41571 729464
rect 41462 729403 41571 729408
rect 41462 729300 41522 729403
rect 41781 728922 41847 728925
rect 41492 728920 41847 728922
rect 41492 728864 41786 728920
rect 41842 728864 41847 728920
rect 41492 728862 41847 728864
rect 41781 728859 41847 728862
rect 43713 728514 43779 728517
rect 44030 728514 44036 728516
rect 41492 728512 44036 728514
rect 41492 728456 43718 728512
rect 43774 728456 44036 728512
rect 41492 728454 44036 728456
rect 43713 728451 43779 728454
rect 44030 728452 44036 728454
rect 44100 728452 44106 728516
rect 39389 728242 39455 728245
rect 58433 728242 58499 728245
rect 39389 728240 39498 728242
rect 39389 728184 39394 728240
rect 39450 728184 39498 728240
rect 39389 728179 39498 728184
rect 58433 728240 64492 728242
rect 58433 728184 58438 728240
rect 58494 728184 64492 728240
rect 58433 728182 64492 728184
rect 58433 728179 58499 728182
rect 39438 728076 39498 728179
rect 44357 727698 44423 727701
rect 41492 727696 44423 727698
rect 41492 727640 44362 727696
rect 44418 727640 44423 727696
rect 41492 727638 44423 727640
rect 44357 727635 44423 727638
rect 42517 727290 42583 727293
rect 41492 727288 42583 727290
rect 41492 727232 42522 727288
rect 42578 727232 42583 727288
rect 41492 727230 42583 727232
rect 42517 727227 42583 727230
rect 43621 726882 43687 726885
rect 41492 726880 43687 726882
rect 41492 726824 43626 726880
rect 43682 726824 43687 726880
rect 41492 726822 43687 726824
rect 43621 726819 43687 726822
rect 43069 726474 43135 726477
rect 41492 726472 43135 726474
rect 41492 726416 43074 726472
rect 43130 726416 43135 726472
rect 41492 726414 43135 726416
rect 43069 726411 43135 726414
rect 43161 726066 43227 726069
rect 41492 726064 43227 726066
rect 41492 726008 43166 726064
rect 43222 726008 43227 726064
rect 41492 726006 43227 726008
rect 43161 726003 43227 726006
rect 43529 725658 43595 725661
rect 41492 725656 43595 725658
rect 41492 725600 43534 725656
rect 43590 725600 43595 725656
rect 41492 725598 43595 725600
rect 43529 725595 43595 725598
rect 43345 725250 43411 725253
rect 41492 725248 43411 725250
rect 41492 725192 43350 725248
rect 43406 725192 43411 725248
rect 41492 725190 43411 725192
rect 43345 725187 43411 725190
rect 41873 724842 41939 724845
rect 41492 724840 41939 724842
rect 41492 724784 41878 724840
rect 41934 724784 41939 724840
rect 41492 724782 41939 724784
rect 41873 724779 41939 724782
rect 42885 724434 42951 724437
rect 41492 724432 42951 724434
rect 41492 724376 42890 724432
rect 42946 724376 42951 724432
rect 41492 724374 42951 724376
rect 42885 724371 42951 724374
rect 41278 723757 41338 723996
rect 41278 723752 41387 723757
rect 41278 723696 41326 723752
rect 41382 723696 41387 723752
rect 41278 723694 41387 723696
rect 41321 723691 41387 723694
rect 42977 723618 43043 723621
rect 41492 723616 43043 723618
rect 41492 723560 42982 723616
rect 43038 723560 43043 723616
rect 41492 723558 43043 723560
rect 42977 723555 43043 723558
rect 655513 723482 655579 723485
rect 650164 723480 655579 723482
rect 650164 723424 655518 723480
rect 655574 723424 655579 723480
rect 650164 723422 655579 723424
rect 655513 723419 655579 723422
rect 42793 723210 42859 723213
rect 41492 723208 42859 723210
rect 41492 723152 42798 723208
rect 42854 723152 42859 723208
rect 41492 723150 42859 723152
rect 42793 723147 42859 723150
rect 43437 722802 43503 722805
rect 41492 722800 43503 722802
rect 41492 722744 43442 722800
rect 43498 722744 43503 722800
rect 41492 722742 43503 722744
rect 43437 722739 43503 722742
rect 43897 722394 43963 722397
rect 41492 722392 43963 722394
rect 41492 722336 43902 722392
rect 43958 722336 43963 722392
rect 41492 722334 43963 722336
rect 43897 722331 43963 722334
rect 44081 721986 44147 721989
rect 41492 721984 44147 721986
rect 41492 721928 44086 721984
rect 44142 721928 44147 721984
rect 41492 721926 44147 721928
rect 44081 721923 44147 721926
rect 43253 721578 43319 721581
rect 41492 721576 43319 721578
rect 41492 721520 43258 721576
rect 43314 721520 43319 721576
rect 41492 721518 43319 721520
rect 43253 721515 43319 721518
rect 41462 720901 41522 721140
rect 41462 720896 41571 720901
rect 41462 720840 41510 720896
rect 41566 720840 41571 720896
rect 41462 720838 41571 720840
rect 41505 720835 41571 720838
rect 30422 720493 30482 720732
rect 30373 720488 30482 720493
rect 30373 720432 30378 720488
rect 30434 720432 30482 720488
rect 30373 720430 30482 720432
rect 30373 720427 30439 720430
rect 41462 720085 41522 720324
rect 30373 720082 30439 720085
rect 30373 720080 30482 720082
rect 30373 720024 30378 720080
rect 30434 720024 30482 720080
rect 30373 720019 30482 720024
rect 41462 720080 41571 720085
rect 41462 720024 41510 720080
rect 41566 720024 41571 720080
rect 41462 720022 41571 720024
rect 41505 720019 41571 720022
rect 30422 719916 30482 720019
rect 676029 716546 676095 716549
rect 676029 716544 676292 716546
rect 676029 716488 676034 716544
rect 676090 716488 676292 716544
rect 676029 716486 676292 716488
rect 676029 716483 676095 716486
rect 676029 716138 676095 716141
rect 676029 716136 676292 716138
rect 676029 716080 676034 716136
rect 676090 716080 676292 716136
rect 676029 716078 676292 716080
rect 676029 716075 676095 716078
rect 676029 715730 676095 715733
rect 676029 715728 676292 715730
rect 676029 715672 676034 715728
rect 676090 715672 676292 715728
rect 676029 715670 676292 715672
rect 676029 715667 676095 715670
rect 58433 715322 58499 715325
rect 676029 715322 676095 715325
rect 58433 715320 64492 715322
rect 58433 715264 58438 715320
rect 58494 715264 64492 715320
rect 58433 715262 64492 715264
rect 676029 715320 676292 715322
rect 676029 715264 676034 715320
rect 676090 715264 676292 715320
rect 676029 715262 676292 715264
rect 58433 715259 58499 715262
rect 676029 715259 676095 715262
rect 676029 714914 676095 714917
rect 676029 714912 676292 714914
rect 676029 714856 676034 714912
rect 676090 714856 676292 714912
rect 676029 714854 676292 714856
rect 676029 714851 676095 714854
rect 678973 714506 679039 714509
rect 678973 714504 679052 714506
rect 678973 714448 678978 714504
rect 679034 714448 679052 714504
rect 678973 714446 679052 714448
rect 678973 714443 679039 714446
rect 676029 714098 676095 714101
rect 676029 714096 676292 714098
rect 676029 714040 676034 714096
rect 676090 714040 676292 714096
rect 676029 714038 676292 714040
rect 676029 714035 676095 714038
rect 676029 713690 676095 713693
rect 676029 713688 676292 713690
rect 676029 713632 676034 713688
rect 676090 713632 676292 713688
rect 676029 713630 676292 713632
rect 676029 713627 676095 713630
rect 676029 713282 676095 713285
rect 676029 713280 676292 713282
rect 676029 713224 676034 713280
rect 676090 713224 676292 713280
rect 676029 713222 676292 713224
rect 676029 713219 676095 713222
rect 676029 712874 676095 712877
rect 676029 712872 676292 712874
rect 676029 712816 676034 712872
rect 676090 712816 676292 712872
rect 676029 712814 676292 712816
rect 676029 712811 676095 712814
rect 676029 712466 676095 712469
rect 676029 712464 676292 712466
rect 676029 712408 676034 712464
rect 676090 712408 676292 712464
rect 676029 712406 676292 712408
rect 676029 712403 676095 712406
rect 675150 711996 675156 712060
rect 675220 712058 675226 712060
rect 675220 711998 676292 712058
rect 675220 711996 675226 711998
rect 675845 711650 675911 711653
rect 675845 711648 676292 711650
rect 675845 711592 675850 711648
rect 675906 711592 676292 711648
rect 675845 711590 676292 711592
rect 675845 711587 675911 711590
rect 674966 711180 674972 711244
rect 675036 711242 675042 711244
rect 675036 711182 676292 711242
rect 675036 711180 675042 711182
rect 676029 710834 676095 710837
rect 676029 710832 676292 710834
rect 676029 710776 676034 710832
rect 676090 710776 676292 710832
rect 676029 710774 676292 710776
rect 676029 710771 676095 710774
rect 676581 710598 676647 710599
rect 676254 710596 676260 710598
rect 675845 710562 675911 710565
rect 676078 710562 676260 710596
rect 675845 710560 676260 710562
rect 675845 710504 675850 710560
rect 675906 710536 676260 710560
rect 675906 710504 676138 710536
rect 676254 710534 676260 710536
rect 676324 710534 676330 710598
rect 676581 710594 676628 710598
rect 676692 710596 676698 710598
rect 676581 710538 676586 710594
rect 676581 710534 676628 710538
rect 676692 710536 676738 710596
rect 676692 710534 676698 710536
rect 676581 710533 676647 710534
rect 675845 710502 676138 710504
rect 675845 710499 675911 710502
rect 675937 710426 676003 710429
rect 675937 710424 676292 710426
rect 675937 710368 675942 710424
rect 675998 710368 676292 710424
rect 675937 710366 676292 710368
rect 675937 710363 676003 710366
rect 655973 710290 656039 710293
rect 650164 710288 656039 710290
rect 650164 710232 655978 710288
rect 656034 710232 656039 710288
rect 650164 710230 656039 710232
rect 655973 710227 656039 710230
rect 676029 710018 676095 710021
rect 676029 710016 676292 710018
rect 676029 709960 676034 710016
rect 676090 709960 676292 710016
rect 676029 709958 676292 709960
rect 676029 709955 676095 709958
rect 674598 709548 674604 709612
rect 674668 709610 674674 709612
rect 674668 709550 676292 709610
rect 674668 709548 674674 709550
rect 674782 709140 674788 709204
rect 674852 709202 674858 709204
rect 674852 709142 676292 709202
rect 674852 709140 674858 709142
rect 674414 708732 674420 708796
rect 674484 708794 674490 708796
rect 674484 708734 676292 708794
rect 674484 708732 674490 708734
rect 676029 708386 676095 708389
rect 676029 708384 676292 708386
rect 676029 708328 676034 708384
rect 676090 708328 676292 708384
rect 676029 708326 676292 708328
rect 676029 708323 676095 708326
rect 676029 707978 676095 707981
rect 676029 707976 676292 707978
rect 676029 707920 676034 707976
rect 676090 707920 676292 707976
rect 676029 707918 676292 707920
rect 676029 707915 676095 707918
rect 676029 707570 676095 707573
rect 676029 707568 676292 707570
rect 676029 707512 676034 707568
rect 676090 707512 676292 707568
rect 676029 707510 676292 707512
rect 676029 707507 676095 707510
rect 675845 707162 675911 707165
rect 675845 707160 676292 707162
rect 675845 707104 675850 707160
rect 675906 707104 676292 707160
rect 675845 707102 676292 707104
rect 675845 707099 675911 707102
rect 676029 706754 676095 706757
rect 676029 706752 676292 706754
rect 676029 706696 676034 706752
rect 676090 706696 676292 706752
rect 676029 706694 676292 706696
rect 676029 706691 676095 706694
rect 675937 706346 676003 706349
rect 675937 706344 676292 706346
rect 675937 706288 675942 706344
rect 675998 706288 676292 706344
rect 675937 706286 676292 706288
rect 675937 706283 676003 706286
rect 676029 705938 676095 705941
rect 676029 705936 676292 705938
rect 676029 705880 676034 705936
rect 676090 705880 676292 705936
rect 676029 705878 676292 705880
rect 676029 705875 676095 705878
rect 675937 705530 676003 705533
rect 675937 705528 676292 705530
rect 675937 705472 675942 705528
rect 675998 705472 676292 705528
rect 675937 705470 676292 705472
rect 675937 705467 676003 705470
rect 676029 705122 676095 705125
rect 676029 705120 676292 705122
rect 676029 705064 676034 705120
rect 676090 705064 676292 705120
rect 676029 705062 676292 705064
rect 676029 705059 676095 705062
rect 58157 702266 58223 702269
rect 58157 702264 64492 702266
rect 58157 702208 58162 702264
rect 58218 702208 64492 702264
rect 58157 702206 64492 702208
rect 58157 702203 58223 702206
rect 673637 699818 673703 699821
rect 676254 699818 676260 699820
rect 673637 699816 676260 699818
rect 673637 699760 673642 699816
rect 673698 699760 676260 699816
rect 673637 699758 676260 699760
rect 673637 699755 673703 699758
rect 676254 699756 676260 699758
rect 676324 699756 676330 699820
rect 674005 699682 674071 699685
rect 676806 699682 676812 699684
rect 674005 699680 676812 699682
rect 674005 699624 674010 699680
rect 674066 699624 676812 699680
rect 674005 699622 676812 699624
rect 674005 699619 674071 699622
rect 676806 699620 676812 699622
rect 676876 699620 676882 699684
rect 675661 699546 675727 699549
rect 676990 699546 676996 699548
rect 675661 699544 676996 699546
rect 675661 699488 675666 699544
rect 675722 699488 676996 699544
rect 675661 699486 676996 699488
rect 675661 699483 675727 699486
rect 676990 699484 676996 699486
rect 677060 699484 677066 699548
rect 675477 698188 675543 698189
rect 675477 698184 675524 698188
rect 675588 698186 675594 698188
rect 675477 698128 675482 698184
rect 675477 698124 675524 698128
rect 675588 698126 675634 698186
rect 675588 698124 675594 698126
rect 675477 698123 675543 698124
rect 673678 697308 673684 697372
rect 673748 697370 673754 697372
rect 675385 697370 675451 697373
rect 673748 697368 675451 697370
rect 673748 697312 675390 697368
rect 675446 697312 675451 697368
rect 673748 697310 675451 697312
rect 673748 697308 673754 697310
rect 675385 697307 675451 697310
rect 654869 696962 654935 696965
rect 650164 696960 654935 696962
rect 650164 696904 654874 696960
rect 654930 696904 654935 696960
rect 650164 696902 654935 696904
rect 654869 696899 654935 696902
rect 674414 696628 674420 696692
rect 674484 696690 674490 696692
rect 675385 696690 675451 696693
rect 674484 696688 675451 696690
rect 674484 696632 675390 696688
rect 675446 696632 675451 696688
rect 674484 696630 675451 696632
rect 674484 696628 674490 696630
rect 675385 696627 675451 696630
rect 674598 694724 674604 694788
rect 674668 694786 674674 694788
rect 675385 694786 675451 694789
rect 674668 694784 675451 694786
rect 674668 694728 675390 694784
rect 675446 694728 675451 694784
rect 674668 694726 675451 694728
rect 674668 694724 674674 694726
rect 675385 694723 675451 694726
rect 673494 694316 673500 694380
rect 673564 694378 673570 694380
rect 675477 694378 675543 694381
rect 673564 694376 675543 694378
rect 673564 694320 675482 694376
rect 675538 694320 675543 694376
rect 673564 694318 675543 694320
rect 673564 694316 673570 694318
rect 675477 694315 675543 694318
rect 674046 693500 674052 693564
rect 674116 693562 674122 693564
rect 675385 693562 675451 693565
rect 674116 693560 675451 693562
rect 674116 693504 675390 693560
rect 675446 693504 675451 693560
rect 674116 693502 675451 693504
rect 674116 693500 674122 693502
rect 675385 693499 675451 693502
rect 675753 693018 675819 693021
rect 677174 693018 677180 693020
rect 675753 693016 677180 693018
rect 675753 692960 675758 693016
rect 675814 692960 677180 693016
rect 675753 692958 677180 692960
rect 675753 692955 675819 692958
rect 677174 692956 677180 692958
rect 677244 692956 677250 693020
rect 675753 690162 675819 690165
rect 676622 690162 676628 690164
rect 675753 690160 676628 690162
rect 675753 690104 675758 690160
rect 675814 690104 676628 690160
rect 675753 690102 676628 690104
rect 675753 690099 675819 690102
rect 676622 690100 676628 690102
rect 676692 690100 676698 690164
rect 58433 689210 58499 689213
rect 58433 689208 64492 689210
rect 58433 689152 58438 689208
rect 58494 689152 64492 689208
rect 58433 689150 64492 689152
rect 58433 689147 58499 689150
rect 41505 688394 41571 688397
rect 41462 688392 41571 688394
rect 41462 688336 41510 688392
rect 41566 688336 41571 688392
rect 41462 688331 41571 688336
rect 41462 688092 41522 688331
rect 41781 687714 41847 687717
rect 41492 687712 41847 687714
rect 41492 687656 41786 687712
rect 41842 687656 41847 687712
rect 41492 687654 41847 687656
rect 41781 687651 41847 687654
rect 41689 687578 41755 687581
rect 41462 687576 41755 687578
rect 41462 687520 41694 687576
rect 41750 687520 41755 687576
rect 41462 687518 41755 687520
rect 41462 687276 41522 687518
rect 41689 687515 41755 687518
rect 41278 686764 41338 686868
rect 41270 686700 41276 686764
rect 41340 686700 41346 686764
rect 44173 686490 44239 686493
rect 41492 686488 44239 686490
rect 41492 686432 44178 686488
rect 44234 686432 44239 686488
rect 41492 686430 44239 686432
rect 44173 686427 44239 686430
rect 44265 686082 44331 686085
rect 41492 686080 44331 686082
rect 41492 686024 44270 686080
rect 44326 686024 44331 686080
rect 41492 686022 44331 686024
rect 44265 686019 44331 686022
rect 43437 685674 43503 685677
rect 41492 685672 43503 685674
rect 41492 685616 43442 685672
rect 43498 685616 43503 685672
rect 41492 685614 43503 685616
rect 43437 685611 43503 685614
rect 42793 685266 42859 685269
rect 41492 685264 42859 685266
rect 41492 685208 42798 685264
rect 42854 685208 42859 685264
rect 41492 685206 42859 685208
rect 42793 685203 42859 685206
rect 43161 684858 43227 684861
rect 41492 684856 43227 684858
rect 41492 684800 43166 684856
rect 43222 684800 43227 684856
rect 41492 684798 43227 684800
rect 43161 684795 43227 684798
rect 42885 684450 42951 684453
rect 41492 684448 42951 684450
rect 41492 684392 42890 684448
rect 42946 684392 42951 684448
rect 41492 684390 42951 684392
rect 42885 684387 42951 684390
rect 39982 684252 39988 684316
rect 40052 684314 40058 684316
rect 41638 684314 41644 684316
rect 40052 684254 41644 684314
rect 40052 684252 40058 684254
rect 41638 684252 41644 684254
rect 41708 684314 41714 684316
rect 62573 684314 62639 684317
rect 41708 684312 62639 684314
rect 41708 684256 62578 684312
rect 62634 684256 62639 684312
rect 41708 684254 62639 684256
rect 41708 684252 41714 684254
rect 62573 684251 62639 684254
rect 44030 684042 44036 684044
rect 41492 683982 44036 684042
rect 44030 683980 44036 683982
rect 44100 684042 44106 684044
rect 44357 684042 44423 684045
rect 44100 684040 44423 684042
rect 44100 683984 44362 684040
rect 44418 683984 44423 684040
rect 44100 683982 44423 683984
rect 44100 683980 44106 683982
rect 44357 683979 44423 683982
rect 43345 683634 43411 683637
rect 654133 683634 654199 683637
rect 41492 683632 43411 683634
rect 41492 683576 43350 683632
rect 43406 683576 43411 683632
rect 41492 683574 43411 683576
rect 650164 683632 654199 683634
rect 650164 683576 654138 683632
rect 654194 683576 654199 683632
rect 650164 683574 654199 683576
rect 43345 683571 43411 683574
rect 654133 683571 654199 683574
rect 43989 683226 44055 683229
rect 41492 683224 44055 683226
rect 41492 683168 43994 683224
rect 44050 683168 44055 683224
rect 41492 683166 44055 683168
rect 43989 683163 44055 683166
rect 42977 682818 43043 682821
rect 41492 682816 43043 682818
rect 41492 682760 42982 682816
rect 43038 682760 43043 682816
rect 41492 682758 43043 682760
rect 42977 682755 43043 682758
rect 43805 682410 43871 682413
rect 41492 682408 43871 682410
rect 41492 682352 43810 682408
rect 43866 682352 43871 682408
rect 41492 682350 43871 682352
rect 43805 682347 43871 682350
rect 41462 681866 41522 681972
rect 41689 681866 41755 681869
rect 41462 681864 41755 681866
rect 41462 681808 41694 681864
rect 41750 681808 41755 681864
rect 41462 681806 41755 681808
rect 41689 681803 41755 681806
rect 41873 681594 41939 681597
rect 41492 681592 41939 681594
rect 41492 681536 41878 681592
rect 41934 681536 41939 681592
rect 41492 681534 41939 681536
rect 41873 681531 41939 681534
rect 43713 681186 43779 681189
rect 41492 681184 43779 681186
rect 41492 681128 43718 681184
rect 43774 681128 43779 681184
rect 41492 681126 43779 681128
rect 43713 681123 43779 681126
rect 43161 680778 43227 680781
rect 41492 680776 43227 680778
rect 41492 680720 43166 680776
rect 43222 680720 43227 680776
rect 41492 680718 43227 680720
rect 43161 680715 43227 680718
rect 43621 680370 43687 680373
rect 41492 680368 43687 680370
rect 41492 680312 43626 680368
rect 43682 680312 43687 680368
rect 41492 680310 43687 680312
rect 43621 680307 43687 680310
rect 43897 679962 43963 679965
rect 41492 679960 43963 679962
rect 41492 679904 43902 679960
rect 43958 679904 43963 679960
rect 41492 679902 43963 679904
rect 43897 679899 43963 679902
rect 43529 679554 43595 679557
rect 41492 679552 43595 679554
rect 41492 679496 43534 679552
rect 43590 679496 43595 679552
rect 41492 679494 43595 679496
rect 43529 679491 43595 679494
rect 44081 679146 44147 679149
rect 41492 679144 44147 679146
rect 41492 679088 44086 679144
rect 44142 679088 44147 679144
rect 41492 679086 44147 679088
rect 44081 679083 44147 679086
rect 41781 678738 41847 678741
rect 41492 678736 41847 678738
rect 41492 678680 41786 678736
rect 41842 678680 41847 678736
rect 41492 678678 41847 678680
rect 41781 678675 41847 678678
rect 41965 678330 42031 678333
rect 41492 678328 42031 678330
rect 41492 678272 41970 678328
rect 42026 678272 42031 678328
rect 41492 678270 42031 678272
rect 41965 678267 42031 678270
rect 41781 677922 41847 677925
rect 41492 677920 41847 677922
rect 41492 677864 41786 677920
rect 41842 677864 41847 677920
rect 41492 677862 41847 677864
rect 41781 677859 41847 677862
rect 30606 677380 30666 677484
rect 30598 677316 30604 677380
rect 30668 677316 30674 677380
rect 41781 677106 41847 677109
rect 41492 677104 41847 677106
rect 41492 677048 41786 677104
rect 41842 677048 41847 677104
rect 41492 677046 41847 677048
rect 41781 677043 41847 677046
rect 30598 676908 30604 676972
rect 30668 676908 30674 676972
rect 30606 676668 30666 676908
rect 58433 676154 58499 676157
rect 58433 676152 64492 676154
rect 58433 676096 58438 676152
rect 58494 676096 64492 676152
rect 58433 676094 64492 676096
rect 58433 676091 58499 676094
rect 676262 671125 676322 671364
rect 676213 671120 676322 671125
rect 676213 671064 676218 671120
rect 676274 671064 676322 671120
rect 676213 671062 676322 671064
rect 676213 671059 676279 671062
rect 676029 670986 676095 670989
rect 676029 670984 676292 670986
rect 676029 670928 676034 670984
rect 676090 670928 676292 670984
rect 676029 670926 676292 670928
rect 676029 670923 676095 670926
rect 676029 670578 676095 670581
rect 676029 670576 676292 670578
rect 676029 670520 676034 670576
rect 676090 670520 676292 670576
rect 676029 670518 676292 670520
rect 676029 670515 676095 670518
rect 655513 670442 655579 670445
rect 650164 670440 655579 670442
rect 650164 670384 655518 670440
rect 655574 670384 655579 670440
rect 650164 670382 655579 670384
rect 655513 670379 655579 670382
rect 676213 670306 676279 670309
rect 676213 670304 676322 670306
rect 676213 670248 676218 670304
rect 676274 670248 676322 670304
rect 676213 670243 676322 670248
rect 676262 670140 676322 670243
rect 676029 669762 676095 669765
rect 676029 669760 676292 669762
rect 676029 669704 676034 669760
rect 676090 669704 676292 669760
rect 676029 669702 676292 669704
rect 676029 669699 676095 669702
rect 678973 669490 679039 669493
rect 678973 669488 679082 669490
rect 678973 669432 678978 669488
rect 679034 669432 679082 669488
rect 678973 669427 679082 669432
rect 679022 669324 679082 669427
rect 676029 668946 676095 668949
rect 676029 668944 676292 668946
rect 676029 668888 676034 668944
rect 676090 668888 676292 668944
rect 676029 668886 676292 668888
rect 676029 668883 676095 668886
rect 676213 668674 676279 668677
rect 676213 668672 676322 668674
rect 676213 668616 676218 668672
rect 676274 668616 676322 668672
rect 676213 668611 676322 668616
rect 676262 668508 676322 668611
rect 675937 668130 676003 668133
rect 675937 668128 676292 668130
rect 675937 668072 675942 668128
rect 675998 668072 676292 668128
rect 675937 668070 676292 668072
rect 675937 668067 676003 668070
rect 675937 667722 676003 667725
rect 675937 667720 676292 667722
rect 675937 667664 675942 667720
rect 675998 667664 676292 667720
rect 675937 667662 676292 667664
rect 675937 667659 676003 667662
rect 668761 667314 668827 667317
rect 668761 667312 677580 667314
rect 668761 667256 668766 667312
rect 668822 667284 677580 667312
rect 668822 667256 677610 667284
rect 668761 667254 677610 667256
rect 668761 667251 668827 667254
rect 677550 667044 677610 667254
rect 677542 666980 677548 667044
rect 677612 666980 677618 667044
rect 674230 666844 674236 666908
rect 674300 666906 674306 666908
rect 674300 666846 676292 666906
rect 674300 666844 674306 666846
rect 676121 666634 676187 666637
rect 676121 666632 676322 666634
rect 676121 666576 676126 666632
rect 676182 666576 676322 666632
rect 676121 666574 676322 666576
rect 676121 666571 676187 666574
rect 676262 666468 676322 666574
rect 675886 666028 675892 666092
rect 675956 666090 675962 666092
rect 675956 666030 676292 666090
rect 675956 666028 675962 666030
rect 675334 665620 675340 665684
rect 675404 665682 675410 665684
rect 675404 665622 676292 665682
rect 675404 665620 675410 665622
rect 676029 665274 676095 665277
rect 676029 665272 676292 665274
rect 676029 665216 676034 665272
rect 676090 665216 676292 665272
rect 676029 665214 676292 665216
rect 676029 665211 676095 665214
rect 676121 665002 676187 665005
rect 676121 665000 676322 665002
rect 676121 664944 676126 665000
rect 676182 664944 676322 665000
rect 676121 664942 676322 664944
rect 676121 664939 676187 664942
rect 676262 664836 676322 664942
rect 676070 664532 676076 664596
rect 676140 664594 676146 664596
rect 676140 664534 676322 664594
rect 676140 664532 676146 664534
rect 676262 664428 676322 664534
rect 673862 663988 673868 664052
rect 673932 664050 673938 664052
rect 673932 663990 676292 664050
rect 673932 663988 673938 663990
rect 675702 663580 675708 663644
rect 675772 663642 675778 663644
rect 675772 663582 676292 663642
rect 675772 663580 675778 663582
rect 676029 663234 676095 663237
rect 676029 663232 676292 663234
rect 676029 663176 676034 663232
rect 676090 663176 676292 663232
rect 676029 663174 676292 663176
rect 676029 663171 676095 663174
rect 58433 663098 58499 663101
rect 58433 663096 64492 663098
rect 58433 663040 58438 663096
rect 58494 663040 64492 663096
rect 58433 663038 64492 663040
rect 58433 663035 58499 663038
rect 676254 662900 676260 662964
rect 676324 662900 676330 662964
rect 676262 662796 676322 662900
rect 676438 662492 676444 662556
rect 676508 662492 676514 662556
rect 676446 662388 676506 662492
rect 676990 662084 676996 662148
rect 677060 662084 677066 662148
rect 676998 661980 677058 662084
rect 676806 661676 676812 661740
rect 676876 661676 676882 661740
rect 676814 661572 676874 661676
rect 679022 660925 679082 661164
rect 678973 660920 679082 660925
rect 678973 660864 678978 660920
rect 679034 660864 679082 660920
rect 678973 660862 679082 660864
rect 678973 660859 679039 660862
rect 684542 660517 684602 660756
rect 678973 660514 679039 660517
rect 678973 660512 679082 660514
rect 678973 660456 678978 660512
rect 679034 660456 679082 660512
rect 678973 660451 679082 660456
rect 684493 660512 684602 660517
rect 684493 660456 684498 660512
rect 684554 660456 684602 660512
rect 684493 660454 684602 660456
rect 684493 660451 684559 660454
rect 679022 660348 679082 660451
rect 684493 660106 684559 660109
rect 684493 660104 684602 660106
rect 684493 660048 684498 660104
rect 684554 660048 684602 660104
rect 684493 660043 684602 660048
rect 684542 659940 684602 660043
rect 656801 657114 656867 657117
rect 650164 657112 656867 657114
rect 650164 657056 656806 657112
rect 656862 657056 656867 657112
rect 650164 657054 656867 657056
rect 656801 657051 656867 657054
rect 674966 652836 674972 652900
rect 675036 652898 675042 652900
rect 675385 652898 675451 652901
rect 675036 652896 675451 652898
rect 675036 652840 675390 652896
rect 675446 652840 675451 652896
rect 675036 652838 675451 652840
rect 675036 652836 675042 652838
rect 675385 652835 675451 652838
rect 674782 652156 674788 652220
rect 674852 652218 674858 652220
rect 675477 652218 675543 652221
rect 674852 652216 675543 652218
rect 674852 652160 675482 652216
rect 675538 652160 675543 652216
rect 674852 652158 675543 652160
rect 674852 652156 674858 652158
rect 675477 652155 675543 652158
rect 675150 651612 675156 651676
rect 675220 651674 675226 651676
rect 675385 651674 675451 651677
rect 675220 651672 675451 651674
rect 675220 651616 675390 651672
rect 675446 651616 675451 651672
rect 675220 651614 675451 651616
rect 675220 651612 675226 651614
rect 675385 651611 675451 651614
rect 59169 650042 59235 650045
rect 59169 650040 64492 650042
rect 59169 649984 59174 650040
rect 59230 649984 64492 650040
rect 59169 649982 64492 649984
rect 59169 649979 59235 649982
rect 675385 648956 675451 648957
rect 675334 648954 675340 648956
rect 675294 648894 675340 648954
rect 675404 648952 675451 648956
rect 675446 648896 675451 648952
rect 675334 648892 675340 648894
rect 675404 648892 675451 648896
rect 675385 648891 675451 648892
rect 675753 648682 675819 648685
rect 675886 648682 675892 648684
rect 675753 648680 675892 648682
rect 675753 648624 675758 648680
rect 675814 648624 675892 648680
rect 675753 648622 675892 648624
rect 675753 648619 675819 648622
rect 675886 648620 675892 648622
rect 675956 648620 675962 648684
rect 41505 645146 41571 645149
rect 41462 645144 41571 645146
rect 41462 645088 41510 645144
rect 41566 645088 41571 645144
rect 41462 645083 41571 645088
rect 41462 644912 41522 645083
rect 41505 644738 41571 644741
rect 41462 644736 41571 644738
rect 41462 644680 41510 644736
rect 41566 644680 41571 644736
rect 41462 644675 41571 644680
rect 41462 644504 41522 644675
rect 41505 644330 41571 644333
rect 41462 644328 41571 644330
rect 41462 644272 41510 644328
rect 41566 644272 41571 644328
rect 41462 644267 41571 644272
rect 41462 644096 41522 644267
rect 654869 643786 654935 643789
rect 650164 643784 654935 643786
rect 650164 643728 654874 643784
rect 654930 643728 654935 643784
rect 650164 643726 654935 643728
rect 654869 643723 654935 643726
rect 41462 643517 41522 643688
rect 39982 643452 39988 643516
rect 40052 643452 40058 643516
rect 41462 643512 41571 643517
rect 41462 643456 41510 643512
rect 41566 643456 41571 643512
rect 41462 643454 41571 643456
rect 39990 643280 40050 643452
rect 41505 643451 41571 643454
rect 43437 643106 43503 643109
rect 41462 643104 43503 643106
rect 41462 643048 43442 643104
rect 43498 643048 43503 643104
rect 41462 643046 43503 643048
rect 41462 642872 41522 643046
rect 43437 643043 43503 643046
rect 41462 642290 41522 642464
rect 44449 642290 44515 642293
rect 41462 642288 44515 642290
rect 41462 642232 44454 642288
rect 44510 642232 44515 642288
rect 41462 642230 44515 642232
rect 44449 642227 44515 642230
rect 41462 642018 41522 642056
rect 44265 642018 44331 642021
rect 41462 642016 44331 642018
rect 41462 641960 44270 642016
rect 44326 641960 44331 642016
rect 41462 641958 44331 641960
rect 44265 641955 44331 641958
rect 42793 641882 42859 641885
rect 41462 641880 42859 641882
rect 41462 641824 42798 641880
rect 42854 641824 42859 641880
rect 41462 641822 42859 641824
rect 41462 641648 41522 641822
rect 42793 641819 42859 641822
rect 44633 641474 44699 641477
rect 46473 641474 46539 641477
rect 41462 641472 46539 641474
rect 41462 641416 44638 641472
rect 44694 641416 46478 641472
rect 46534 641416 46539 641472
rect 41462 641414 46539 641416
rect 41462 641240 41522 641414
rect 44633 641411 44699 641414
rect 46473 641411 46539 641414
rect 42885 641066 42951 641069
rect 41462 641064 42951 641066
rect 41462 641008 42890 641064
rect 42946 641008 42951 641064
rect 41462 641006 42951 641008
rect 41462 640832 41522 641006
rect 42885 641003 42951 641006
rect 41462 640386 41522 640424
rect 43069 640386 43135 640389
rect 41462 640384 43135 640386
rect 41462 640328 43074 640384
rect 43130 640328 43135 640384
rect 41462 640326 43135 640328
rect 43069 640323 43135 640326
rect 41462 639842 41522 640016
rect 43529 639842 43595 639845
rect 41462 639840 43595 639842
rect 41462 639784 43534 639840
rect 43590 639784 43595 639840
rect 41462 639782 43595 639784
rect 43529 639779 43595 639782
rect 41462 639434 41522 639608
rect 42793 639434 42859 639437
rect 41462 639432 42859 639434
rect 41462 639376 42798 639432
rect 42854 639376 42859 639432
rect 41462 639374 42859 639376
rect 42793 639371 42859 639374
rect 41462 639026 41522 639200
rect 43161 639026 43227 639029
rect 41462 639024 43227 639026
rect 41462 638968 43166 639024
rect 43222 638968 43227 639024
rect 41462 638966 43227 638968
rect 43161 638963 43227 638966
rect 41462 638618 41522 638792
rect 43437 638618 43503 638621
rect 41462 638616 43503 638618
rect 41462 638560 43442 638616
rect 43498 638560 43503 638616
rect 41462 638558 43503 638560
rect 43437 638555 43503 638558
rect 41781 638414 41847 638417
rect 41492 638412 41847 638414
rect 41492 638356 41786 638412
rect 41842 638356 41847 638412
rect 41492 638354 41847 638356
rect 41781 638351 41847 638354
rect 41462 637802 41522 637976
rect 42977 637802 43043 637805
rect 41462 637800 43043 637802
rect 41462 637744 42982 637800
rect 43038 637744 43043 637800
rect 41462 637742 43043 637744
rect 42977 637739 43043 637742
rect 43713 637666 43779 637669
rect 41462 637664 43779 637666
rect 41462 637608 43718 637664
rect 43774 637608 43779 637664
rect 41462 637606 43779 637608
rect 41462 637568 41522 637606
rect 43713 637603 43779 637606
rect 41462 636986 41522 637160
rect 58433 637122 58499 637125
rect 58433 637120 64492 637122
rect 58433 637064 58438 637120
rect 58494 637064 64492 637120
rect 58433 637062 64492 637064
rect 58433 637059 58499 637062
rect 43805 636986 43871 636989
rect 41462 636984 43871 636986
rect 41462 636928 43810 636984
rect 43866 636928 43871 636984
rect 41462 636926 43871 636928
rect 43805 636923 43871 636926
rect 41462 636578 41522 636752
rect 42885 636578 42951 636581
rect 41462 636576 42951 636578
rect 41462 636520 42890 636576
rect 42946 636520 42951 636576
rect 41462 636518 42951 636520
rect 42885 636515 42951 636518
rect 41462 636170 41522 636344
rect 43345 636170 43411 636173
rect 41462 636168 43411 636170
rect 41462 636112 43350 636168
rect 43406 636112 43411 636168
rect 41462 636110 43411 636112
rect 43345 636107 43411 636110
rect 41462 635762 41522 635936
rect 43621 635762 43687 635765
rect 41462 635760 43687 635762
rect 41462 635704 43626 635760
rect 43682 635704 43687 635760
rect 41462 635702 43687 635704
rect 43621 635699 43687 635702
rect 41462 635354 41522 635528
rect 43253 635354 43319 635357
rect 41462 635352 43319 635354
rect 41462 635296 43258 635352
rect 43314 635296 43319 635352
rect 41462 635294 43319 635296
rect 43253 635291 43319 635294
rect 32998 634949 33058 635120
rect 32998 634944 33107 634949
rect 32998 634888 33046 634944
rect 33102 634888 33107 634944
rect 32998 634886 33107 634888
rect 33041 634883 33107 634886
rect 41462 634541 41522 634712
rect 41462 634536 41571 634541
rect 41462 634480 41510 634536
rect 41566 634480 41571 634536
rect 41462 634478 41571 634480
rect 41505 634475 41571 634478
rect 30422 634133 30482 634304
rect 30373 634128 30482 634133
rect 30373 634072 30378 634128
rect 30434 634072 30482 634128
rect 30373 634070 30482 634072
rect 30373 634067 30439 634070
rect 41462 633725 41522 633896
rect 30373 633722 30439 633725
rect 30373 633720 30482 633722
rect 30373 633664 30378 633720
rect 30434 633664 30482 633720
rect 30373 633659 30482 633664
rect 41462 633720 41571 633725
rect 41462 633664 41510 633720
rect 41566 633664 41571 633720
rect 41462 633662 41571 633664
rect 41505 633659 41571 633662
rect 30422 633488 30482 633659
rect 654133 630594 654199 630597
rect 650164 630592 654199 630594
rect 650164 630536 654138 630592
rect 654194 630536 654199 630592
rect 650164 630534 654199 630536
rect 654133 630531 654199 630534
rect 679022 626109 679082 626348
rect 678973 626104 679082 626109
rect 678973 626048 678978 626104
rect 679034 626048 679082 626104
rect 678973 626046 679082 626048
rect 678973 626043 679039 626046
rect 676121 625698 676187 625701
rect 676262 625698 676322 625940
rect 676121 625696 676322 625698
rect 676121 625640 676126 625696
rect 676182 625640 676322 625696
rect 676121 625638 676322 625640
rect 676121 625635 676187 625638
rect 676262 625293 676322 625532
rect 676262 625288 676371 625293
rect 676262 625232 676310 625288
rect 676366 625232 676371 625288
rect 676262 625230 676371 625232
rect 676305 625227 676371 625230
rect 676029 625154 676095 625157
rect 676029 625152 676292 625154
rect 676029 625096 676034 625152
rect 676090 625096 676292 625152
rect 676029 625094 676292 625096
rect 676029 625091 676095 625094
rect 676262 624477 676322 624716
rect 676213 624472 676322 624477
rect 679065 624474 679131 624477
rect 676213 624416 676218 624472
rect 676274 624416 676322 624472
rect 676213 624414 676322 624416
rect 679022 624472 679131 624474
rect 679022 624416 679070 624472
rect 679126 624416 679131 624472
rect 676213 624411 676279 624414
rect 679022 624411 679131 624416
rect 679022 624308 679082 624411
rect 58433 624066 58499 624069
rect 58433 624064 64492 624066
rect 58433 624008 58438 624064
rect 58494 624008 64492 624064
rect 58433 624006 64492 624008
rect 58433 624003 58499 624006
rect 676029 623930 676095 623933
rect 676029 623928 676292 623930
rect 676029 623872 676034 623928
rect 676090 623872 676292 623928
rect 676029 623870 676292 623872
rect 676029 623867 676095 623870
rect 679157 623658 679223 623661
rect 679022 623656 679223 623658
rect 679022 623600 679162 623656
rect 679218 623600 679223 623656
rect 679022 623598 679223 623600
rect 679022 623253 679082 623598
rect 679157 623595 679223 623598
rect 678973 623248 679082 623253
rect 678973 623192 678978 623248
rect 679034 623192 679082 623248
rect 678973 623190 679082 623192
rect 678973 623187 679039 623190
rect 673862 623052 673868 623116
rect 673932 623114 673938 623116
rect 673932 623054 676292 623114
rect 673932 623052 673938 623054
rect 677358 622780 677364 622844
rect 677428 622780 677434 622844
rect 677366 622676 677426 622780
rect 676262 622029 676322 622268
rect 676213 622024 676322 622029
rect 676213 621968 676218 622024
rect 676274 621968 676322 622024
rect 676213 621966 676322 621968
rect 676213 621963 676279 621966
rect 674414 621828 674420 621892
rect 674484 621890 674490 621892
rect 674484 621830 676292 621890
rect 674484 621828 674490 621830
rect 668669 621618 668735 621621
rect 673862 621618 673868 621620
rect 668669 621616 673868 621618
rect 668669 621560 668674 621616
rect 668730 621560 673868 621616
rect 668669 621558 673868 621560
rect 668669 621555 668735 621558
rect 673862 621556 673868 621558
rect 673932 621556 673938 621620
rect 676029 621482 676095 621485
rect 676029 621480 676292 621482
rect 676029 621424 676034 621480
rect 676090 621424 676292 621480
rect 676029 621422 676292 621424
rect 676029 621419 676095 621422
rect 675518 621012 675524 621076
rect 675588 621074 675594 621076
rect 675588 621014 676292 621074
rect 675588 621012 675594 621014
rect 674598 620604 674604 620668
rect 674668 620666 674674 620668
rect 674668 620606 676292 620666
rect 674668 620604 674674 620606
rect 676121 620394 676187 620397
rect 676121 620392 676322 620394
rect 676121 620336 676126 620392
rect 676182 620336 676322 620392
rect 676121 620334 676322 620336
rect 676121 620331 676187 620334
rect 676262 620228 676322 620334
rect 676029 619850 676095 619853
rect 676029 619848 676292 619850
rect 676029 619792 676034 619848
rect 676090 619792 676292 619848
rect 676029 619790 676292 619792
rect 676029 619787 676095 619790
rect 673678 619380 673684 619444
rect 673748 619442 673754 619444
rect 673748 619382 676292 619442
rect 673748 619380 673754 619382
rect 673494 618972 673500 619036
rect 673564 619034 673570 619036
rect 673564 618974 676292 619034
rect 673564 618972 673570 618974
rect 674046 618564 674052 618628
rect 674116 618626 674122 618628
rect 674116 618566 676292 618626
rect 674116 618564 674122 618566
rect 676029 618218 676095 618221
rect 676029 618216 676292 618218
rect 676029 618160 676034 618216
rect 676090 618160 676292 618216
rect 676029 618158 676292 618160
rect 676029 618155 676095 618158
rect 676213 617946 676279 617949
rect 676213 617944 676322 617946
rect 676213 617888 676218 617944
rect 676274 617888 676322 617944
rect 676213 617883 676322 617888
rect 676262 617780 676322 617883
rect 677174 617476 677180 617540
rect 677244 617476 677250 617540
rect 677182 617372 677242 617476
rect 654593 617266 654659 617269
rect 650164 617264 654659 617266
rect 650164 617208 654598 617264
rect 654654 617208 654659 617264
rect 650164 617206 654659 617208
rect 654593 617203 654659 617206
rect 676622 617068 676628 617132
rect 676692 617068 676698 617132
rect 676630 616964 676690 617068
rect 676213 616722 676279 616725
rect 676213 616720 676322 616722
rect 676213 616664 676218 616720
rect 676274 616664 676322 616720
rect 676213 616659 676322 616664
rect 676262 616556 676322 616659
rect 679206 615909 679266 616148
rect 679206 615904 679315 615909
rect 679206 615848 679254 615904
rect 679310 615848 679315 615904
rect 679206 615846 679315 615848
rect 679249 615843 679315 615846
rect 679022 615501 679082 615740
rect 678973 615496 679082 615501
rect 679249 615498 679315 615501
rect 678973 615440 678978 615496
rect 679034 615440 679082 615496
rect 678973 615438 679082 615440
rect 679206 615496 679315 615498
rect 679206 615440 679254 615496
rect 679310 615440 679315 615496
rect 678973 615435 679039 615438
rect 679206 615435 679315 615440
rect 679206 615332 679266 615435
rect 678973 615090 679039 615093
rect 678973 615088 679082 615090
rect 678973 615032 678978 615088
rect 679034 615032 679082 615088
rect 678973 615027 679082 615032
rect 679022 614924 679082 615027
rect 58433 611010 58499 611013
rect 58433 611008 64492 611010
rect 58433 610952 58438 611008
rect 58494 610952 64492 611008
rect 58433 610950 64492 610952
rect 58433 610947 58499 610950
rect 674373 608970 674439 608973
rect 676438 608970 676444 608972
rect 674373 608968 676444 608970
rect 674373 608912 674378 608968
rect 674434 608912 676444 608968
rect 674373 608910 676444 608912
rect 674373 608907 674439 608910
rect 676438 608908 676444 608910
rect 676508 608908 676514 608972
rect 675477 608834 675543 608837
rect 676622 608834 676628 608836
rect 675477 608832 676628 608834
rect 675477 608776 675482 608832
rect 675538 608776 676628 608832
rect 675477 608774 676628 608776
rect 675477 608771 675543 608774
rect 676622 608772 676628 608774
rect 676692 608772 676698 608836
rect 675661 607612 675727 607613
rect 675661 607608 675708 607612
rect 675772 607610 675778 607612
rect 675661 607552 675666 607608
rect 675661 607548 675708 607552
rect 675772 607550 675818 607610
rect 675772 607548 675778 607550
rect 675661 607547 675727 607548
rect 675753 607338 675819 607341
rect 676070 607338 676076 607340
rect 675753 607336 676076 607338
rect 675753 607280 675758 607336
rect 675814 607280 676076 607336
rect 675753 607278 676076 607280
rect 675753 607275 675819 607278
rect 676070 607276 676076 607278
rect 676140 607276 676146 607340
rect 674598 606460 674604 606524
rect 674668 606522 674674 606524
rect 675385 606522 675451 606525
rect 674668 606520 675451 606522
rect 674668 606464 675390 606520
rect 675446 606464 675451 606520
rect 674668 606462 675451 606464
rect 674668 606460 674674 606462
rect 675385 606459 675451 606462
rect 674414 604692 674420 604756
rect 674484 604754 674490 604756
rect 675385 604754 675451 604757
rect 674484 604752 675451 604754
rect 674484 604696 675390 604752
rect 675446 604696 675451 604752
rect 674484 604694 675451 604696
rect 674484 604692 674490 604694
rect 675385 604691 675451 604694
rect 675477 604348 675543 604349
rect 675477 604344 675524 604348
rect 675588 604346 675594 604348
rect 675477 604288 675482 604344
rect 675477 604284 675524 604288
rect 675588 604286 675634 604346
rect 675588 604284 675594 604286
rect 675477 604283 675543 604284
rect 654317 603938 654383 603941
rect 650164 603936 654383 603938
rect 650164 603880 654322 603936
rect 654378 603880 654383 603936
rect 650164 603878 654383 603880
rect 654317 603875 654383 603878
rect 674230 603468 674236 603532
rect 674300 603530 674306 603532
rect 675477 603530 675543 603533
rect 674300 603528 675543 603530
rect 674300 603472 675482 603528
rect 675538 603472 675543 603528
rect 674300 603470 675543 603472
rect 674300 603468 674306 603470
rect 675477 603467 675543 603470
rect 675753 602986 675819 602989
rect 676254 602986 676260 602988
rect 675753 602984 676260 602986
rect 675753 602928 675758 602984
rect 675814 602928 676260 602984
rect 675753 602926 676260 602928
rect 675753 602923 675819 602926
rect 676254 602924 676260 602926
rect 676324 602924 676330 602988
rect 41505 601898 41571 601901
rect 41462 601896 41571 601898
rect 41462 601840 41510 601896
rect 41566 601840 41571 601896
rect 41462 601835 41571 601840
rect 41462 601732 41522 601835
rect 41505 601490 41571 601493
rect 41462 601488 41571 601490
rect 41462 601432 41510 601488
rect 41566 601432 41571 601488
rect 41462 601427 41571 601432
rect 41462 601324 41522 601427
rect 53833 600946 53899 600949
rect 41492 600944 53899 600946
rect 41492 600888 53838 600944
rect 53894 600888 53899 600944
rect 41492 600886 53899 600888
rect 53833 600883 53899 600886
rect 43069 600538 43135 600541
rect 43846 600538 43852 600540
rect 41492 600536 43852 600538
rect 41492 600480 43074 600536
rect 43130 600480 43852 600536
rect 41492 600478 43852 600480
rect 43069 600475 43135 600478
rect 43846 600476 43852 600478
rect 43916 600476 43922 600540
rect 44357 600130 44423 600133
rect 46473 600130 46539 600133
rect 41492 600128 46539 600130
rect 41492 600072 44362 600128
rect 44418 600072 46478 600128
rect 46534 600072 46539 600128
rect 41492 600070 46539 600072
rect 44357 600067 44423 600070
rect 46473 600067 46539 600070
rect 41505 599858 41571 599861
rect 41462 599856 41571 599858
rect 41462 599800 41510 599856
rect 41566 599800 41571 599856
rect 41462 599795 41571 599800
rect 41462 599692 41522 599795
rect 41462 599045 41522 599284
rect 41462 599040 41571 599045
rect 41462 598984 41510 599040
rect 41566 598984 41571 599040
rect 41462 598982 41571 598984
rect 41505 598979 41571 598982
rect 40174 598636 40234 598876
rect 40166 598572 40172 598636
rect 40236 598572 40242 598636
rect 44265 598498 44331 598501
rect 46565 598498 46631 598501
rect 41492 598496 46631 598498
rect 41492 598440 44270 598496
rect 44326 598440 46570 598496
rect 46626 598440 46631 598496
rect 41492 598438 46631 598440
rect 44265 598435 44331 598438
rect 46565 598435 46631 598438
rect 42425 598090 42491 598093
rect 43662 598090 43668 598092
rect 41492 598088 43668 598090
rect 41492 598032 42430 598088
rect 42486 598032 43668 598088
rect 41492 598030 43668 598032
rect 42425 598027 42491 598030
rect 43662 598028 43668 598030
rect 43732 598028 43738 598092
rect 59169 597954 59235 597957
rect 59169 597952 64492 597954
rect 59169 597896 59174 597952
rect 59230 597896 64492 597952
rect 59169 597894 64492 597896
rect 59169 597891 59235 597894
rect 44633 597682 44699 597685
rect 41492 597680 44699 597682
rect 41492 597624 44638 597680
rect 44694 597624 44699 597680
rect 41492 597622 44699 597624
rect 44633 597619 44699 597622
rect 43805 597274 43871 597277
rect 41492 597272 43871 597274
rect 41492 597216 43810 597272
rect 43866 597216 43871 597272
rect 41492 597214 43871 597216
rect 43805 597211 43871 597214
rect 42885 596866 42951 596869
rect 41492 596864 42951 596866
rect 41492 596808 42890 596864
rect 42946 596808 42951 596864
rect 41492 596806 42951 596808
rect 42885 596803 42951 596806
rect 43253 596458 43319 596461
rect 41492 596456 43319 596458
rect 41492 596400 43258 596456
rect 43314 596400 43319 596456
rect 41492 596398 43319 596400
rect 43253 596395 43319 596398
rect 40166 596124 40172 596188
rect 40236 596186 40242 596188
rect 62389 596186 62455 596189
rect 40236 596184 62455 596186
rect 40236 596128 62394 596184
rect 62450 596128 62455 596184
rect 40236 596126 62455 596128
rect 40236 596124 40242 596126
rect 62389 596123 62455 596126
rect 43897 596050 43963 596053
rect 41492 596048 43963 596050
rect 41492 595992 43902 596048
rect 43958 595992 43963 596048
rect 41492 595990 43963 595992
rect 43897 595987 43963 595990
rect 43437 595642 43503 595645
rect 41492 595640 43503 595642
rect 41492 595584 43442 595640
rect 43498 595584 43503 595640
rect 41492 595582 43503 595584
rect 43437 595579 43503 595582
rect 41873 595234 41939 595237
rect 41492 595232 41939 595234
rect 41492 595176 41878 595232
rect 41934 595176 41939 595232
rect 41492 595174 41939 595176
rect 41873 595171 41939 595174
rect 43161 594826 43227 594829
rect 41492 594824 43227 594826
rect 41492 594768 43166 594824
rect 43222 594768 43227 594824
rect 41492 594766 43227 594768
rect 43161 594763 43227 594766
rect 41278 594149 41338 594388
rect 41278 594144 41387 594149
rect 41278 594088 41326 594144
rect 41382 594088 41387 594144
rect 41278 594086 41387 594088
rect 41321 594083 41387 594086
rect 42977 594010 43043 594013
rect 41492 594008 43043 594010
rect 41492 593952 42982 594008
rect 43038 593952 43043 594008
rect 41492 593950 43043 593952
rect 42977 593947 43043 593950
rect 42793 593602 42859 593605
rect 41492 593600 42859 593602
rect 41492 593544 42798 593600
rect 42854 593544 42859 593600
rect 41492 593542 42859 593544
rect 42793 593539 42859 593542
rect 43621 593194 43687 593197
rect 41492 593192 43687 593194
rect 41492 593136 43626 593192
rect 43682 593136 43687 593192
rect 41492 593134 43687 593136
rect 43621 593131 43687 593134
rect 43713 592786 43779 592789
rect 41492 592784 43779 592786
rect 41492 592728 43718 592784
rect 43774 592728 43779 592784
rect 41492 592726 43779 592728
rect 43713 592723 43779 592726
rect 43253 592378 43319 592381
rect 41492 592376 43319 592378
rect 41492 592320 43258 592376
rect 43314 592320 43319 592376
rect 41492 592318 43319 592320
rect 43253 592315 43319 592318
rect 42701 591970 42767 591973
rect 41492 591968 42767 591970
rect 41492 591912 42706 591968
rect 42762 591912 42767 591968
rect 41492 591910 42767 591912
rect 42701 591907 42767 591910
rect 29870 591293 29930 591532
rect 29870 591288 29979 591293
rect 29870 591232 29918 591288
rect 29974 591232 29979 591288
rect 29870 591230 29979 591232
rect 29913 591227 29979 591230
rect 30422 590885 30482 591124
rect 29913 590882 29979 590885
rect 29870 590880 29979 590882
rect 29870 590824 29918 590880
rect 29974 590824 29979 590880
rect 29870 590819 29979 590824
rect 30373 590880 30482 590885
rect 30373 590824 30378 590880
rect 30434 590824 30482 590880
rect 30373 590822 30482 590824
rect 30373 590819 30439 590822
rect 29870 590716 29930 590819
rect 48865 590746 48931 590749
rect 656801 590746 656867 590749
rect 41492 590744 48931 590746
rect 41492 590688 48870 590744
rect 48926 590688 48931 590744
rect 41492 590686 48931 590688
rect 650164 590744 656867 590746
rect 650164 590688 656806 590744
rect 656862 590688 656867 590744
rect 650164 590686 656867 590688
rect 48865 590683 48931 590686
rect 656801 590683 656867 590686
rect 30373 590474 30439 590477
rect 30373 590472 30482 590474
rect 30373 590416 30378 590472
rect 30434 590416 30482 590472
rect 30373 590411 30482 590416
rect 30422 590308 30482 590411
rect 58433 584898 58499 584901
rect 58433 584896 64492 584898
rect 58433 584840 58438 584896
rect 58494 584840 64492 584896
rect 58433 584838 64492 584840
rect 58433 584835 58499 584838
rect 676121 580954 676187 580957
rect 676262 580954 676322 581060
rect 676121 580952 676322 580954
rect 676121 580896 676126 580952
rect 676182 580896 676322 580952
rect 676121 580894 676322 580896
rect 676121 580891 676187 580894
rect 676262 580549 676322 580652
rect 676262 580544 676371 580549
rect 676262 580488 676310 580544
rect 676366 580488 676371 580544
rect 676262 580486 676371 580488
rect 676305 580483 676371 580486
rect 676262 580141 676322 580244
rect 676213 580136 676322 580141
rect 676213 580080 676218 580136
rect 676274 580080 676322 580136
rect 676213 580078 676322 580080
rect 676213 580075 676279 580078
rect 676029 579866 676095 579869
rect 676029 579864 676292 579866
rect 676029 579808 676034 579864
rect 676090 579808 676292 579864
rect 676029 579806 676292 579808
rect 676029 579803 676095 579806
rect 676262 579325 676322 579428
rect 676213 579320 676322 579325
rect 676213 579264 676218 579320
rect 676274 579264 676322 579320
rect 676213 579262 676322 579264
rect 678973 579322 679039 579325
rect 678973 579320 679082 579322
rect 678973 579264 678978 579320
rect 679034 579264 679082 579320
rect 676213 579259 676279 579262
rect 678973 579259 679082 579264
rect 679022 579020 679082 579259
rect 676262 578509 676322 578612
rect 676213 578504 676322 578509
rect 676213 578448 676218 578504
rect 676274 578448 676322 578504
rect 676213 578446 676322 578448
rect 676213 578443 676279 578446
rect 673862 578172 673868 578236
rect 673932 578234 673938 578236
rect 673932 578174 676292 578234
rect 673932 578172 673938 578174
rect 676262 577693 676322 577796
rect 676213 577688 676322 577693
rect 676213 577632 676218 577688
rect 676274 577632 676322 577688
rect 676213 577630 676322 577632
rect 676213 577627 676279 577630
rect 654501 577418 654567 577421
rect 650164 577416 654567 577418
rect 650164 577360 654506 577416
rect 654562 577360 654567 577416
rect 650164 577358 654567 577360
rect 654501 577355 654567 577358
rect 676262 577285 676322 577388
rect 676213 577280 676322 577285
rect 676213 577224 676218 577280
rect 676274 577224 676322 577280
rect 676213 577222 676322 577224
rect 676213 577219 676279 577222
rect 676029 577010 676095 577013
rect 676029 577008 676292 577010
rect 676029 576952 676034 577008
rect 676090 576952 676292 577008
rect 676029 576950 676292 576952
rect 676029 576947 676095 576950
rect 675150 576540 675156 576604
rect 675220 576602 675226 576604
rect 675220 576542 676292 576602
rect 675220 576540 675226 576542
rect 676029 576194 676095 576197
rect 676029 576192 676292 576194
rect 676029 576136 676034 576192
rect 676090 576136 676292 576192
rect 676029 576134 676292 576136
rect 676029 576131 676095 576134
rect 674966 575724 674972 575788
rect 675036 575786 675042 575788
rect 675036 575726 676292 575786
rect 675036 575724 675042 575726
rect 675569 575378 675635 575381
rect 675569 575376 676292 575378
rect 675569 575320 675574 575376
rect 675630 575320 676292 575376
rect 675569 575318 676292 575320
rect 675569 575315 675635 575318
rect 676029 574970 676095 574973
rect 676029 574968 676292 574970
rect 676029 574912 676034 574968
rect 676090 574912 676292 574968
rect 676029 574910 676292 574912
rect 676029 574907 676095 574910
rect 675385 574562 675451 574565
rect 675385 574560 676292 574562
rect 675385 574504 675390 574560
rect 675446 574504 676292 574560
rect 675385 574502 676292 574504
rect 675385 574499 675451 574502
rect 674782 574092 674788 574156
rect 674852 574154 674858 574156
rect 674852 574094 676292 574154
rect 674852 574092 674858 574094
rect 675334 573684 675340 573748
rect 675404 573746 675410 573748
rect 675404 573686 676292 573746
rect 675404 573684 675410 573686
rect 675886 573276 675892 573340
rect 675956 573338 675962 573340
rect 675956 573278 676292 573338
rect 675956 573276 675962 573278
rect 676029 572930 676095 572933
rect 676029 572928 676292 572930
rect 676029 572872 676034 572928
rect 676090 572872 676292 572928
rect 676029 572870 676292 572872
rect 676029 572867 676095 572870
rect 676029 572522 676095 572525
rect 676029 572520 676292 572522
rect 676029 572464 676034 572520
rect 676090 572464 676292 572520
rect 676029 572462 676292 572464
rect 676029 572459 676095 572462
rect 676029 572114 676095 572117
rect 676029 572112 676292 572114
rect 676029 572056 676034 572112
rect 676090 572056 676292 572112
rect 676029 572054 676292 572056
rect 676029 572051 676095 572054
rect 676622 571916 676628 571980
rect 676692 571916 676698 571980
rect 58433 571842 58499 571845
rect 58433 571840 64492 571842
rect 58433 571784 58438 571840
rect 58494 571784 64492 571840
rect 58433 571782 64492 571784
rect 58433 571779 58499 571782
rect 676630 571676 676690 571916
rect 676438 571508 676444 571572
rect 676508 571508 676514 571572
rect 676446 571268 676506 571508
rect 679022 570757 679082 570860
rect 678973 570752 679082 570757
rect 678973 570696 678978 570752
rect 679034 570696 679082 570752
rect 678973 570694 679082 570696
rect 678973 570691 679039 570694
rect 684542 570349 684602 570452
rect 678973 570346 679039 570349
rect 678973 570344 679082 570346
rect 678973 570288 678978 570344
rect 679034 570288 679082 570344
rect 678973 570283 679082 570288
rect 684493 570344 684602 570349
rect 684493 570288 684498 570344
rect 684554 570288 684602 570344
rect 684493 570286 684602 570288
rect 684493 570283 684559 570286
rect 679022 570044 679082 570283
rect 684493 569938 684559 569941
rect 684493 569936 684602 569938
rect 684493 569880 684498 569936
rect 684554 569880 684602 569936
rect 684493 569875 684602 569880
rect 684542 569636 684602 569875
rect 675477 564498 675543 564501
rect 676806 564498 676812 564500
rect 675477 564496 676812 564498
rect 675477 564440 675482 564496
rect 675538 564440 676812 564496
rect 675477 564438 676812 564440
rect 675477 564435 675543 564438
rect 676806 564436 676812 564438
rect 676876 564436 676882 564500
rect 654317 564090 654383 564093
rect 650164 564088 654383 564090
rect 650164 564032 654322 564088
rect 654378 564032 654383 564088
rect 650164 564030 654383 564032
rect 654317 564027 654383 564030
rect 675334 562396 675340 562460
rect 675404 562458 675410 562460
rect 675477 562458 675543 562461
rect 675404 562456 675543 562458
rect 675404 562400 675482 562456
rect 675538 562400 675543 562456
rect 675404 562398 675543 562400
rect 675404 562396 675410 562398
rect 675477 562395 675543 562398
rect 675753 562050 675819 562053
rect 675886 562050 675892 562052
rect 675753 562048 675892 562050
rect 675753 561992 675758 562048
rect 675814 561992 675892 562048
rect 675753 561990 675892 561992
rect 675753 561987 675819 561990
rect 675886 561988 675892 561990
rect 675956 561988 675962 562052
rect 675150 561172 675156 561236
rect 675220 561234 675226 561236
rect 675477 561234 675543 561237
rect 675220 561232 675543 561234
rect 675220 561176 675482 561232
rect 675538 561176 675543 561232
rect 675220 561174 675543 561176
rect 675220 561172 675226 561174
rect 675477 561171 675543 561174
rect 41505 558786 41571 558789
rect 41462 558784 41571 558786
rect 41462 558728 41510 558784
rect 41566 558728 41571 558784
rect 41462 558723 41571 558728
rect 57973 558786 58039 558789
rect 57973 558784 64492 558786
rect 57973 558728 57978 558784
rect 58034 558728 64492 558784
rect 57973 558726 64492 558728
rect 57973 558723 58039 558726
rect 674966 558724 674972 558788
rect 675036 558786 675042 558788
rect 675385 558786 675451 558789
rect 675036 558784 675451 558786
rect 675036 558728 675390 558784
rect 675446 558728 675451 558784
rect 675036 558726 675451 558728
rect 675036 558724 675042 558726
rect 675385 558723 675451 558726
rect 41462 558484 41522 558723
rect 675753 558378 675819 558381
rect 676438 558378 676444 558380
rect 675753 558376 676444 558378
rect 675753 558320 675758 558376
rect 675814 558320 676444 558376
rect 675753 558318 676444 558320
rect 675753 558315 675819 558318
rect 676438 558316 676444 558318
rect 676508 558316 676514 558380
rect 41781 558106 41847 558109
rect 41492 558104 41847 558106
rect 41492 558048 41786 558104
rect 41842 558048 41847 558104
rect 41492 558046 41847 558048
rect 41781 558043 41847 558046
rect 41505 557970 41571 557973
rect 41462 557968 41571 557970
rect 41462 557912 41510 557968
rect 41566 557912 41571 557968
rect 41462 557907 41571 557912
rect 41462 557668 41522 557907
rect 675753 557562 675819 557565
rect 676622 557562 676628 557564
rect 675753 557560 676628 557562
rect 675753 557504 675758 557560
rect 675814 557504 676628 557560
rect 675753 557502 676628 557504
rect 675753 557499 675819 557502
rect 676622 557500 676628 557502
rect 676692 557500 676698 557564
rect 41462 557154 41522 557260
rect 41638 557154 41644 557156
rect 41462 557094 41644 557154
rect 41638 557092 41644 557094
rect 41708 557092 41714 557156
rect 43069 556882 43135 556885
rect 41492 556880 43135 556882
rect 41492 556824 43074 556880
rect 43130 556824 43135 556880
rect 41492 556822 43135 556824
rect 43069 556819 43135 556822
rect 43345 556474 43411 556477
rect 41492 556472 43411 556474
rect 41492 556416 43350 556472
rect 43406 556416 43411 556472
rect 41492 556414 43411 556416
rect 43345 556411 43411 556414
rect 43846 556066 43852 556068
rect 41492 556006 43852 556066
rect 43846 556004 43852 556006
rect 43916 556004 43922 556068
rect 39990 555524 40050 555628
rect 39982 555460 39988 555524
rect 40052 555460 40058 555524
rect 40166 555460 40172 555524
rect 40236 555460 40242 555524
rect 40174 555220 40234 555460
rect 41822 554842 41828 554844
rect 41492 554782 41828 554842
rect 41822 554780 41828 554782
rect 41892 554780 41898 554844
rect 43161 554434 43227 554437
rect 41492 554432 43227 554434
rect 41492 554376 43166 554432
rect 43222 554376 43227 554432
rect 41492 554374 43227 554376
rect 43161 554371 43227 554374
rect 43529 554026 43595 554029
rect 41492 554024 43595 554026
rect 41492 553968 43534 554024
rect 43590 553968 43595 554024
rect 41492 553966 43595 553968
rect 43529 553963 43595 553966
rect 42701 553618 42767 553621
rect 41492 553616 42767 553618
rect 41492 553560 42706 553616
rect 42762 553560 42767 553616
rect 41492 553558 42767 553560
rect 42701 553555 42767 553558
rect 43345 553210 43411 553213
rect 41492 553208 43411 553210
rect 41492 553152 43350 553208
rect 43406 553152 43411 553208
rect 41492 553150 43411 553152
rect 43345 553147 43411 553150
rect 42977 552802 43043 552805
rect 41492 552800 43043 552802
rect 41492 552744 42982 552800
rect 43038 552744 43043 552800
rect 41492 552742 43043 552744
rect 42977 552739 43043 552742
rect 43161 552394 43227 552397
rect 41492 552392 43227 552394
rect 41492 552336 43166 552392
rect 43222 552336 43227 552392
rect 41492 552334 43227 552336
rect 43161 552331 43227 552334
rect 41781 551986 41847 551989
rect 41492 551984 41847 551986
rect 41492 551928 41786 551984
rect 41842 551928 41847 551984
rect 41492 551926 41847 551928
rect 41781 551923 41847 551926
rect 43621 551578 43687 551581
rect 41492 551576 43687 551578
rect 41492 551520 43626 551576
rect 43682 551520 43687 551576
rect 41492 551518 43687 551520
rect 43621 551515 43687 551518
rect 43069 551170 43135 551173
rect 41492 551168 43135 551170
rect 41492 551112 43074 551168
rect 43130 551112 43135 551168
rect 41492 551110 43135 551112
rect 43069 551107 43135 551110
rect 655053 550898 655119 550901
rect 650164 550896 655119 550898
rect 650164 550840 655058 550896
rect 655114 550840 655119 550896
rect 650164 550838 655119 550840
rect 655053 550835 655119 550838
rect 43713 550762 43779 550765
rect 41492 550760 43779 550762
rect 41492 550704 43718 550760
rect 43774 550704 43779 550760
rect 41492 550702 43779 550704
rect 43713 550699 43779 550702
rect 42885 550354 42951 550357
rect 41492 550352 42951 550354
rect 41492 550296 42890 550352
rect 42946 550296 42951 550352
rect 41492 550294 42951 550296
rect 42885 550291 42951 550294
rect 43437 549946 43503 549949
rect 41492 549944 43503 549946
rect 41492 549888 43442 549944
rect 43498 549888 43503 549944
rect 41492 549886 43503 549888
rect 43437 549883 43503 549886
rect 43805 549538 43871 549541
rect 41492 549536 43871 549538
rect 41492 549480 43810 549536
rect 43866 549480 43871 549536
rect 41492 549478 43871 549480
rect 43805 549475 43871 549478
rect 41462 548994 41522 549100
rect 41597 548994 41663 548997
rect 41462 548992 41663 548994
rect 41462 548936 41602 548992
rect 41658 548936 41663 548992
rect 41462 548934 41663 548936
rect 41597 548931 41663 548934
rect 41462 548589 41522 548692
rect 41462 548584 41571 548589
rect 41462 548528 41510 548584
rect 41566 548528 41571 548584
rect 41462 548526 41571 548528
rect 41505 548523 41571 548526
rect 41462 548181 41522 548284
rect 41413 548176 41522 548181
rect 41413 548120 41418 548176
rect 41474 548120 41522 548176
rect 41413 548118 41522 548120
rect 41413 548115 41479 548118
rect 30422 547773 30482 547876
rect 30422 547768 30531 547773
rect 30422 547712 30470 547768
rect 30526 547712 30531 547768
rect 30422 547710 30531 547712
rect 30465 547707 30531 547710
rect 41462 547365 41522 547468
rect 30465 547362 30531 547365
rect 30422 547360 30531 547362
rect 30422 547304 30470 547360
rect 30526 547304 30531 547360
rect 30422 547299 30531 547304
rect 41413 547360 41522 547365
rect 41413 547304 41418 547360
rect 41474 547304 41522 547360
rect 41413 547302 41522 547304
rect 41413 547299 41479 547302
rect 30422 547060 30482 547299
rect 59169 545866 59235 545869
rect 59169 545864 64492 545866
rect 59169 545808 59174 545864
rect 59230 545808 64492 545864
rect 59169 545806 64492 545808
rect 59169 545803 59235 545806
rect 41822 540908 41828 540972
rect 41892 540970 41898 540972
rect 44081 540970 44147 540973
rect 41892 540968 44147 540970
rect 41892 540912 44086 540968
rect 44142 540912 44147 540968
rect 41892 540910 44147 540912
rect 41892 540908 41898 540910
rect 44081 540907 44147 540910
rect 41638 540772 41644 540836
rect 41708 540834 41714 540836
rect 43989 540834 44055 540837
rect 41708 540832 44055 540834
rect 41708 540776 43994 540832
rect 44050 540776 44055 540832
rect 41708 540774 44055 540776
rect 41708 540772 41714 540774
rect 43989 540771 44055 540774
rect 654685 537570 654751 537573
rect 650164 537568 654751 537570
rect 650164 537512 654690 537568
rect 654746 537512 654751 537568
rect 650164 537510 654751 537512
rect 654685 537507 654751 537510
rect 676262 535941 676322 536112
rect 676213 535936 676322 535941
rect 676213 535880 676218 535936
rect 676274 535880 676322 535936
rect 676213 535878 676322 535880
rect 676213 535875 676279 535878
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 679022 535125 679082 535296
rect 678973 535120 679082 535125
rect 678973 535064 678978 535120
rect 679034 535064 679082 535120
rect 678973 535062 679082 535064
rect 678973 535059 679039 535062
rect 676029 534918 676095 534921
rect 676029 534916 676292 534918
rect 676029 534860 676034 534916
rect 676090 534860 676292 534916
rect 676029 534858 676292 534860
rect 676029 534855 676095 534858
rect 676121 534306 676187 534309
rect 676262 534306 676322 534480
rect 679065 534306 679131 534309
rect 676121 534304 676322 534306
rect 676121 534248 676126 534304
rect 676182 534248 676322 534304
rect 676121 534246 676322 534248
rect 679022 534304 679131 534306
rect 679022 534248 679070 534304
rect 679126 534248 679131 534304
rect 676121 534243 676187 534246
rect 679022 534243 679131 534248
rect 679022 534072 679082 534243
rect 679022 533493 679082 533664
rect 679022 533488 679131 533493
rect 679022 533432 679070 533488
rect 679126 533432 679131 533488
rect 679022 533430 679131 533432
rect 679065 533427 679131 533430
rect 676029 533286 676095 533289
rect 676029 533284 676292 533286
rect 676029 533228 676034 533284
rect 676090 533228 676292 533284
rect 676029 533226 676292 533228
rect 676029 533223 676095 533226
rect 675937 532878 676003 532881
rect 675937 532876 676292 532878
rect 675937 532820 675942 532876
rect 675998 532820 676292 532876
rect 675937 532818 676292 532820
rect 675937 532815 676003 532818
rect 59261 532810 59327 532813
rect 59261 532808 64492 532810
rect 59261 532752 59266 532808
rect 59322 532752 64492 532808
rect 59261 532750 64492 532752
rect 59261 532747 59327 532750
rect 676213 532674 676279 532677
rect 676213 532672 676322 532674
rect 676213 532616 676218 532672
rect 676274 532616 676322 532672
rect 676213 532611 676322 532616
rect 676262 532440 676322 532611
rect 675753 532062 675819 532065
rect 675753 532060 676292 532062
rect 675753 532004 675758 532060
rect 675814 532004 676292 532060
rect 675753 532002 676292 532004
rect 675753 531999 675819 532002
rect 674598 531796 674604 531860
rect 674668 531858 674674 531860
rect 674668 531798 676322 531858
rect 674668 531796 674674 531798
rect 676262 531624 676322 531798
rect 676029 531246 676095 531249
rect 676029 531244 676292 531246
rect 676029 531188 676034 531244
rect 676090 531188 676292 531244
rect 676029 531186 676292 531188
rect 676029 531183 676095 531186
rect 675702 530776 675708 530840
rect 675772 530838 675778 530840
rect 675772 530778 676292 530838
rect 675772 530776 675778 530778
rect 674414 530572 674420 530636
rect 674484 530634 674490 530636
rect 674484 530574 676322 530634
rect 674484 530572 674490 530574
rect 676262 530400 676322 530574
rect 676029 530022 676095 530025
rect 676029 530020 676292 530022
rect 676029 529964 676034 530020
rect 676090 529964 676292 530020
rect 676029 529962 676292 529964
rect 676029 529959 676095 529962
rect 676029 529614 676095 529617
rect 676029 529612 676292 529614
rect 676029 529556 676034 529612
rect 676090 529556 676292 529612
rect 676029 529554 676292 529556
rect 676029 529551 676095 529554
rect 676070 529348 676076 529412
rect 676140 529410 676146 529412
rect 676140 529350 676322 529410
rect 676140 529348 676146 529350
rect 676262 529176 676322 529350
rect 675518 528940 675524 529004
rect 675588 529002 675594 529004
rect 675588 528942 676322 529002
rect 675588 528940 675594 528942
rect 676262 528768 676322 528942
rect 674230 528532 674236 528596
rect 674300 528594 674306 528596
rect 674300 528534 676322 528594
rect 674300 528532 674306 528534
rect 676262 528360 676322 528534
rect 676029 527982 676095 527985
rect 676029 527980 676292 527982
rect 676029 527924 676034 527980
rect 676090 527924 676292 527980
rect 676029 527922 676292 527924
rect 676029 527919 676095 527922
rect 676029 527574 676095 527577
rect 676029 527572 676292 527574
rect 676029 527516 676034 527572
rect 676090 527516 676292 527572
rect 676029 527514 676292 527516
rect 676029 527511 676095 527514
rect 676254 527308 676260 527372
rect 676324 527308 676330 527372
rect 676262 527136 676322 527308
rect 676806 526900 676812 526964
rect 676876 526900 676882 526964
rect 676814 526728 676874 526900
rect 676029 526350 676095 526353
rect 676029 526348 676292 526350
rect 676029 526292 676034 526348
rect 676090 526292 676292 526348
rect 676029 526290 676292 526292
rect 676029 526287 676095 526290
rect 679022 525741 679082 525912
rect 678973 525736 679082 525741
rect 678973 525680 678978 525736
rect 679034 525680 679082 525736
rect 678973 525678 679082 525680
rect 678973 525675 679039 525678
rect 684542 525333 684602 525504
rect 678973 525330 679039 525333
rect 678973 525328 679082 525330
rect 678973 525272 678978 525328
rect 679034 525272 679082 525328
rect 678973 525267 679082 525272
rect 684542 525328 684651 525333
rect 684542 525272 684590 525328
rect 684646 525272 684651 525328
rect 684542 525270 684651 525272
rect 684585 525267 684651 525270
rect 679022 525096 679082 525267
rect 684585 524922 684651 524925
rect 684542 524920 684651 524922
rect 684542 524864 684590 524920
rect 684646 524864 684651 524920
rect 684542 524859 684651 524864
rect 684542 524688 684602 524859
rect 654133 524242 654199 524245
rect 650164 524240 654199 524242
rect 650164 524184 654138 524240
rect 654194 524184 654199 524240
rect 650164 524182 654199 524184
rect 654133 524179 654199 524182
rect 58433 519754 58499 519757
rect 58433 519752 64492 519754
rect 58433 519696 58438 519752
rect 58494 519696 64492 519752
rect 58433 519694 64492 519696
rect 58433 519691 58499 519694
rect 654777 511050 654843 511053
rect 650164 511048 654843 511050
rect 650164 510992 654782 511048
rect 654838 510992 654843 511048
rect 650164 510990 654843 510992
rect 654777 510987 654843 510990
rect 58433 506698 58499 506701
rect 58433 506696 64492 506698
rect 58433 506640 58438 506696
rect 58494 506640 64492 506696
rect 58433 506638 64492 506640
rect 58433 506635 58499 506638
rect 656801 497722 656867 497725
rect 650164 497720 656867 497722
rect 650164 497664 656806 497720
rect 656862 497664 656867 497720
rect 650164 497662 656867 497664
rect 656801 497659 656867 497662
rect 57973 493642 58039 493645
rect 57973 493640 64492 493642
rect 57973 493584 57978 493640
rect 58034 493584 64492 493640
rect 57973 493582 64492 493584
rect 57973 493579 58039 493582
rect 676029 492146 676095 492149
rect 676029 492144 676292 492146
rect 676029 492088 676034 492144
rect 676090 492088 676292 492144
rect 676029 492086 676292 492088
rect 676029 492083 676095 492086
rect 675937 491738 676003 491741
rect 675937 491736 676292 491738
rect 675937 491680 675942 491736
rect 675998 491680 676292 491736
rect 675937 491678 676292 491680
rect 675937 491675 676003 491678
rect 676029 491330 676095 491333
rect 676029 491328 676292 491330
rect 676029 491272 676034 491328
rect 676090 491272 676292 491328
rect 676029 491270 676292 491272
rect 676029 491267 676095 491270
rect 675845 490922 675911 490925
rect 675845 490920 676292 490922
rect 675845 490864 675850 490920
rect 675906 490864 676292 490920
rect 675845 490862 676292 490864
rect 675845 490859 675911 490862
rect 675937 490514 676003 490517
rect 675937 490512 676292 490514
rect 675937 490456 675942 490512
rect 675998 490456 676292 490512
rect 675937 490454 676292 490456
rect 675937 490451 676003 490454
rect 676029 490106 676095 490109
rect 676029 490104 676292 490106
rect 676029 490048 676034 490104
rect 676090 490048 676292 490104
rect 676029 490046 676292 490048
rect 676029 490043 676095 490046
rect 675845 489698 675911 489701
rect 675845 489696 676292 489698
rect 675845 489640 675850 489696
rect 675906 489640 676292 489696
rect 675845 489638 676292 489640
rect 675845 489635 675911 489638
rect 673494 489228 673500 489292
rect 673564 489290 673570 489292
rect 676029 489290 676095 489293
rect 673564 489288 676292 489290
rect 673564 489232 676034 489288
rect 676090 489232 676292 489288
rect 673564 489230 676292 489232
rect 673564 489228 673570 489230
rect 676029 489227 676095 489230
rect 675661 488882 675727 488885
rect 675661 488880 676292 488882
rect 675661 488824 675666 488880
rect 675722 488824 676292 488880
rect 675661 488822 676292 488824
rect 675661 488819 675727 488822
rect 673862 488412 673868 488476
rect 673932 488474 673938 488476
rect 675753 488474 675819 488477
rect 673932 488472 676292 488474
rect 673932 488416 675758 488472
rect 675814 488416 676292 488472
rect 673932 488414 676292 488416
rect 673932 488412 673938 488414
rect 675753 488411 675819 488414
rect 675201 488066 675267 488069
rect 676029 488066 676095 488069
rect 675201 488064 676292 488066
rect 675201 488008 675206 488064
rect 675262 488008 676034 488064
rect 676090 488008 676292 488064
rect 675201 488006 676292 488008
rect 675201 488003 675267 488006
rect 676029 488003 676095 488006
rect 675150 487596 675156 487660
rect 675220 487658 675226 487660
rect 675220 487598 676292 487658
rect 675220 487596 675226 487598
rect 676029 487250 676095 487253
rect 676029 487248 676292 487250
rect 676029 487192 676034 487248
rect 676090 487192 676292 487248
rect 676029 487190 676292 487192
rect 676029 487187 676095 487190
rect 675334 486780 675340 486844
rect 675404 486842 675410 486844
rect 675404 486782 676292 486842
rect 675404 486780 675410 486782
rect 675937 486434 676003 486437
rect 675937 486432 676292 486434
rect 675937 486376 675942 486432
rect 675998 486376 676292 486432
rect 675937 486374 676292 486376
rect 675937 486371 676003 486374
rect 676029 486026 676095 486029
rect 676029 486024 676292 486026
rect 676029 485968 676034 486024
rect 676090 485968 676292 486024
rect 676029 485966 676292 485968
rect 676029 485963 676095 485966
rect 676029 485618 676095 485621
rect 676029 485616 676292 485618
rect 676029 485560 676034 485616
rect 676090 485560 676292 485616
rect 676029 485558 676292 485560
rect 676029 485555 676095 485558
rect 675886 485148 675892 485212
rect 675956 485210 675962 485212
rect 675956 485150 676292 485210
rect 675956 485148 675962 485150
rect 674966 484740 674972 484804
rect 675036 484802 675042 484804
rect 675036 484742 676292 484802
rect 675036 484740 675042 484742
rect 676070 484468 676076 484532
rect 676140 484468 676146 484532
rect 655053 484394 655119 484397
rect 650164 484392 655119 484394
rect 650164 484336 655058 484392
rect 655114 484336 655119 484392
rect 650164 484334 655119 484336
rect 676078 484394 676138 484468
rect 676078 484334 676292 484394
rect 655053 484331 655119 484334
rect 676029 483986 676095 483989
rect 676029 483984 676292 483986
rect 676029 483928 676034 483984
rect 676090 483928 676292 483984
rect 676029 483926 676292 483928
rect 676029 483923 676095 483926
rect 676029 483578 676095 483581
rect 676029 483576 676292 483578
rect 676029 483520 676034 483576
rect 676090 483520 676292 483576
rect 676029 483518 676292 483520
rect 676029 483515 676095 483518
rect 676070 483442 676076 483444
rect 676032 483380 676076 483442
rect 676140 483380 676146 483444
rect 676032 483306 676092 483380
rect 676032 483246 676230 483306
rect 676170 483170 676230 483246
rect 676170 483110 676292 483170
rect 675937 482762 676003 482765
rect 675937 482760 676292 482762
rect 675937 482704 675942 482760
rect 675998 482704 676292 482760
rect 675937 482702 676292 482704
rect 675937 482699 676003 482702
rect 676029 482354 676095 482357
rect 676029 482352 676292 482354
rect 676029 482296 676034 482352
rect 676090 482296 676292 482352
rect 676029 482294 676292 482296
rect 676029 482291 676095 482294
rect 676029 481946 676095 481949
rect 676029 481944 676292 481946
rect 676029 481888 676034 481944
rect 676090 481888 676292 481944
rect 676029 481886 676292 481888
rect 676029 481883 676095 481886
rect 675937 481538 676003 481541
rect 675937 481536 676292 481538
rect 675937 481480 675942 481536
rect 675998 481480 676292 481536
rect 675937 481478 676292 481480
rect 675937 481475 676003 481478
rect 676029 481130 676095 481133
rect 676029 481128 676292 481130
rect 676029 481072 676034 481128
rect 676090 481072 676292 481128
rect 676029 481070 676292 481072
rect 676029 481067 676095 481070
rect 675937 480722 676003 480725
rect 675937 480720 676292 480722
rect 675937 480664 675942 480720
rect 675998 480664 676292 480720
rect 675937 480662 676292 480664
rect 675937 480659 676003 480662
rect 58433 480586 58499 480589
rect 58433 480584 64492 480586
rect 58433 480528 58438 480584
rect 58494 480528 64492 480584
rect 58433 480526 64492 480528
rect 58433 480523 58499 480526
rect 654869 471202 654935 471205
rect 650164 471200 654935 471202
rect 650164 471144 654874 471200
rect 654930 471144 654935 471200
rect 650164 471142 654935 471144
rect 654869 471139 654935 471142
rect 58617 467530 58683 467533
rect 58617 467528 64492 467530
rect 58617 467472 58622 467528
rect 58678 467472 64492 467528
rect 58617 467470 64492 467472
rect 58617 467467 58683 467470
rect 654133 457874 654199 457877
rect 650164 457872 654199 457874
rect 650164 457816 654138 457872
rect 654194 457816 654199 457872
rect 650164 457814 654199 457816
rect 654133 457811 654199 457814
rect 59169 454610 59235 454613
rect 59169 454608 64492 454610
rect 59169 454552 59174 454608
rect 59230 454552 64492 454608
rect 59169 454550 64492 454552
rect 59169 454547 59235 454550
rect 656801 444546 656867 444549
rect 650164 444544 656867 444546
rect 650164 444488 656806 444544
rect 656862 444488 656867 444544
rect 650164 444486 656867 444488
rect 656801 444483 656867 444486
rect 58433 441554 58499 441557
rect 58433 441552 64492 441554
rect 58433 441496 58438 441552
rect 58494 441496 64492 441552
rect 58433 441494 64492 441496
rect 58433 441491 58499 441494
rect 654869 431354 654935 431357
rect 650164 431352 654935 431354
rect 650164 431296 654874 431352
rect 654930 431296 654935 431352
rect 650164 431294 654935 431296
rect 654869 431291 654935 431294
rect 41781 430946 41847 430949
rect 41492 430944 41847 430946
rect 41492 430888 41786 430944
rect 41842 430888 41847 430944
rect 41492 430886 41847 430888
rect 41781 430883 41847 430886
rect 51257 430538 51323 430541
rect 41492 430536 51323 430538
rect 41492 430480 51262 430536
rect 51318 430480 51323 430536
rect 41492 430478 51323 430480
rect 51257 430475 51323 430478
rect 53833 430130 53899 430133
rect 41492 430128 53899 430130
rect 41492 430072 53838 430128
rect 53894 430072 53899 430128
rect 41492 430070 53899 430072
rect 53833 430067 53899 430070
rect 43529 429722 43595 429725
rect 41492 429720 43595 429722
rect 41492 429664 43534 429720
rect 43590 429664 43595 429720
rect 41492 429662 43595 429664
rect 43529 429659 43595 429662
rect 43989 429314 44055 429317
rect 41492 429312 44055 429314
rect 41492 429256 43994 429312
rect 44050 429256 44055 429312
rect 41492 429254 44055 429256
rect 43989 429251 44055 429254
rect 43846 428906 43852 428908
rect 41492 428846 43852 428906
rect 43846 428844 43852 428846
rect 43916 428844 43922 428908
rect 43713 428498 43779 428501
rect 41492 428496 43779 428498
rect 41492 428440 43718 428496
rect 43774 428440 43779 428496
rect 41492 428438 43779 428440
rect 43713 428435 43779 428438
rect 57973 428498 58039 428501
rect 57973 428496 64492 428498
rect 57973 428440 57978 428496
rect 58034 428440 64492 428496
rect 57973 428438 64492 428440
rect 57973 428435 58039 428438
rect 39990 427854 40050 428060
rect 41822 427954 41828 427956
rect 41700 427894 41828 427954
rect 41784 427892 41828 427894
rect 41892 427954 41898 427956
rect 62757 427954 62823 427957
rect 41892 427952 62823 427954
rect 41892 427896 62762 427952
rect 62818 427896 62823 427952
rect 41892 427894 62823 427896
rect 41892 427892 41898 427894
rect 39982 427790 39988 427854
rect 40052 427790 40058 427854
rect 41784 427682 41844 427892
rect 62757 427891 62823 427894
rect 41492 427622 41844 427682
rect 41822 427274 41828 427276
rect 41492 427214 41828 427274
rect 41822 427212 41828 427214
rect 41892 427212 41898 427276
rect 41781 426866 41847 426869
rect 41492 426864 41847 426866
rect 41492 426808 41786 426864
rect 41842 426808 41847 426864
rect 41492 426806 41847 426808
rect 41781 426803 41847 426806
rect 43253 426458 43319 426461
rect 41492 426456 43319 426458
rect 41492 426400 43258 426456
rect 43314 426400 43319 426456
rect 41492 426398 43319 426400
rect 43253 426395 43319 426398
rect 42793 426050 42859 426053
rect 41492 426048 42859 426050
rect 41492 425992 42798 426048
rect 42854 425992 42859 426048
rect 41492 425990 42859 425992
rect 42793 425987 42859 425990
rect 42885 425642 42951 425645
rect 41492 425640 42951 425642
rect 41492 425584 42890 425640
rect 42946 425584 42951 425640
rect 41492 425582 42951 425584
rect 42885 425579 42951 425582
rect 43161 425234 43227 425237
rect 41492 425232 43227 425234
rect 41492 425176 43166 425232
rect 43222 425176 43227 425232
rect 41492 425174 43227 425176
rect 43161 425171 43227 425174
rect 43437 424826 43503 424829
rect 41492 424824 43503 424826
rect 41492 424768 43442 424824
rect 43498 424768 43503 424824
rect 41492 424766 43503 424768
rect 43437 424763 43503 424766
rect 41873 424418 41939 424421
rect 41492 424416 41939 424418
rect 41492 424360 41878 424416
rect 41934 424360 41939 424416
rect 41492 424358 41939 424360
rect 41873 424355 41939 424358
rect 43897 424010 43963 424013
rect 41492 424008 43963 424010
rect 41492 423952 43902 424008
rect 43958 423952 43963 424008
rect 41492 423950 43963 423952
rect 43897 423947 43963 423950
rect 43805 423602 43871 423605
rect 41492 423600 43871 423602
rect 41492 423544 43810 423600
rect 43866 423544 43871 423600
rect 41492 423542 43871 423544
rect 43805 423539 43871 423542
rect 43621 423194 43687 423197
rect 41492 423192 43687 423194
rect 41492 423136 43626 423192
rect 43682 423136 43687 423192
rect 41492 423134 43687 423136
rect 43621 423131 43687 423134
rect 42977 422786 43043 422789
rect 41492 422784 43043 422786
rect 41492 422728 42982 422784
rect 43038 422728 43043 422784
rect 41492 422726 43043 422728
rect 42977 422723 43043 422726
rect 43345 422378 43411 422381
rect 41492 422376 43411 422378
rect 41492 422320 43350 422376
rect 43406 422320 43411 422376
rect 41492 422318 43411 422320
rect 43345 422315 43411 422318
rect 43989 421970 44055 421973
rect 41492 421968 44055 421970
rect 41492 421912 43994 421968
rect 44050 421912 44055 421968
rect 41492 421910 44055 421912
rect 43989 421907 44055 421910
rect 41781 421562 41847 421565
rect 41492 421560 41847 421562
rect 41492 421504 41786 421560
rect 41842 421504 41847 421560
rect 41492 421502 41847 421504
rect 41781 421499 41847 421502
rect 42517 421154 42583 421157
rect 41492 421152 42583 421154
rect 41492 421096 42522 421152
rect 42578 421096 42583 421152
rect 41492 421094 42583 421096
rect 42517 421091 42583 421094
rect 41492 420686 41844 420746
rect 22694 419492 22754 420308
rect 41784 419930 41844 420686
rect 46657 419930 46723 419933
rect 41492 419928 46723 419930
rect 41492 419872 46662 419928
rect 46718 419872 46723 419928
rect 41492 419870 46723 419872
rect 46657 419867 46723 419870
rect 655053 418026 655119 418029
rect 650164 418024 655119 418026
rect 650164 417968 655058 418024
rect 655114 417968 655119 418024
rect 650164 417966 655119 417968
rect 655053 417963 655119 417966
rect 58433 415442 58499 415445
rect 58433 415440 64492 415442
rect 58433 415384 58438 415440
rect 58494 415384 64492 415440
rect 58433 415382 64492 415384
rect 58433 415379 58499 415382
rect 43529 411498 43595 411501
rect 42934 411496 43595 411498
rect 42934 411440 43534 411496
rect 43590 411440 43595 411496
rect 42934 411438 43595 411440
rect 42793 411270 42859 411273
rect 42934 411270 42994 411438
rect 43529 411435 43595 411438
rect 42793 411268 42994 411270
rect 42793 411212 42798 411268
rect 42854 411212 42994 411268
rect 42793 411210 42994 411212
rect 42793 411207 42859 411210
rect 654869 404698 654935 404701
rect 650164 404696 654935 404698
rect 650164 404640 654874 404696
rect 654930 404640 654935 404696
rect 650164 404638 654935 404640
rect 654869 404635 654935 404638
rect 676262 403749 676322 403852
rect 676213 403744 676322 403749
rect 676213 403688 676218 403744
rect 676274 403688 676322 403744
rect 676213 403686 676322 403688
rect 676213 403683 676279 403686
rect 675937 403474 676003 403477
rect 675937 403472 676292 403474
rect 675937 403416 675942 403472
rect 675998 403416 676292 403472
rect 675937 403414 676292 403416
rect 675937 403411 676003 403414
rect 675937 403066 676003 403069
rect 675937 403064 676292 403066
rect 675937 403008 675942 403064
rect 675998 403008 676292 403064
rect 675937 403006 676292 403008
rect 675937 403003 676003 403006
rect 676121 402930 676187 402933
rect 676121 402928 676322 402930
rect 676121 402872 676126 402928
rect 676182 402872 676322 402928
rect 676121 402870 676322 402872
rect 676121 402867 676187 402870
rect 676262 402628 676322 402870
rect 58433 402386 58499 402389
rect 58433 402384 64492 402386
rect 58433 402328 58438 402384
rect 58494 402328 64492 402384
rect 58433 402326 64492 402328
rect 58433 402323 58499 402326
rect 676121 402114 676187 402117
rect 676262 402114 676322 402220
rect 676121 402112 676322 402114
rect 676121 402056 676126 402112
rect 676182 402056 676322 402112
rect 676121 402054 676322 402056
rect 676121 402051 676187 402054
rect 675845 401842 675911 401845
rect 675845 401840 676292 401842
rect 675845 401784 675850 401840
rect 675906 401784 676292 401840
rect 675845 401782 676292 401784
rect 675845 401779 675911 401782
rect 675661 401434 675727 401437
rect 675661 401432 676292 401434
rect 675661 401376 675666 401432
rect 675722 401376 676292 401432
rect 675661 401374 676292 401376
rect 675661 401371 675727 401374
rect 673862 400964 673868 401028
rect 673932 401026 673938 401028
rect 675569 401026 675635 401029
rect 673932 401024 676292 401026
rect 673932 400968 675574 401024
rect 675630 400968 676292 401024
rect 673932 400966 676292 400968
rect 673932 400964 673938 400966
rect 675569 400963 675635 400966
rect 675753 400618 675819 400621
rect 675753 400616 676292 400618
rect 675753 400560 675758 400616
rect 675814 400560 676292 400616
rect 675753 400558 676292 400560
rect 675753 400555 675819 400558
rect 676029 400210 676095 400213
rect 676029 400208 676292 400210
rect 676029 400152 676034 400208
rect 676090 400152 676292 400208
rect 676029 400150 676292 400152
rect 676029 400147 676095 400150
rect 676029 399802 676095 399805
rect 676029 399800 676292 399802
rect 676029 399744 676034 399800
rect 676090 399744 676292 399800
rect 676029 399742 676292 399744
rect 676029 399739 676095 399742
rect 676029 399394 676095 399397
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 676121 398850 676187 398853
rect 676262 398850 676322 398956
rect 676121 398848 676322 398850
rect 676121 398792 676126 398848
rect 676182 398792 676322 398848
rect 676121 398790 676322 398792
rect 676121 398787 676187 398790
rect 675845 398578 675911 398581
rect 675845 398576 676292 398578
rect 675845 398520 675850 398576
rect 675906 398520 676292 398576
rect 675845 398518 676292 398520
rect 675845 398515 675911 398518
rect 676029 398170 676095 398173
rect 676029 398168 676292 398170
rect 676029 398112 676034 398168
rect 676090 398112 676292 398168
rect 676029 398110 676292 398112
rect 676029 398107 676095 398110
rect 675937 397762 676003 397765
rect 675937 397760 676292 397762
rect 675937 397704 675942 397760
rect 675998 397704 676292 397760
rect 675937 397702 676292 397704
rect 675937 397699 676003 397702
rect 676029 397354 676095 397357
rect 676029 397352 676292 397354
rect 676029 397296 676034 397352
rect 676090 397296 676292 397352
rect 676029 397294 676292 397296
rect 676029 397291 676095 397294
rect 675293 396946 675359 396949
rect 675293 396944 676292 396946
rect 675293 396888 675298 396944
rect 675354 396888 676292 396944
rect 675293 396886 676292 396888
rect 675293 396883 675359 396886
rect 676029 396538 676095 396541
rect 676029 396536 676292 396538
rect 676029 396480 676034 396536
rect 676090 396480 676292 396536
rect 676029 396478 676292 396480
rect 676029 396475 676095 396478
rect 676121 395994 676187 395997
rect 676262 395994 676322 396100
rect 676121 395992 676322 395994
rect 676121 395936 676126 395992
rect 676182 395936 676322 395992
rect 676121 395934 676322 395936
rect 676121 395931 676187 395934
rect 675937 395722 676003 395725
rect 675937 395720 676292 395722
rect 675937 395664 675942 395720
rect 675998 395664 676292 395720
rect 675937 395662 676292 395664
rect 675937 395659 676003 395662
rect 675937 395314 676003 395317
rect 675937 395312 676292 395314
rect 675937 395256 675942 395312
rect 675998 395256 676292 395312
rect 675937 395254 676292 395256
rect 675937 395251 676003 395254
rect 676029 394906 676095 394909
rect 676029 394904 676292 394906
rect 676029 394848 676034 394904
rect 676090 394848 676292 394904
rect 676029 394846 676292 394848
rect 676029 394843 676095 394846
rect 676029 394498 676095 394501
rect 676029 394496 676292 394498
rect 676029 394440 676034 394496
rect 676090 394440 676292 394496
rect 676029 394438 676292 394440
rect 676029 394435 676095 394438
rect 676029 394090 676095 394093
rect 676029 394088 676292 394090
rect 676029 394032 676034 394088
rect 676090 394032 676292 394088
rect 676029 394030 676292 394032
rect 676029 394027 676095 394030
rect 679022 393549 679082 393652
rect 678973 393544 679082 393549
rect 678973 393488 678978 393544
rect 679034 393488 679082 393544
rect 678973 393486 679082 393488
rect 678973 393483 679039 393486
rect 684542 393141 684602 393244
rect 678973 393138 679039 393141
rect 678973 393136 679082 393138
rect 678973 393080 678978 393136
rect 679034 393080 679082 393136
rect 678973 393075 679082 393080
rect 684493 393136 684602 393141
rect 684493 393080 684498 393136
rect 684554 393080 684602 393136
rect 684493 393078 684602 393080
rect 684493 393075 684559 393078
rect 679022 392836 679082 393075
rect 684493 392730 684559 392733
rect 684493 392728 684602 392730
rect 684493 392672 684498 392728
rect 684554 392672 684602 392728
rect 684493 392667 684602 392672
rect 684542 392428 684602 392667
rect 654133 391506 654199 391509
rect 650164 391504 654199 391506
rect 650164 391448 654138 391504
rect 654194 391448 654199 391504
rect 650164 391446 654199 391448
rect 654133 391443 654199 391446
rect 57973 389330 58039 389333
rect 57973 389328 64492 389330
rect 57973 389272 57978 389328
rect 58034 389272 64492 389328
rect 57973 389270 64492 389272
rect 57973 389267 58039 389270
rect 41505 387970 41571 387973
rect 41462 387968 41571 387970
rect 41462 387912 41510 387968
rect 41566 387912 41571 387968
rect 41462 387907 41571 387912
rect 41462 387668 41522 387907
rect 41781 387290 41847 387293
rect 41492 387288 41847 387290
rect 41492 387232 41786 387288
rect 41842 387232 41847 387288
rect 41492 387230 41847 387232
rect 41781 387227 41847 387230
rect 41505 387154 41571 387157
rect 41462 387152 41571 387154
rect 41462 387096 41510 387152
rect 41566 387096 41571 387152
rect 41462 387091 41571 387096
rect 41462 386852 41522 387091
rect 41462 386338 41522 386444
rect 42926 386338 42932 386340
rect 41462 386278 42932 386338
rect 42926 386276 42932 386278
rect 42996 386338 43002 386340
rect 62113 386338 62179 386341
rect 42996 386336 62179 386338
rect 42996 386280 62118 386336
rect 62174 386280 62179 386336
rect 42996 386278 62179 386280
rect 42996 386276 43002 386278
rect 62113 386275 62179 386278
rect 42793 386066 42859 386069
rect 41492 386064 42859 386066
rect 41492 386008 42798 386064
rect 42854 386008 42859 386064
rect 41492 386006 42859 386008
rect 42793 386003 42859 386006
rect 43713 385658 43779 385661
rect 41492 385656 43779 385658
rect 41492 385600 43718 385656
rect 43774 385600 43779 385656
rect 41492 385598 43779 385600
rect 43713 385595 43779 385598
rect 43529 385250 43595 385253
rect 41492 385248 43595 385250
rect 41492 385192 43534 385248
rect 43590 385192 43595 385248
rect 41492 385190 43595 385192
rect 43529 385187 43595 385190
rect 40174 384708 40234 384812
rect 39982 384644 39988 384708
rect 40052 384644 40058 384708
rect 40166 384644 40172 384708
rect 40236 384644 40242 384708
rect 39990 384404 40050 384644
rect 42742 384026 42748 384028
rect 41492 383966 42748 384026
rect 42742 383964 42748 383966
rect 42812 383964 42818 384028
rect 40350 383828 40356 383892
rect 40420 383890 40426 383892
rect 63309 383890 63375 383893
rect 40420 383888 63375 383890
rect 40420 383832 63314 383888
rect 63370 383832 63375 383888
rect 40420 383830 63375 383832
rect 40420 383828 40426 383830
rect 41278 383588 41338 383830
rect 63309 383827 63375 383830
rect 42742 383420 42748 383484
rect 42812 383482 42818 383484
rect 62021 383482 62087 383485
rect 42812 383480 62087 383482
rect 42812 383424 62026 383480
rect 62082 383424 62087 383480
rect 42812 383422 62087 383424
rect 42812 383420 42818 383422
rect 62021 383419 62087 383422
rect 42977 383210 43043 383213
rect 41492 383208 43043 383210
rect 41492 383152 42982 383208
rect 43038 383152 43043 383208
rect 41492 383150 43043 383152
rect 42977 383147 43043 383150
rect 40166 383012 40172 383076
rect 40236 383074 40242 383076
rect 62205 383074 62271 383077
rect 40236 383072 62271 383074
rect 40236 383016 62210 383072
rect 62266 383016 62271 383072
rect 40236 383014 62271 383016
rect 40236 383012 40242 383014
rect 62205 383011 62271 383014
rect 42701 382802 42767 382805
rect 41492 382800 42767 382802
rect 41492 382744 42706 382800
rect 42762 382744 42767 382800
rect 41492 382742 42767 382744
rect 42701 382739 42767 382742
rect 41462 382260 41522 382364
rect 41454 382196 41460 382260
rect 41524 382196 41530 382260
rect 42885 381986 42951 381989
rect 41492 381984 42951 381986
rect 41492 381928 42890 381984
rect 42946 381928 42951 381984
rect 41492 381926 42951 381928
rect 42885 381923 42951 381926
rect 42793 381578 42859 381581
rect 41492 381576 42859 381578
rect 41492 381520 42798 381576
rect 42854 381520 42859 381576
rect 41492 381518 42859 381520
rect 42793 381515 42859 381518
rect 42333 381170 42399 381173
rect 41492 381168 42399 381170
rect 41492 381112 42338 381168
rect 42394 381112 42399 381168
rect 41492 381110 42399 381112
rect 42333 381107 42399 381110
rect 43621 380762 43687 380765
rect 41492 380760 43687 380762
rect 41492 380704 43626 380760
rect 43682 380704 43687 380760
rect 41492 380702 43687 380704
rect 43621 380699 43687 380702
rect 43713 380354 43779 380357
rect 41492 380352 43779 380354
rect 41492 380296 43718 380352
rect 43774 380296 43779 380352
rect 41492 380294 43779 380296
rect 43713 380291 43779 380294
rect 43805 379946 43871 379949
rect 41492 379944 43871 379946
rect 41492 379888 43810 379944
rect 43866 379888 43871 379944
rect 41492 379886 43871 379888
rect 43805 379883 43871 379886
rect 43069 379538 43135 379541
rect 41492 379536 43135 379538
rect 41492 379480 43074 379536
rect 43130 379480 43135 379536
rect 41492 379478 43135 379480
rect 43069 379475 43135 379478
rect 43253 379130 43319 379133
rect 41492 379128 43319 379130
rect 41492 379072 43258 379128
rect 43314 379072 43319 379128
rect 41492 379070 43319 379072
rect 43253 379067 43319 379070
rect 43437 378722 43503 378725
rect 41492 378720 43503 378722
rect 41492 378664 43442 378720
rect 43498 378664 43503 378720
rect 41492 378662 43503 378664
rect 43437 378659 43503 378662
rect 43161 378314 43227 378317
rect 41492 378312 43227 378314
rect 41492 378256 43166 378312
rect 43222 378256 43227 378312
rect 41492 378254 43227 378256
rect 43161 378251 43227 378254
rect 656801 378178 656867 378181
rect 650164 378176 656867 378178
rect 650164 378120 656806 378176
rect 656862 378120 656867 378176
rect 650164 378118 656867 378120
rect 656801 378115 656867 378118
rect 41462 377773 41522 377876
rect 41462 377768 41571 377773
rect 41462 377712 41510 377768
rect 41566 377712 41571 377768
rect 41462 377710 41571 377712
rect 41505 377707 41571 377710
rect 41462 377365 41522 377468
rect 41413 377360 41522 377365
rect 41413 377304 41418 377360
rect 41474 377304 41522 377360
rect 41413 377302 41522 377304
rect 41413 377299 41479 377302
rect 30422 376957 30482 377060
rect 30422 376952 30531 376957
rect 30422 376896 30470 376952
rect 30526 376896 30531 376952
rect 30422 376894 30531 376896
rect 30465 376891 30531 376894
rect 41462 376549 41522 376652
rect 30465 376546 30531 376549
rect 30422 376544 30531 376546
rect 30422 376488 30470 376544
rect 30526 376488 30531 376544
rect 30422 376483 30531 376488
rect 41413 376544 41522 376549
rect 41413 376488 41418 376544
rect 41474 376488 41522 376544
rect 41413 376486 41522 376488
rect 41413 376483 41479 376486
rect 30422 376244 30482 376483
rect 58433 376274 58499 376277
rect 58433 376272 64492 376274
rect 58433 376216 58438 376272
rect 58494 376216 64492 376272
rect 58433 376214 64492 376216
rect 58433 376211 58499 376214
rect 656801 364850 656867 364853
rect 650164 364848 656867 364850
rect 650164 364792 656806 364848
rect 656862 364792 656867 364848
rect 650164 364790 656867 364792
rect 656801 364787 656867 364790
rect 58433 363354 58499 363357
rect 58433 363352 64492 363354
rect 58433 363296 58438 363352
rect 58494 363296 64492 363352
rect 58433 363294 64492 363296
rect 58433 363291 58499 363294
rect 675845 358730 675911 358733
rect 675845 358728 676292 358730
rect 675845 358672 675850 358728
rect 675906 358672 676292 358728
rect 675845 358670 676292 358672
rect 675845 358667 675911 358670
rect 675937 358322 676003 358325
rect 675937 358320 676292 358322
rect 675937 358264 675942 358320
rect 675998 358264 676292 358320
rect 675937 358262 676292 358264
rect 675937 358259 676003 358262
rect 676029 357914 676095 357917
rect 676029 357912 676292 357914
rect 676029 357856 676034 357912
rect 676090 357856 676292 357912
rect 676029 357854 676292 357856
rect 676029 357851 676095 357854
rect 674046 357444 674052 357508
rect 674116 357506 674122 357508
rect 674741 357506 674807 357509
rect 674116 357504 676292 357506
rect 674116 357448 674746 357504
rect 674802 357448 676292 357504
rect 674116 357446 676292 357448
rect 674116 357444 674122 357446
rect 674741 357443 674807 357446
rect 675569 357098 675635 357101
rect 675569 357096 676292 357098
rect 675569 357040 675574 357096
rect 675630 357040 676292 357096
rect 675569 357038 676292 357040
rect 675569 357035 675635 357038
rect 675661 356690 675727 356693
rect 675661 356688 676292 356690
rect 675661 356632 675666 356688
rect 675722 356632 676292 356688
rect 675661 356630 676292 356632
rect 675661 356627 675727 356630
rect 676029 356282 676095 356285
rect 676029 356280 676292 356282
rect 676029 356224 676034 356280
rect 676090 356224 676292 356280
rect 676029 356222 676292 356224
rect 676029 356219 676095 356222
rect 674414 355812 674420 355876
rect 674484 355874 674490 355876
rect 675753 355874 675819 355877
rect 674484 355872 676292 355874
rect 674484 355816 675758 355872
rect 675814 355816 676292 355872
rect 674484 355814 676292 355816
rect 674484 355812 674490 355814
rect 675753 355811 675819 355814
rect 41454 355676 41460 355740
rect 41524 355738 41530 355740
rect 41781 355738 41847 355741
rect 41524 355736 41847 355738
rect 41524 355680 41786 355736
rect 41842 355680 41847 355736
rect 41524 355678 41847 355680
rect 41524 355676 41530 355678
rect 41781 355675 41847 355678
rect 676029 355466 676095 355469
rect 676029 355464 676292 355466
rect 676029 355408 676034 355464
rect 676090 355408 676292 355464
rect 676029 355406 676292 355408
rect 676029 355403 676095 355406
rect 674230 354996 674236 355060
rect 674300 355058 674306 355060
rect 675293 355058 675359 355061
rect 674300 355056 676292 355058
rect 674300 355000 675298 355056
rect 675354 355000 676292 355056
rect 674300 354998 676292 355000
rect 674300 354996 674306 354998
rect 675293 354995 675359 354998
rect 676029 354650 676095 354653
rect 676029 354648 676292 354650
rect 676029 354592 676034 354648
rect 676090 354592 676292 354648
rect 676029 354590 676292 354592
rect 676029 354587 676095 354590
rect 676029 354242 676095 354245
rect 676029 354240 676292 354242
rect 676029 354184 676034 354240
rect 676090 354184 676292 354240
rect 676029 354182 676292 354184
rect 676029 354179 676095 354182
rect 676078 353774 676292 353834
rect 676078 353700 676138 353774
rect 676070 353636 676076 353700
rect 676140 353636 676146 353700
rect 676029 353426 676095 353429
rect 676029 353424 676292 353426
rect 676029 353368 676034 353424
rect 676090 353368 676292 353424
rect 676029 353366 676292 353368
rect 676029 353363 676095 353366
rect 676029 353018 676095 353021
rect 676029 353016 676292 353018
rect 676029 352960 676034 353016
rect 676090 352960 676292 353016
rect 676029 352958 676292 352960
rect 676029 352955 676095 352958
rect 675937 352610 676003 352613
rect 675937 352608 676292 352610
rect 675937 352552 675942 352608
rect 675998 352552 676292 352608
rect 675937 352550 676292 352552
rect 675937 352547 676003 352550
rect 675886 352140 675892 352204
rect 675956 352202 675962 352204
rect 675956 352142 676292 352202
rect 675956 352140 675962 352142
rect 33041 351930 33107 351933
rect 42926 351930 42932 351932
rect 33041 351928 42932 351930
rect 33041 351872 33046 351928
rect 33102 351872 42932 351928
rect 33041 351870 42932 351872
rect 33041 351867 33107 351870
rect 42926 351868 42932 351870
rect 42996 351868 43002 351932
rect 675293 351794 675359 351797
rect 675293 351792 676292 351794
rect 675293 351736 675298 351792
rect 675354 351736 676292 351792
rect 675293 351734 676292 351736
rect 675293 351731 675359 351734
rect 654869 351658 654935 351661
rect 650164 351656 654935 351658
rect 650164 351600 654874 351656
rect 654930 351600 654935 351656
rect 650164 351598 654935 351600
rect 654869 351595 654935 351598
rect 676029 351386 676095 351389
rect 676029 351384 676292 351386
rect 676029 351328 676034 351384
rect 676090 351328 676292 351384
rect 676029 351326 676292 351328
rect 676029 351323 676095 351326
rect 675937 350978 676003 350981
rect 675937 350976 676292 350978
rect 675937 350920 675942 350976
rect 675998 350920 676292 350976
rect 675937 350918 676292 350920
rect 675937 350915 676003 350918
rect 675702 350508 675708 350572
rect 675772 350570 675778 350572
rect 675772 350510 676292 350570
rect 675772 350508 675778 350510
rect 58433 350298 58499 350301
rect 58433 350296 64492 350298
rect 58433 350240 58438 350296
rect 58494 350240 64492 350296
rect 58433 350238 64492 350240
rect 58433 350235 58499 350238
rect 676029 350162 676095 350165
rect 676029 350160 676292 350162
rect 676029 350104 676034 350160
rect 676090 350104 676292 350160
rect 676029 350102 676292 350104
rect 676029 350099 676095 350102
rect 676029 349754 676095 349757
rect 676029 349752 676292 349754
rect 676029 349696 676034 349752
rect 676090 349696 676292 349752
rect 676029 349694 676292 349696
rect 676029 349691 676095 349694
rect 675937 349346 676003 349349
rect 675937 349344 676292 349346
rect 675937 349288 675942 349344
rect 675998 349288 676292 349344
rect 675937 349286 676292 349288
rect 675937 349283 676003 349286
rect 675845 348938 675911 348941
rect 675845 348936 676292 348938
rect 675845 348880 675850 348936
rect 675906 348880 676292 348936
rect 675845 348878 676292 348880
rect 675845 348875 675911 348878
rect 675753 348530 675819 348533
rect 675753 348528 676292 348530
rect 675753 348472 675758 348528
rect 675814 348472 676292 348528
rect 675753 348470 676292 348472
rect 675753 348467 675819 348470
rect 675661 348122 675727 348125
rect 675661 348120 676292 348122
rect 675661 348064 675666 348120
rect 675722 348064 676292 348120
rect 675661 348062 676292 348064
rect 675661 348059 675727 348062
rect 675753 347714 675819 347717
rect 675753 347712 676292 347714
rect 675753 347656 675758 347712
rect 675814 347656 676292 347712
rect 675753 347654 676292 347656
rect 675753 347651 675819 347654
rect 675661 347306 675727 347309
rect 675661 347304 676292 347306
rect 675661 347248 675666 347304
rect 675722 347248 676292 347304
rect 675661 347246 676292 347248
rect 675661 347243 675727 347246
rect 41462 344317 41522 344556
rect 41462 344312 41571 344317
rect 41462 344256 41510 344312
rect 41566 344256 41571 344312
rect 41462 344254 41571 344256
rect 41505 344251 41571 344254
rect 41781 344178 41847 344181
rect 41492 344176 41847 344178
rect 41492 344120 41786 344176
rect 41842 344120 41847 344176
rect 41492 344118 41847 344120
rect 41781 344115 41847 344118
rect 41597 343906 41663 343909
rect 41462 343904 41663 343906
rect 41462 343848 41602 343904
rect 41658 343848 41663 343904
rect 41462 343846 41663 343848
rect 41462 343740 41522 343846
rect 41597 343843 41663 343846
rect 672993 343634 673059 343637
rect 673177 343634 673243 343637
rect 672993 343632 673243 343634
rect 672993 343576 672998 343632
rect 673054 343576 673182 343632
rect 673238 343576 673243 343632
rect 672993 343574 673243 343576
rect 672993 343571 673059 343574
rect 673177 343571 673243 343574
rect 41781 343362 41847 343365
rect 41492 343360 41847 343362
rect 41492 343304 41786 343360
rect 41842 343304 41847 343360
rect 41492 343302 41847 343304
rect 41781 343299 41847 343302
rect 33041 343090 33107 343093
rect 32998 343088 33107 343090
rect 32998 343032 33046 343088
rect 33102 343032 33107 343088
rect 32998 343027 33107 343032
rect 32998 342924 33058 343027
rect 41505 342682 41571 342685
rect 41462 342680 41571 342682
rect 41462 342624 41510 342680
rect 41566 342624 41571 342680
rect 41462 342619 41571 342624
rect 41462 342516 41522 342619
rect 43253 342138 43319 342141
rect 41492 342136 43319 342138
rect 41492 342080 43258 342136
rect 43314 342080 43319 342136
rect 41492 342078 43319 342080
rect 43253 342075 43319 342078
rect 44265 341730 44331 341733
rect 41492 341728 44331 341730
rect 41492 341672 44270 341728
rect 44326 341672 44331 341728
rect 41492 341670 44331 341672
rect 44265 341667 44331 341670
rect 40166 341396 40172 341460
rect 40236 341396 40242 341460
rect 40174 341292 40234 341396
rect 44173 340914 44239 340917
rect 46197 340914 46263 340917
rect 41492 340912 46263 340914
rect 41492 340856 44178 340912
rect 44234 340856 46202 340912
rect 46258 340856 46263 340912
rect 41492 340854 46263 340856
rect 44173 340851 44239 340854
rect 46197 340851 46263 340854
rect 42742 340506 42748 340508
rect 41492 340446 42748 340506
rect 42742 340444 42748 340446
rect 42812 340444 42818 340508
rect 44265 340098 44331 340101
rect 46381 340098 46447 340101
rect 44265 340096 46447 340098
rect 32673 339826 32739 339829
rect 32630 339824 32739 339826
rect 32630 339768 32678 339824
rect 32734 339768 32739 339824
rect 32630 339763 32739 339768
rect 41462 339826 41522 340068
rect 44265 340040 44270 340096
rect 44326 340040 46386 340096
rect 46442 340040 46447 340096
rect 44265 340038 46447 340040
rect 44265 340035 44331 340038
rect 46381 340035 46447 340038
rect 41462 339766 41890 339826
rect 32630 339660 32690 339763
rect 41830 339418 41890 339766
rect 42558 339418 42564 339420
rect 41830 339358 42564 339418
rect 42558 339356 42564 339358
rect 42628 339356 42634 339420
rect 41822 339282 41828 339284
rect 41492 339222 41828 339282
rect 41822 339220 41828 339222
rect 41892 339220 41898 339284
rect 32630 338605 32690 338844
rect 32581 338600 32690 338605
rect 32581 338544 32586 338600
rect 32642 338544 32690 338600
rect 32581 338542 32690 338544
rect 32581 338539 32647 338542
rect 32814 338197 32874 338436
rect 654317 338330 654383 338333
rect 650164 338328 654383 338330
rect 650164 338272 654322 338328
rect 654378 338272 654383 338328
rect 650164 338270 654383 338272
rect 654317 338267 654383 338270
rect 32765 338192 32874 338197
rect 32765 338136 32770 338192
rect 32826 338136 32874 338192
rect 32765 338134 32874 338136
rect 32765 338131 32831 338134
rect 32998 337789 33058 338028
rect 32998 337784 33107 337789
rect 32998 337728 33046 337784
rect 33102 337728 33107 337784
rect 32998 337726 33107 337728
rect 33041 337723 33107 337726
rect 41462 337378 41522 337620
rect 41638 337378 41644 337380
rect 41462 337318 41644 337378
rect 41638 337316 41644 337318
rect 41708 337316 41714 337380
rect 42190 337242 42196 337244
rect 41492 337182 42196 337242
rect 42190 337180 42196 337182
rect 42260 337180 42266 337244
rect 58433 337242 58499 337245
rect 58433 337240 64492 337242
rect 58433 337184 58438 337240
rect 58494 337184 64492 337240
rect 58433 337182 64492 337184
rect 58433 337179 58499 337182
rect 42006 336834 42012 336836
rect 41492 336774 42012 336834
rect 42006 336772 42012 336774
rect 42076 336772 42082 336836
rect 32998 336157 33058 336396
rect 32949 336152 33058 336157
rect 32949 336096 32954 336152
rect 33010 336096 33058 336152
rect 32949 336094 33058 336096
rect 32949 336091 33015 336094
rect 32814 335749 32874 335988
rect 32814 335744 32923 335749
rect 32814 335688 32862 335744
rect 32918 335688 32923 335744
rect 32814 335686 32923 335688
rect 32857 335683 32923 335686
rect 43069 335610 43135 335613
rect 41492 335608 43135 335610
rect 41492 335552 43074 335608
rect 43130 335552 43135 335608
rect 41492 335550 43135 335552
rect 43069 335547 43135 335550
rect 42977 335202 43043 335205
rect 41492 335200 43043 335202
rect 41492 335144 42982 335200
rect 43038 335144 43043 335200
rect 41492 335142 43043 335144
rect 42977 335139 43043 335142
rect 43161 334794 43227 334797
rect 41492 334792 43227 334794
rect 41492 334736 43166 334792
rect 43222 334736 43227 334792
rect 41492 334734 43227 334736
rect 43161 334731 43227 334734
rect 41462 334117 41522 334356
rect 41462 334112 41571 334117
rect 41462 334056 41510 334112
rect 41566 334056 41571 334112
rect 41462 334054 41571 334056
rect 41505 334051 41571 334054
rect 30422 333709 30482 333948
rect 30373 333704 30482 333709
rect 30373 333648 30378 333704
rect 30434 333648 30482 333704
rect 30373 333646 30482 333648
rect 30373 333643 30439 333646
rect 41462 333301 41522 333540
rect 30373 333298 30439 333301
rect 30373 333296 30482 333298
rect 30373 333240 30378 333296
rect 30434 333240 30482 333296
rect 30373 333235 30482 333240
rect 41462 333296 41571 333301
rect 41462 333240 41510 333296
rect 41566 333240 41571 333296
rect 41462 333238 41571 333240
rect 41505 333235 41571 333238
rect 30422 333132 30482 333235
rect 675661 330580 675727 330581
rect 675661 330576 675708 330580
rect 675772 330578 675778 330580
rect 675661 330520 675666 330576
rect 675661 330516 675708 330520
rect 675772 330518 675818 330578
rect 675772 330516 675778 330518
rect 675661 330515 675727 330516
rect 32765 329898 32831 329901
rect 41454 329898 41460 329900
rect 32765 329896 41460 329898
rect 32765 329840 32770 329896
rect 32826 329840 41460 329896
rect 32765 329838 41460 329840
rect 32765 329835 32831 329838
rect 41454 329836 41460 329838
rect 41524 329836 41530 329900
rect 32581 329762 32647 329765
rect 42374 329762 42380 329764
rect 32581 329760 42380 329762
rect 32581 329704 32586 329760
rect 32642 329704 42380 329760
rect 32581 329702 42380 329704
rect 32581 329699 32647 329702
rect 42374 329700 42380 329702
rect 42444 329700 42450 329764
rect 675753 328402 675819 328405
rect 676070 328402 676076 328404
rect 675753 328400 676076 328402
rect 675753 328344 675758 328400
rect 675814 328344 676076 328400
rect 675753 328342 676076 328344
rect 675753 328339 675819 328342
rect 676070 328340 676076 328342
rect 676140 328340 676146 328404
rect 675753 326906 675819 326909
rect 675886 326906 675892 326908
rect 675753 326904 675892 326906
rect 675753 326848 675758 326904
rect 675814 326848 675892 326904
rect 675753 326846 675892 326848
rect 675753 326843 675819 326846
rect 675886 326844 675892 326846
rect 675956 326844 675962 326908
rect 654317 325002 654383 325005
rect 650164 325000 654383 325002
rect 650164 324944 654322 325000
rect 654378 324944 654383 325000
rect 650164 324942 654383 324944
rect 654317 324939 654383 324942
rect 58157 324186 58223 324189
rect 58157 324184 64492 324186
rect 58157 324128 58162 324184
rect 58218 324128 64492 324184
rect 58157 324126 64492 324128
rect 58157 324123 58223 324126
rect 41454 319908 41460 319972
rect 41524 319970 41530 319972
rect 41781 319970 41847 319973
rect 41524 319968 41847 319970
rect 41524 319912 41786 319968
rect 41842 319912 41847 319968
rect 41524 319910 41847 319912
rect 41524 319908 41530 319910
rect 41781 319907 41847 319910
rect 41965 316980 42031 316981
rect 41965 316976 42012 316980
rect 42076 316978 42082 316980
rect 41965 316920 41970 316976
rect 41965 316916 42012 316920
rect 42076 316918 42122 316978
rect 42076 316916 42082 316918
rect 41965 316915 42031 316916
rect 40350 316100 40356 316164
rect 40420 316162 40426 316164
rect 62021 316162 62087 316165
rect 40420 316160 62087 316162
rect 40420 316104 62026 316160
rect 62082 316104 62087 316160
rect 40420 316102 62087 316104
rect 40420 316100 40426 316102
rect 62021 316099 62087 316102
rect 42149 316028 42215 316029
rect 42149 316026 42196 316028
rect 42104 316024 42196 316026
rect 42104 315968 42154 316024
rect 42104 315966 42196 315968
rect 42149 315964 42196 315966
rect 42260 315964 42266 316028
rect 42149 315963 42215 315964
rect 42149 315482 42215 315485
rect 42374 315482 42380 315484
rect 42149 315480 42380 315482
rect 42149 315424 42154 315480
rect 42210 315424 42380 315480
rect 42149 315422 42380 315424
rect 42149 315419 42215 315422
rect 42374 315420 42380 315422
rect 42444 315420 42450 315484
rect 42149 313850 42215 313853
rect 42558 313850 42564 313852
rect 42149 313848 42564 313850
rect 42149 313792 42154 313848
rect 42210 313792 42564 313848
rect 42149 313790 42564 313792
rect 42149 313787 42215 313790
rect 42558 313788 42564 313790
rect 42628 313788 42634 313852
rect 676262 313581 676322 313684
rect 676213 313576 676322 313581
rect 676213 313520 676218 313576
rect 676274 313520 676322 313576
rect 676213 313518 676322 313520
rect 676213 313515 676279 313518
rect 676029 313306 676095 313309
rect 676029 313304 676292 313306
rect 676029 313248 676034 313304
rect 676090 313248 676292 313304
rect 676029 313246 676292 313248
rect 676029 313243 676095 313246
rect 41638 313108 41644 313172
rect 41708 313170 41714 313172
rect 41781 313170 41847 313173
rect 41708 313168 41847 313170
rect 41708 313112 41786 313168
rect 41842 313112 41847 313168
rect 41708 313110 41847 313112
rect 41708 313108 41714 313110
rect 41781 313107 41847 313110
rect 676029 312898 676095 312901
rect 676029 312896 676292 312898
rect 676029 312840 676034 312896
rect 676090 312840 676292 312896
rect 676029 312838 676292 312840
rect 676029 312835 676095 312838
rect 676029 312490 676095 312493
rect 676029 312488 676292 312490
rect 676029 312432 676034 312488
rect 676090 312432 676292 312488
rect 676029 312430 676292 312432
rect 676029 312427 676095 312430
rect 41781 312356 41847 312357
rect 41781 312352 41828 312356
rect 41892 312354 41898 312356
rect 41781 312296 41786 312352
rect 41781 312292 41828 312296
rect 41892 312294 41938 312354
rect 41892 312292 41898 312294
rect 41781 312291 41847 312292
rect 676029 312082 676095 312085
rect 676029 312080 676292 312082
rect 676029 312024 676034 312080
rect 676090 312024 676292 312080
rect 676029 312022 676292 312024
rect 676029 312019 676095 312022
rect 654133 311810 654199 311813
rect 650164 311808 654199 311810
rect 650164 311752 654138 311808
rect 654194 311752 654199 311808
rect 650164 311750 654199 311752
rect 654133 311747 654199 311750
rect 676029 311674 676095 311677
rect 676029 311672 676292 311674
rect 676029 311616 676034 311672
rect 676090 311616 676292 311672
rect 676029 311614 676292 311616
rect 676029 311611 676095 311614
rect 676029 311266 676095 311269
rect 676029 311264 676292 311266
rect 676029 311208 676034 311264
rect 676090 311208 676292 311264
rect 676029 311206 676292 311208
rect 676029 311203 676095 311206
rect 59261 311130 59327 311133
rect 59261 311128 64492 311130
rect 59261 311072 59266 311128
rect 59322 311072 64492 311128
rect 59261 311070 64492 311072
rect 59261 311067 59327 311070
rect 676029 310858 676095 310861
rect 676029 310856 676292 310858
rect 676029 310800 676034 310856
rect 676090 310800 676292 310856
rect 676029 310798 676292 310800
rect 676029 310795 676095 310798
rect 676029 310450 676095 310453
rect 676029 310448 676292 310450
rect 676029 310392 676034 310448
rect 676090 310392 676292 310448
rect 676029 310390 676292 310392
rect 676029 310387 676095 310390
rect 676029 310042 676095 310045
rect 676029 310040 676292 310042
rect 676029 309984 676034 310040
rect 676090 309984 676292 310040
rect 676029 309982 676292 309984
rect 676029 309979 676095 309982
rect 676029 309634 676095 309637
rect 676029 309632 676292 309634
rect 676029 309576 676034 309632
rect 676090 309576 676292 309632
rect 676029 309574 676292 309576
rect 676029 309571 676095 309574
rect 676029 309226 676095 309229
rect 676029 309224 676292 309226
rect 676029 309168 676034 309224
rect 676090 309168 676292 309224
rect 676029 309166 676292 309168
rect 676029 309163 676095 309166
rect 676029 308818 676095 308821
rect 676029 308816 676292 308818
rect 676029 308760 676034 308816
rect 676090 308760 676292 308816
rect 676029 308758 676292 308760
rect 676029 308755 676095 308758
rect 675753 308410 675819 308413
rect 675753 308408 676292 308410
rect 675753 308352 675758 308408
rect 675814 308352 676292 308408
rect 675753 308350 676292 308352
rect 675753 308347 675819 308350
rect 676029 308002 676095 308005
rect 676029 308000 676292 308002
rect 676029 307944 676034 308000
rect 676090 307944 676292 308000
rect 676029 307942 676292 307944
rect 676029 307939 676095 307942
rect 676121 307458 676187 307461
rect 676262 307458 676322 307564
rect 676121 307456 676322 307458
rect 676121 307400 676126 307456
rect 676182 307400 676322 307456
rect 676121 307398 676322 307400
rect 676121 307395 676187 307398
rect 675937 307186 676003 307189
rect 675937 307184 676292 307186
rect 675937 307128 675942 307184
rect 675998 307128 676292 307184
rect 675937 307126 676292 307128
rect 675937 307123 676003 307126
rect 676029 306778 676095 306781
rect 676029 306776 676292 306778
rect 676029 306720 676034 306776
rect 676090 306720 676292 306776
rect 676029 306718 676292 306720
rect 676029 306715 676095 306718
rect 675886 306308 675892 306372
rect 675956 306370 675962 306372
rect 675956 306310 676292 306370
rect 675956 306308 675962 306310
rect 676029 305962 676095 305965
rect 676029 305960 676292 305962
rect 676029 305904 676034 305960
rect 676090 305904 676292 305960
rect 676029 305902 676292 305904
rect 676029 305899 676095 305902
rect 676121 305418 676187 305421
rect 676262 305418 676322 305524
rect 676121 305416 676322 305418
rect 676121 305360 676126 305416
rect 676182 305360 676322 305416
rect 676121 305358 676322 305360
rect 676121 305355 676187 305358
rect 676121 305010 676187 305013
rect 676262 305010 676322 305116
rect 676121 305008 676322 305010
rect 676121 304952 676126 305008
rect 676182 304952 676322 305008
rect 676121 304950 676322 304952
rect 676121 304947 676187 304950
rect 676029 304738 676095 304741
rect 676029 304736 676292 304738
rect 676029 304680 676034 304736
rect 676090 304680 676292 304736
rect 676029 304678 676292 304680
rect 676029 304675 676095 304678
rect 676121 304194 676187 304197
rect 676262 304194 676322 304300
rect 676121 304192 676322 304194
rect 676121 304136 676126 304192
rect 676182 304136 676322 304192
rect 676121 304134 676322 304136
rect 676121 304131 676187 304134
rect 675937 303922 676003 303925
rect 675937 303920 676292 303922
rect 675937 303864 675942 303920
rect 675998 303864 676292 303920
rect 675937 303862 676292 303864
rect 675937 303859 676003 303862
rect 679022 303381 679082 303484
rect 679022 303376 679131 303381
rect 679022 303320 679070 303376
rect 679126 303320 679131 303376
rect 679022 303318 679131 303320
rect 679065 303315 679131 303318
rect 684542 302973 684602 303076
rect 679065 302970 679131 302973
rect 679022 302968 679131 302970
rect 679022 302912 679070 302968
rect 679126 302912 679131 302968
rect 679022 302907 679131 302912
rect 684493 302968 684602 302973
rect 684493 302912 684498 302968
rect 684554 302912 684602 302968
rect 684493 302910 684602 302912
rect 684493 302907 684559 302910
rect 679022 302668 679082 302907
rect 684493 302562 684559 302565
rect 684493 302560 684602 302562
rect 684493 302504 684498 302560
rect 684554 302504 684602 302560
rect 684493 302499 684602 302504
rect 684542 302260 684602 302499
rect 41505 301610 41571 301613
rect 41462 301608 41571 301610
rect 41462 301552 41510 301608
rect 41566 301552 41571 301608
rect 41462 301547 41571 301552
rect 41462 301308 41522 301547
rect 41781 300930 41847 300933
rect 41492 300928 41847 300930
rect 41492 300872 41786 300928
rect 41842 300872 41847 300928
rect 41492 300870 41847 300872
rect 41781 300867 41847 300870
rect 53833 300522 53899 300525
rect 41492 300520 53899 300522
rect 41492 300464 53838 300520
rect 53894 300464 53899 300520
rect 41492 300462 53899 300464
rect 53833 300459 53899 300462
rect 41822 300114 41828 300116
rect 41492 300054 41828 300114
rect 41822 300052 41828 300054
rect 41892 300114 41898 300116
rect 48313 300114 48379 300117
rect 41892 300112 48379 300114
rect 41892 300056 48318 300112
rect 48374 300056 48379 300112
rect 41892 300054 48379 300056
rect 41892 300052 41898 300054
rect 48313 300051 48379 300054
rect 44357 299706 44423 299709
rect 41492 299704 44423 299706
rect 41492 299648 44362 299704
rect 44418 299648 44423 299704
rect 41492 299646 44423 299648
rect 44357 299643 44423 299646
rect 43253 299298 43319 299301
rect 41492 299296 43319 299298
rect 41492 299240 43258 299296
rect 43314 299240 43319 299296
rect 41492 299238 43319 299240
rect 43253 299235 43319 299238
rect 43529 298890 43595 298893
rect 41492 298888 43595 298890
rect 41492 298832 43534 298888
rect 43590 298832 43595 298888
rect 41492 298830 43595 298832
rect 43529 298827 43595 298830
rect 41822 298482 41828 298484
rect 41492 298422 41828 298482
rect 41822 298420 41828 298422
rect 41892 298482 41898 298484
rect 46105 298482 46171 298485
rect 656801 298482 656867 298485
rect 41892 298480 46171 298482
rect 41892 298424 46110 298480
rect 46166 298424 46171 298480
rect 41892 298422 46171 298424
rect 650164 298480 656867 298482
rect 650164 298424 656806 298480
rect 656862 298424 656867 298480
rect 650164 298422 656867 298424
rect 41892 298420 41898 298422
rect 46105 298419 46171 298422
rect 656801 298419 656867 298422
rect 59353 298210 59419 298213
rect 59353 298208 64492 298210
rect 59353 298152 59358 298208
rect 59414 298152 64492 298208
rect 59353 298150 64492 298152
rect 59353 298147 59419 298150
rect 44265 298074 44331 298077
rect 41492 298072 44331 298074
rect 41492 298016 44270 298072
rect 44326 298016 44331 298072
rect 41492 298014 44331 298016
rect 44265 298011 44331 298014
rect 42006 297666 42012 297668
rect 41492 297606 42012 297666
rect 42006 297604 42012 297606
rect 42076 297666 42082 297668
rect 48221 297666 48287 297669
rect 42076 297664 48287 297666
rect 42076 297608 48226 297664
rect 48282 297608 48287 297664
rect 42076 297606 48287 297608
rect 42076 297604 42082 297606
rect 48221 297603 48287 297606
rect 44173 297258 44239 297261
rect 41492 297256 44239 297258
rect 41492 297200 44178 297256
rect 44234 297200 44239 297256
rect 41492 297198 44239 297200
rect 44173 297195 44239 297198
rect 32765 296850 32831 296853
rect 32765 296848 32844 296850
rect 32765 296792 32770 296848
rect 32826 296792 32844 296848
rect 32765 296790 32844 296792
rect 32765 296787 32831 296790
rect 35801 296442 35867 296445
rect 35788 296440 35867 296442
rect 35788 296384 35806 296440
rect 35862 296384 35867 296440
rect 35788 296382 35867 296384
rect 35801 296379 35867 296382
rect 32581 296034 32647 296037
rect 32581 296032 32660 296034
rect 32581 295976 32586 296032
rect 32642 295976 32660 296032
rect 32581 295974 32660 295976
rect 32581 295971 32647 295974
rect 41492 295566 41890 295626
rect 32857 295218 32923 295221
rect 32844 295216 32923 295218
rect 32844 295160 32862 295216
rect 32918 295160 32923 295216
rect 32844 295158 32923 295160
rect 41830 295218 41890 295566
rect 42006 295218 42012 295220
rect 41830 295158 42012 295218
rect 32857 295155 32923 295158
rect 42006 295156 42012 295158
rect 42076 295156 42082 295220
rect 32673 294810 32739 294813
rect 32660 294808 32739 294810
rect 32660 294752 32678 294808
rect 32734 294752 32739 294808
rect 32660 294750 32739 294752
rect 32673 294747 32739 294750
rect 33041 294402 33107 294405
rect 33028 294400 33107 294402
rect 33028 294344 33046 294400
rect 33102 294344 33107 294400
rect 33028 294342 33107 294344
rect 33041 294339 33107 294342
rect 32949 293994 33015 293997
rect 32949 293992 33028 293994
rect 32949 293936 32954 293992
rect 33010 293936 33028 293992
rect 32949 293934 33028 293936
rect 32949 293931 33015 293934
rect 42885 293586 42951 293589
rect 41492 293584 42951 293586
rect 41492 293528 42890 293584
rect 42946 293528 42951 293584
rect 41492 293526 42951 293528
rect 42885 293523 42951 293526
rect 42977 293178 43043 293181
rect 41492 293176 43043 293178
rect 41492 293120 42982 293176
rect 43038 293120 43043 293176
rect 41492 293118 43043 293120
rect 42977 293115 43043 293118
rect 43161 292770 43227 292773
rect 41492 292768 43227 292770
rect 41492 292712 43166 292768
rect 43222 292712 43227 292768
rect 41492 292710 43227 292712
rect 43161 292707 43227 292710
rect 43069 292362 43135 292365
rect 41492 292360 43135 292362
rect 41492 292304 43074 292360
rect 43130 292304 43135 292360
rect 41492 292302 43135 292304
rect 43069 292299 43135 292302
rect 675753 292226 675819 292229
rect 675886 292226 675892 292228
rect 675753 292224 675892 292226
rect 675753 292168 675758 292224
rect 675814 292168 675892 292224
rect 675753 292166 675892 292168
rect 675753 292163 675819 292166
rect 675886 292164 675892 292166
rect 675956 292164 675962 292228
rect 43621 291954 43687 291957
rect 41492 291952 43687 291954
rect 41492 291896 43626 291952
rect 43682 291896 43687 291952
rect 41492 291894 43687 291896
rect 43621 291891 43687 291894
rect 43345 291546 43411 291549
rect 41492 291544 43411 291546
rect 41492 291488 43350 291544
rect 43406 291488 43411 291544
rect 41492 291486 43411 291488
rect 43345 291483 43411 291486
rect 46105 291138 46171 291141
rect 41492 291136 46171 291138
rect 41492 291080 46110 291136
rect 46166 291080 46171 291136
rect 41492 291078 46171 291080
rect 46105 291075 46171 291078
rect 46381 290730 46447 290733
rect 41492 290728 46447 290730
rect 41492 290672 46386 290728
rect 46442 290672 46447 290728
rect 41492 290670 46447 290672
rect 46381 290667 46447 290670
rect 46841 290322 46907 290325
rect 41492 290320 46907 290322
rect 41492 290264 46846 290320
rect 46902 290264 46907 290320
rect 41492 290262 46907 290264
rect 46841 290259 46907 290262
rect 33041 285970 33107 285973
rect 42190 285970 42196 285972
rect 33041 285968 42196 285970
rect 33041 285912 33046 285968
rect 33102 285912 42196 285968
rect 33041 285910 42196 285912
rect 33041 285907 33107 285910
rect 42190 285908 42196 285910
rect 42260 285908 42266 285972
rect 32765 285834 32831 285837
rect 42374 285834 42380 285836
rect 32765 285832 42380 285834
rect 32765 285776 32770 285832
rect 32826 285776 42380 285832
rect 32765 285774 42380 285776
rect 32765 285771 32831 285774
rect 42374 285772 42380 285774
rect 42444 285772 42450 285836
rect 32581 285698 32647 285701
rect 42558 285698 42564 285700
rect 32581 285696 42564 285698
rect 32581 285640 32586 285696
rect 32642 285640 42564 285696
rect 32581 285638 42564 285640
rect 32581 285635 32647 285638
rect 42558 285636 42564 285638
rect 42628 285636 42634 285700
rect 655697 285290 655763 285293
rect 650164 285288 655763 285290
rect 650164 285232 655702 285288
rect 655758 285232 655763 285288
rect 650164 285230 655763 285232
rect 655697 285227 655763 285230
rect 59445 285154 59511 285157
rect 59445 285152 64492 285154
rect 59445 285096 59450 285152
rect 59506 285096 64492 285152
rect 59445 285094 64492 285096
rect 59445 285091 59511 285094
rect 44030 278428 44036 278492
rect 44100 278490 44106 278492
rect 672809 278490 672875 278493
rect 44100 278488 672875 278490
rect 44100 278432 672814 278488
rect 672870 278432 672875 278488
rect 44100 278430 672875 278432
rect 44100 278428 44106 278430
rect 672809 278427 672875 278430
rect 62297 278354 62363 278357
rect 674414 278354 674420 278356
rect 62297 278352 674420 278354
rect 62297 278296 62302 278352
rect 62358 278296 674420 278352
rect 62297 278294 674420 278296
rect 62297 278291 62363 278294
rect 674414 278292 674420 278294
rect 674484 278292 674490 278356
rect 62481 278218 62547 278221
rect 674046 278218 674052 278220
rect 62481 278216 674052 278218
rect 62481 278160 62486 278216
rect 62542 278160 674052 278216
rect 62481 278158 674052 278160
rect 62481 278155 62547 278158
rect 674046 278156 674052 278158
rect 674116 278156 674122 278220
rect 62665 278082 62731 278085
rect 674230 278082 674236 278084
rect 62665 278080 674236 278082
rect 62665 278024 62670 278080
rect 62726 278024 674236 278080
rect 62665 278022 674236 278024
rect 62665 278019 62731 278022
rect 674230 278020 674236 278022
rect 674300 278020 674306 278084
rect 62849 277946 62915 277949
rect 673862 277946 673868 277948
rect 62849 277944 673868 277946
rect 62849 277888 62854 277944
rect 62910 277888 673868 277944
rect 62849 277886 673868 277888
rect 62849 277883 62915 277886
rect 673862 277884 673868 277886
rect 673932 277884 673938 277948
rect 63033 277810 63099 277813
rect 673678 277810 673684 277812
rect 63033 277808 673684 277810
rect 63033 277752 63038 277808
rect 63094 277752 673684 277808
rect 63033 277750 673684 277752
rect 63033 277747 63099 277750
rect 673678 277748 673684 277750
rect 673748 277748 673754 277812
rect 63217 277674 63283 277677
rect 673494 277674 673500 277676
rect 63217 277672 673500 277674
rect 63217 277616 63222 277672
rect 63278 277616 673500 277672
rect 63217 277614 673500 277616
rect 63217 277611 63283 277614
rect 673494 277612 673500 277614
rect 673564 277612 673570 277676
rect 388253 275906 388319 275909
rect 586053 275906 586119 275909
rect 388253 275904 586119 275906
rect 388253 275848 388258 275904
rect 388314 275848 586058 275904
rect 586114 275848 586119 275904
rect 388253 275846 586119 275848
rect 388253 275843 388319 275846
rect 586053 275843 586119 275846
rect 391289 275770 391355 275773
rect 593137 275770 593203 275773
rect 391289 275768 593203 275770
rect 391289 275712 391294 275768
rect 391350 275712 593142 275768
rect 593198 275712 593203 275768
rect 391289 275710 593203 275712
rect 391289 275707 391355 275710
rect 593137 275707 593203 275710
rect 393589 275634 393655 275637
rect 600221 275634 600287 275637
rect 393589 275632 600287 275634
rect 393589 275576 393594 275632
rect 393650 275576 600226 275632
rect 600282 275576 600287 275632
rect 393589 275574 600287 275576
rect 393589 275571 393655 275574
rect 600221 275571 600287 275574
rect 396257 275498 396323 275501
rect 607305 275498 607371 275501
rect 396257 275496 607371 275498
rect 396257 275440 396262 275496
rect 396318 275440 607310 275496
rect 607366 275440 607371 275496
rect 396257 275438 607371 275440
rect 396257 275435 396323 275438
rect 607305 275435 607371 275438
rect 398925 275362 398991 275365
rect 614389 275362 614455 275365
rect 398925 275360 614455 275362
rect 398925 275304 398930 275360
rect 398986 275304 614394 275360
rect 614450 275304 614455 275360
rect 398925 275302 614455 275304
rect 398925 275299 398991 275302
rect 614389 275299 614455 275302
rect 401685 275226 401751 275229
rect 621473 275226 621539 275229
rect 401685 275224 621539 275226
rect 401685 275168 401690 275224
rect 401746 275168 621478 275224
rect 621534 275168 621539 275224
rect 401685 275166 621539 275168
rect 401685 275163 401751 275166
rect 621473 275163 621539 275166
rect 404261 275090 404327 275093
rect 628557 275090 628623 275093
rect 404261 275088 628623 275090
rect 404261 275032 404266 275088
rect 404322 275032 628562 275088
rect 628618 275032 628623 275088
rect 404261 275030 628623 275032
rect 404261 275027 404327 275030
rect 628557 275027 628623 275030
rect 402697 274954 402763 274957
rect 623865 274954 623931 274957
rect 402697 274952 623931 274954
rect 402697 274896 402702 274952
rect 402758 274896 623870 274952
rect 623926 274896 623931 274952
rect 402697 274894 623931 274896
rect 402697 274891 402763 274894
rect 623865 274891 623931 274894
rect 405365 274818 405431 274821
rect 630949 274818 631015 274821
rect 405365 274816 631015 274818
rect 405365 274760 405370 274816
rect 405426 274760 630954 274816
rect 631010 274760 631015 274816
rect 405365 274758 631015 274760
rect 405365 274755 405431 274758
rect 630949 274755 631015 274758
rect 406929 274682 406995 274685
rect 635641 274682 635707 274685
rect 406929 274680 635707 274682
rect 406929 274624 406934 274680
rect 406990 274624 635646 274680
rect 635702 274624 635707 274680
rect 406929 274622 635707 274624
rect 406929 274619 406995 274622
rect 635641 274619 635707 274622
rect 408217 274546 408283 274549
rect 638033 274546 638099 274549
rect 408217 274544 638099 274546
rect 408217 274488 408222 274544
rect 408278 274488 638038 274544
rect 638094 274488 638099 274544
rect 408217 274486 638099 274488
rect 408217 274483 408283 274486
rect 638033 274483 638099 274486
rect 111977 273186 112043 273189
rect 209221 273186 209287 273189
rect 111977 273184 209287 273186
rect 111977 273128 111982 273184
rect 112038 273128 209226 273184
rect 209282 273128 209287 273184
rect 111977 273126 209287 273128
rect 111977 273123 112043 273126
rect 209221 273123 209287 273126
rect 368657 273186 368723 273189
rect 533981 273186 534047 273189
rect 368657 273184 534047 273186
rect 368657 273128 368662 273184
rect 368718 273128 533986 273184
rect 534042 273128 534047 273184
rect 368657 273126 534047 273128
rect 368657 273123 368723 273126
rect 533981 273123 534047 273126
rect 107193 273050 107259 273053
rect 203425 273050 203491 273053
rect 107193 273048 203491 273050
rect 107193 272992 107198 273048
rect 107254 272992 203430 273048
rect 203486 272992 203491 273048
rect 107193 272990 203491 272992
rect 107193 272987 107259 272990
rect 203425 272987 203491 272990
rect 371233 273050 371299 273053
rect 539869 273050 539935 273053
rect 371233 273048 539935 273050
rect 371233 272992 371238 273048
rect 371294 272992 539874 273048
rect 539930 272992 539935 273048
rect 371233 272990 539935 272992
rect 371233 272987 371299 272990
rect 539869 272987 539935 272990
rect 105997 272914 106063 272917
rect 207473 272914 207539 272917
rect 105997 272912 207539 272914
rect 105997 272856 106002 272912
rect 106058 272856 207478 272912
rect 207534 272856 207539 272912
rect 105997 272854 207539 272856
rect 105997 272851 106063 272854
rect 207473 272851 207539 272854
rect 371325 272914 371391 272917
rect 541065 272914 541131 272917
rect 371325 272912 541131 272914
rect 371325 272856 371330 272912
rect 371386 272856 541070 272912
rect 541126 272856 541131 272912
rect 371325 272854 541131 272856
rect 371325 272851 371391 272854
rect 541065 272851 541131 272854
rect 97717 272778 97783 272781
rect 201309 272778 201375 272781
rect 97717 272776 201375 272778
rect 97717 272720 97722 272776
rect 97778 272720 201314 272776
rect 201370 272720 201375 272776
rect 97717 272718 201375 272720
rect 97717 272715 97783 272718
rect 201309 272715 201375 272718
rect 373993 272778 374059 272781
rect 548149 272778 548215 272781
rect 373993 272776 548215 272778
rect 373993 272720 373998 272776
rect 374054 272720 548154 272776
rect 548210 272720 548215 272776
rect 373993 272718 548215 272720
rect 373993 272715 374059 272718
rect 548149 272715 548215 272718
rect 100109 272642 100175 272645
rect 205725 272642 205791 272645
rect 100109 272640 205791 272642
rect 100109 272584 100114 272640
rect 100170 272584 205730 272640
rect 205786 272584 205791 272640
rect 100109 272582 205791 272584
rect 100109 272579 100175 272582
rect 205725 272579 205791 272582
rect 379329 272642 379395 272645
rect 562409 272642 562475 272645
rect 379329 272640 562475 272642
rect 379329 272584 379334 272640
rect 379390 272584 562414 272640
rect 562470 272584 562475 272640
rect 379329 272582 562475 272584
rect 379329 272579 379395 272582
rect 562409 272579 562475 272582
rect 98913 272506 98979 272509
rect 204805 272506 204871 272509
rect 98913 272504 204871 272506
rect 98913 272448 98918 272504
rect 98974 272448 204810 272504
rect 204866 272448 204871 272504
rect 98913 272446 204871 272448
rect 98913 272443 98979 272446
rect 204805 272443 204871 272446
rect 392761 272506 392827 272509
rect 597829 272506 597895 272509
rect 392761 272504 597895 272506
rect 392761 272448 392766 272504
rect 392822 272448 597834 272504
rect 597890 272448 597895 272504
rect 392761 272446 597895 272448
rect 392761 272443 392827 272446
rect 597829 272443 597895 272446
rect 41965 272372 42031 272373
rect 41965 272368 42012 272372
rect 42076 272370 42082 272372
rect 91829 272370 91895 272373
rect 202137 272370 202203 272373
rect 41965 272312 41970 272368
rect 41965 272308 42012 272312
rect 42076 272310 42122 272370
rect 91829 272368 202203 272370
rect 91829 272312 91834 272368
rect 91890 272312 202142 272368
rect 202198 272312 202203 272368
rect 91829 272310 202203 272312
rect 42076 272308 42082 272310
rect 41965 272307 42031 272308
rect 91829 272307 91895 272310
rect 202137 272307 202203 272310
rect 398097 272370 398163 272373
rect 611997 272370 612063 272373
rect 398097 272368 612063 272370
rect 398097 272312 398102 272368
rect 398158 272312 612002 272368
rect 612058 272312 612063 272368
rect 398097 272310 612063 272312
rect 398097 272307 398163 272310
rect 611997 272307 612063 272310
rect 85941 272234 86007 272237
rect 199929 272234 199995 272237
rect 85941 272232 199995 272234
rect 85941 272176 85946 272232
rect 86002 272176 199934 272232
rect 199990 272176 199995 272232
rect 85941 272174 199995 272176
rect 85941 272171 86007 272174
rect 199929 272171 199995 272174
rect 403433 272234 403499 272237
rect 626165 272234 626231 272237
rect 403433 272232 626231 272234
rect 403433 272176 403438 272232
rect 403494 272176 626170 272232
rect 626226 272176 626231 272232
rect 403433 272174 626231 272176
rect 403433 272171 403499 272174
rect 626165 272171 626231 272174
rect 83549 272098 83615 272101
rect 199101 272098 199167 272101
rect 83549 272096 199167 272098
rect 83549 272040 83554 272096
rect 83610 272040 199106 272096
rect 199162 272040 199167 272096
rect 83549 272038 199167 272040
rect 83549 272035 83615 272038
rect 199101 272035 199167 272038
rect 408769 272098 408835 272101
rect 640425 272098 640491 272101
rect 408769 272096 640491 272098
rect 408769 272040 408774 272096
rect 408830 272040 640430 272096
rect 640486 272040 640491 272096
rect 408769 272038 640491 272040
rect 408769 272035 408835 272038
rect 640425 272035 640491 272038
rect 76465 271962 76531 271965
rect 196341 271962 196407 271965
rect 76465 271960 196407 271962
rect 76465 271904 76470 271960
rect 76526 271904 196346 271960
rect 196402 271904 196407 271960
rect 76465 271902 196407 271904
rect 76465 271899 76531 271902
rect 196341 271899 196407 271902
rect 410885 271962 410951 271965
rect 645117 271962 645183 271965
rect 410885 271960 645183 271962
rect 410885 271904 410890 271960
rect 410946 271904 645122 271960
rect 645178 271904 645183 271960
rect 410885 271902 645183 271904
rect 410885 271899 410951 271902
rect 645117 271899 645183 271902
rect 70577 271826 70643 271829
rect 194133 271826 194199 271829
rect 70577 271824 194199 271826
rect 70577 271768 70582 271824
rect 70638 271768 194138 271824
rect 194194 271768 194199 271824
rect 70577 271766 194199 271768
rect 70577 271763 70643 271766
rect 194133 271763 194199 271766
rect 194501 271826 194567 271829
rect 208485 271826 208551 271829
rect 194501 271824 208551 271826
rect 194501 271768 194506 271824
rect 194562 271768 208490 271824
rect 208546 271768 208551 271824
rect 194501 271766 208551 271768
rect 194501 271763 194567 271766
rect 208485 271763 208551 271766
rect 411069 271826 411135 271829
rect 646313 271826 646379 271829
rect 411069 271824 646379 271826
rect 411069 271768 411074 271824
rect 411130 271768 646318 271824
rect 646374 271768 646379 271824
rect 411069 271766 646379 271768
rect 411069 271763 411135 271766
rect 646313 271763 646379 271766
rect 115473 271690 115539 271693
rect 210601 271690 210667 271693
rect 115473 271688 210667 271690
rect 115473 271632 115478 271688
rect 115534 271632 210606 271688
rect 210662 271632 210667 271688
rect 115473 271630 210667 271632
rect 115473 271627 115539 271630
rect 210601 271627 210667 271630
rect 365529 271690 365595 271693
rect 525701 271690 525767 271693
rect 365529 271688 525767 271690
rect 365529 271632 365534 271688
rect 365590 271632 525706 271688
rect 525762 271632 525767 271688
rect 365529 271630 525767 271632
rect 365529 271627 365595 271630
rect 525701 271627 525767 271630
rect 122557 271554 122623 271557
rect 213269 271554 213335 271557
rect 122557 271552 213335 271554
rect 122557 271496 122562 271552
rect 122618 271496 213274 271552
rect 213330 271496 213335 271552
rect 122557 271494 213335 271496
rect 122557 271491 122623 271494
rect 213269 271491 213335 271494
rect 365989 271554 366055 271557
rect 526897 271554 526963 271557
rect 365989 271552 526963 271554
rect 365989 271496 365994 271552
rect 366050 271496 526902 271552
rect 526958 271496 526963 271552
rect 365989 271494 526963 271496
rect 365989 271491 366055 271494
rect 526897 271491 526963 271494
rect 363321 271418 363387 271421
rect 519813 271418 519879 271421
rect 363321 271416 519879 271418
rect 363321 271360 363326 271416
rect 363382 271360 519818 271416
rect 519874 271360 519879 271416
rect 363321 271358 519879 271360
rect 363321 271355 363387 271358
rect 519813 271355 519879 271358
rect 42149 270466 42215 270469
rect 42374 270466 42380 270468
rect 42149 270464 42380 270466
rect 42149 270408 42154 270464
rect 42210 270408 42380 270464
rect 42149 270406 42380 270408
rect 42149 270403 42215 270406
rect 42374 270404 42380 270406
rect 42444 270404 42450 270468
rect 121361 270466 121427 270469
rect 213729 270466 213795 270469
rect 121361 270464 213795 270466
rect 121361 270408 121366 270464
rect 121422 270408 213734 270464
rect 213790 270408 213795 270464
rect 121361 270406 213795 270408
rect 121361 270403 121427 270406
rect 213729 270403 213795 270406
rect 366909 270466 366975 270469
rect 529289 270466 529355 270469
rect 366909 270464 529355 270466
rect 366909 270408 366914 270464
rect 366970 270408 529294 270464
rect 529350 270408 529355 270464
rect 366909 270406 529355 270408
rect 366909 270403 366975 270406
rect 529289 270403 529355 270406
rect 108389 270330 108455 270333
rect 207933 270330 207999 270333
rect 108389 270328 207999 270330
rect 108389 270272 108394 270328
rect 108450 270272 207938 270328
rect 207994 270272 207999 270328
rect 108389 270270 207999 270272
rect 108389 270267 108455 270270
rect 207933 270267 207999 270270
rect 369577 270330 369643 270333
rect 536373 270330 536439 270333
rect 369577 270328 536439 270330
rect 369577 270272 369582 270328
rect 369638 270272 536378 270328
rect 536434 270272 536439 270328
rect 369577 270270 536439 270272
rect 369577 270267 369643 270270
rect 536373 270267 536439 270270
rect 103697 270194 103763 270197
rect 207013 270194 207079 270197
rect 103697 270192 207079 270194
rect 103697 270136 103702 270192
rect 103758 270136 207018 270192
rect 207074 270136 207079 270192
rect 103697 270134 207079 270136
rect 103697 270131 103763 270134
rect 207013 270131 207079 270134
rect 372245 270194 372311 270197
rect 543457 270194 543523 270197
rect 372245 270192 543523 270194
rect 372245 270136 372250 270192
rect 372306 270136 543462 270192
rect 543518 270136 543523 270192
rect 372245 270134 543523 270136
rect 372245 270131 372311 270134
rect 543457 270131 543523 270134
rect 42149 270060 42215 270061
rect 42149 270058 42196 270060
rect 42104 270056 42196 270058
rect 42104 270000 42154 270056
rect 42104 269998 42196 270000
rect 42149 269996 42196 269998
rect 42260 269996 42266 270060
rect 101305 270058 101371 270061
rect 205265 270058 205331 270061
rect 101305 270056 205331 270058
rect 101305 270000 101310 270056
rect 101366 270000 205270 270056
rect 205326 270000 205331 270056
rect 101305 269998 205331 270000
rect 42149 269995 42215 269996
rect 101305 269995 101371 269998
rect 205265 269995 205331 269998
rect 378041 270058 378107 270061
rect 558821 270058 558887 270061
rect 378041 270056 558887 270058
rect 378041 270000 378046 270056
rect 378102 270000 558826 270056
rect 558882 270000 558887 270056
rect 378041 269998 558887 270000
rect 378041 269995 378107 269998
rect 558821 269995 558887 269998
rect 96613 269922 96679 269925
rect 204345 269922 204411 269925
rect 96613 269920 204411 269922
rect 96613 269864 96618 269920
rect 96674 269864 204350 269920
rect 204406 269864 204411 269920
rect 96613 269862 204411 269864
rect 96613 269859 96679 269862
rect 204345 269859 204411 269862
rect 383377 269922 383443 269925
rect 572989 269922 573055 269925
rect 383377 269920 573055 269922
rect 383377 269864 383382 269920
rect 383438 269864 572994 269920
rect 573050 269864 573055 269920
rect 383377 269862 573055 269864
rect 383377 269859 383443 269862
rect 572989 269859 573055 269862
rect 87137 269786 87203 269789
rect 200389 269786 200455 269789
rect 87137 269784 200455 269786
rect 87137 269728 87142 269784
rect 87198 269728 200394 269784
rect 200450 269728 200455 269784
rect 87137 269726 200455 269728
rect 87137 269723 87203 269726
rect 200389 269723 200455 269726
rect 391381 269786 391447 269789
rect 594333 269786 594399 269789
rect 391381 269784 594399 269786
rect 391381 269728 391386 269784
rect 391442 269728 594338 269784
rect 594394 269728 594399 269784
rect 391381 269726 594399 269728
rect 391381 269723 391447 269726
rect 594333 269723 594399 269726
rect 90633 269650 90699 269653
rect 201677 269650 201743 269653
rect 90633 269648 201743 269650
rect 90633 269592 90638 269648
rect 90694 269592 201682 269648
rect 201738 269592 201743 269648
rect 90633 269590 201743 269592
rect 90633 269587 90699 269590
rect 201677 269587 201743 269590
rect 402053 269650 402119 269653
rect 622669 269650 622735 269653
rect 402053 269648 622735 269650
rect 402053 269592 402058 269648
rect 402114 269592 622674 269648
rect 622730 269592 622735 269648
rect 402053 269590 622735 269592
rect 402053 269587 402119 269590
rect 622669 269587 622735 269590
rect 84745 269514 84811 269517
rect 199009 269514 199075 269517
rect 84745 269512 199075 269514
rect 84745 269456 84750 269512
rect 84806 269456 199014 269512
rect 199070 269456 199075 269512
rect 84745 269454 199075 269456
rect 84745 269451 84811 269454
rect 199009 269451 199075 269454
rect 404721 269514 404787 269517
rect 629753 269514 629819 269517
rect 404721 269512 629819 269514
rect 404721 269456 404726 269512
rect 404782 269456 629758 269512
rect 629814 269456 629819 269512
rect 404721 269454 629819 269456
rect 404721 269451 404787 269454
rect 629753 269451 629819 269454
rect 78857 269378 78923 269381
rect 197721 269378 197787 269381
rect 78857 269376 197787 269378
rect 78857 269320 78862 269376
rect 78918 269320 197726 269376
rect 197782 269320 197787 269376
rect 78857 269318 197787 269320
rect 78857 269315 78923 269318
rect 197721 269315 197787 269318
rect 407389 269378 407455 269381
rect 636837 269378 636903 269381
rect 407389 269376 636903 269378
rect 407389 269320 407394 269376
rect 407450 269320 636842 269376
rect 636898 269320 636903 269376
rect 407389 269318 636903 269320
rect 407389 269315 407455 269318
rect 636837 269315 636903 269318
rect 42149 269242 42215 269245
rect 42558 269242 42564 269244
rect 42149 269240 42564 269242
rect 42149 269184 42154 269240
rect 42210 269184 42564 269240
rect 42149 269182 42564 269184
rect 42149 269179 42215 269182
rect 42558 269180 42564 269182
rect 42628 269180 42634 269244
rect 77661 269242 77727 269245
rect 196801 269242 196867 269245
rect 77661 269240 196867 269242
rect 77661 269184 77666 269240
rect 77722 269184 196806 269240
rect 196862 269184 196867 269240
rect 77661 269182 196867 269184
rect 77661 269179 77727 269182
rect 196801 269179 196867 269182
rect 409597 269242 409663 269245
rect 642725 269242 642791 269245
rect 409597 269240 642791 269242
rect 409597 269184 409602 269240
rect 409658 269184 642730 269240
rect 642786 269184 642791 269240
rect 409597 269182 642791 269184
rect 409597 269179 409663 269182
rect 642725 269179 642791 269182
rect 69381 269106 69447 269109
rect 193673 269106 193739 269109
rect 69381 269104 193739 269106
rect 69381 269048 69386 269104
rect 69442 269048 193678 269104
rect 193734 269048 193739 269104
rect 69381 269046 193739 269048
rect 69381 269043 69447 269046
rect 193673 269043 193739 269046
rect 410057 269106 410123 269109
rect 643921 269106 643987 269109
rect 410057 269104 643987 269106
rect 410057 269048 410062 269104
rect 410118 269048 643926 269104
rect 643982 269048 643987 269104
rect 410057 269046 643987 269048
rect 410057 269043 410123 269046
rect 643921 269043 643987 269046
rect 128537 268970 128603 268973
rect 216397 268970 216463 268973
rect 128537 268968 216463 268970
rect 128537 268912 128542 268968
rect 128598 268912 216402 268968
rect 216458 268912 216463 268968
rect 128537 268910 216463 268912
rect 128537 268907 128603 268910
rect 216397 268907 216463 268910
rect 364241 268970 364307 268973
rect 522205 268970 522271 268973
rect 364241 268968 522271 268970
rect 364241 268912 364246 268968
rect 364302 268912 522210 268968
rect 522266 268912 522271 268968
rect 364241 268910 522271 268912
rect 364241 268907 364307 268910
rect 522205 268907 522271 268910
rect 127341 268834 127407 268837
rect 215477 268834 215543 268837
rect 127341 268832 215543 268834
rect 127341 268776 127346 268832
rect 127402 268776 215482 268832
rect 215538 268776 215543 268832
rect 127341 268774 215543 268776
rect 127341 268771 127407 268774
rect 215477 268771 215543 268774
rect 362033 268834 362099 268837
rect 516225 268834 516291 268837
rect 362033 268832 516291 268834
rect 362033 268776 362038 268832
rect 362094 268776 516230 268832
rect 516286 268776 516291 268832
rect 362033 268774 516291 268776
rect 362033 268771 362099 268774
rect 516225 268771 516291 268774
rect 142705 268698 142771 268701
rect 221733 268698 221799 268701
rect 142705 268696 221799 268698
rect 142705 268640 142710 268696
rect 142766 268640 221738 268696
rect 221794 268640 221799 268696
rect 142705 268638 221799 268640
rect 142705 268635 142771 268638
rect 221733 268635 221799 268638
rect 358905 268698 358971 268701
rect 507945 268698 508011 268701
rect 358905 268696 508011 268698
rect 358905 268640 358910 268696
rect 358966 268640 507950 268696
rect 508006 268640 508011 268696
rect 358905 268638 508011 268640
rect 358905 268635 358971 268638
rect 507945 268635 508011 268638
rect 153285 268562 153351 268565
rect 225781 268562 225847 268565
rect 153285 268560 225847 268562
rect 153285 268504 153290 268560
rect 153346 268504 225786 268560
rect 225842 268504 225847 268560
rect 153285 268502 225847 268504
rect 153285 268499 153351 268502
rect 225781 268499 225847 268502
rect 359365 268562 359431 268565
rect 509141 268562 509207 268565
rect 359365 268560 509207 268562
rect 359365 268504 359370 268560
rect 359426 268504 509146 268560
rect 509202 268504 509207 268560
rect 359365 268502 509207 268504
rect 359365 268499 359431 268502
rect 509141 268499 509207 268502
rect 676121 268562 676187 268565
rect 676262 268562 676322 268668
rect 676121 268560 676322 268562
rect 676121 268504 676126 268560
rect 676182 268504 676322 268560
rect 676121 268502 676322 268504
rect 676121 268499 676187 268502
rect 184933 268426 184999 268429
rect 203057 268426 203123 268429
rect 184933 268424 203123 268426
rect 184933 268368 184938 268424
rect 184994 268368 203062 268424
rect 203118 268368 203123 268424
rect 184933 268366 203123 268368
rect 184933 268363 184999 268366
rect 203057 268363 203123 268366
rect 356605 268426 356671 268429
rect 502057 268426 502123 268429
rect 356605 268424 502123 268426
rect 356605 268368 356610 268424
rect 356666 268368 502062 268424
rect 502118 268368 502123 268424
rect 356605 268366 502123 268368
rect 356605 268363 356671 268366
rect 502057 268363 502123 268366
rect 353937 268290 354003 268293
rect 494973 268290 495039 268293
rect 353937 268288 495039 268290
rect 353937 268232 353942 268288
rect 353998 268232 494978 268288
rect 495034 268232 495039 268288
rect 353937 268230 495039 268232
rect 353937 268227 354003 268230
rect 494973 268227 495039 268230
rect 676262 268157 676322 268260
rect 203425 268154 203491 268157
rect 208393 268154 208459 268157
rect 203425 268152 208459 268154
rect 203425 268096 203430 268152
rect 203486 268096 208398 268152
rect 208454 268096 208459 268152
rect 203425 268094 208459 268096
rect 203425 268091 203491 268094
rect 208393 268091 208459 268094
rect 676213 268152 676322 268157
rect 676213 268096 676218 268152
rect 676274 268096 676322 268152
rect 676213 268094 676322 268096
rect 676213 268091 676279 268094
rect 676029 267882 676095 267885
rect 676029 267880 676292 267882
rect 676029 267824 676034 267880
rect 676090 267824 676292 267880
rect 676029 267822 676292 267824
rect 676029 267819 676095 267822
rect 387793 267746 387859 267749
rect 584857 267746 584923 267749
rect 387793 267744 584923 267746
rect 387793 267688 387798 267744
rect 387854 267688 584862 267744
rect 584918 267688 584923 267744
rect 387793 267686 584923 267688
rect 387793 267683 387859 267686
rect 584857 267683 584923 267686
rect 386965 267610 387031 267613
rect 582465 267610 582531 267613
rect 386965 267608 582531 267610
rect 386965 267552 386970 267608
rect 387026 267552 582470 267608
rect 582526 267552 582531 267608
rect 386965 267550 582531 267552
rect 386965 267547 387031 267550
rect 582465 267547 582531 267550
rect 389633 267474 389699 267477
rect 589549 267474 589615 267477
rect 389633 267472 589615 267474
rect 389633 267416 389638 267472
rect 389694 267416 589554 267472
rect 589610 267416 589615 267472
rect 389633 267414 589615 267416
rect 389633 267411 389699 267414
rect 589549 267411 589615 267414
rect 675937 267474 676003 267477
rect 675937 267472 676292 267474
rect 675937 267416 675942 267472
rect 675998 267416 676292 267472
rect 675937 267414 676292 267416
rect 675937 267411 676003 267414
rect 390461 267338 390527 267341
rect 591941 267338 592007 267341
rect 390461 267336 592007 267338
rect 390461 267280 390466 267336
rect 390522 267280 591946 267336
rect 592002 267280 592007 267336
rect 390461 267278 592007 267280
rect 390461 267275 390527 267278
rect 591941 267275 592007 267278
rect 391841 267202 391907 267205
rect 595437 267202 595503 267205
rect 391841 267200 595503 267202
rect 391841 267144 391846 267200
rect 391902 267144 595442 267200
rect 595498 267144 595503 267200
rect 391841 267142 595503 267144
rect 391841 267139 391907 267142
rect 595437 267139 595503 267142
rect 393129 267066 393195 267069
rect 599025 267066 599091 267069
rect 393129 267064 599091 267066
rect 393129 267008 393134 267064
rect 393190 267008 599030 267064
rect 599086 267008 599091 267064
rect 393129 267006 599091 267008
rect 393129 267003 393195 267006
rect 599025 267003 599091 267006
rect 675753 267066 675819 267069
rect 675753 267064 676292 267066
rect 675753 267008 675758 267064
rect 675814 267008 676292 267064
rect 675753 267006 676292 267008
rect 675753 267003 675819 267006
rect 394509 266930 394575 266933
rect 602521 266930 602587 266933
rect 394509 266928 602587 266930
rect 394509 266872 394514 266928
rect 394570 266872 602526 266928
rect 602582 266872 602587 266928
rect 394509 266870 602587 266872
rect 394509 266867 394575 266870
rect 602521 266867 602587 266870
rect 395797 266794 395863 266797
rect 606109 266794 606175 266797
rect 395797 266792 606175 266794
rect 395797 266736 395802 266792
rect 395858 266736 606114 266792
rect 606170 266736 606175 266792
rect 395797 266734 606175 266736
rect 395797 266731 395863 266734
rect 606109 266731 606175 266734
rect 397177 266658 397243 266661
rect 609697 266658 609763 266661
rect 397177 266656 609763 266658
rect 397177 266600 397182 266656
rect 397238 266600 609702 266656
rect 609758 266600 609763 266656
rect 397177 266598 609763 266600
rect 397177 266595 397243 266598
rect 609697 266595 609763 266598
rect 676029 266658 676095 266661
rect 676029 266656 676292 266658
rect 676029 266600 676034 266656
rect 676090 266600 676292 266656
rect 676029 266598 676292 266600
rect 676029 266595 676095 266598
rect 398465 266522 398531 266525
rect 613193 266522 613259 266525
rect 398465 266520 613259 266522
rect 398465 266464 398470 266520
rect 398526 266464 613198 266520
rect 613254 266464 613259 266520
rect 398465 266462 613259 266464
rect 398465 266459 398531 266462
rect 613193 266459 613259 266462
rect 399845 266386 399911 266389
rect 616781 266386 616847 266389
rect 399845 266384 616847 266386
rect 399845 266328 399850 266384
rect 399906 266328 616786 266384
rect 616842 266328 616847 266384
rect 399845 266326 616847 266328
rect 399845 266323 399911 266326
rect 616781 266323 616847 266326
rect 386505 266250 386571 266253
rect 581269 266250 581335 266253
rect 386505 266248 581335 266250
rect 386505 266192 386510 266248
rect 386566 266192 581274 266248
rect 581330 266192 581335 266248
rect 386505 266190 581335 266192
rect 386505 266187 386571 266190
rect 581269 266187 581335 266190
rect 676029 266250 676095 266253
rect 676029 266248 676292 266250
rect 676029 266192 676034 266248
rect 676090 266192 676292 266248
rect 676029 266190 676292 266192
rect 676029 266187 676095 266190
rect 385125 266114 385191 266117
rect 577773 266114 577839 266117
rect 385125 266112 577839 266114
rect 385125 266056 385130 266112
rect 385186 266056 577778 266112
rect 577834 266056 577839 266112
rect 385125 266054 577839 266056
rect 385125 266051 385191 266054
rect 577773 266051 577839 266054
rect 676213 266114 676279 266117
rect 676213 266112 676322 266114
rect 676213 266056 676218 266112
rect 676274 266056 676322 266112
rect 676213 266051 676322 266056
rect 405457 265978 405523 265981
rect 465901 265978 465967 265981
rect 405457 265976 465967 265978
rect 405457 265920 405462 265976
rect 405518 265920 465906 265976
rect 465962 265920 465967 265976
rect 405457 265918 465967 265920
rect 405457 265915 405523 265918
rect 465901 265915 465967 265918
rect 408309 265842 408375 265845
rect 459461 265842 459527 265845
rect 408309 265840 459527 265842
rect 408309 265784 408314 265840
rect 408370 265784 459466 265840
rect 459522 265784 459527 265840
rect 676262 265812 676322 266051
rect 408309 265782 459527 265784
rect 408309 265779 408375 265782
rect 459461 265779 459527 265782
rect 675661 265434 675727 265437
rect 675661 265432 676292 265434
rect 675661 265376 675666 265432
rect 675722 265376 676292 265432
rect 675661 265374 676292 265376
rect 675661 265371 675727 265374
rect 676262 264893 676322 264996
rect 676213 264888 676322 264893
rect 676213 264832 676218 264888
rect 676274 264832 676322 264888
rect 676213 264830 676322 264832
rect 676213 264827 676279 264830
rect 674230 264556 674236 264620
rect 674300 264618 674306 264620
rect 674300 264558 676292 264618
rect 674300 264556 674306 264558
rect 676029 264210 676095 264213
rect 676029 264208 676292 264210
rect 676029 264152 676034 264208
rect 676090 264152 676292 264208
rect 676029 264150 676292 264152
rect 676029 264147 676095 264150
rect 676121 263666 676187 263669
rect 676262 263666 676322 263772
rect 676121 263664 676322 263666
rect 676121 263608 676126 263664
rect 676182 263608 676322 263664
rect 676121 263606 676322 263608
rect 676121 263603 676187 263606
rect 675845 263394 675911 263397
rect 675845 263392 676292 263394
rect 675845 263336 675850 263392
rect 675906 263336 676292 263392
rect 675845 263334 676292 263336
rect 675845 263331 675911 263334
rect 676029 262986 676095 262989
rect 676029 262984 676292 262986
rect 676029 262928 676034 262984
rect 676090 262928 676292 262984
rect 676029 262926 676292 262928
rect 676029 262923 676095 262926
rect 418061 262714 418127 262717
rect 412436 262712 418127 262714
rect 412436 262656 418066 262712
rect 418122 262656 418127 262712
rect 412436 262654 418127 262656
rect 418061 262651 418127 262654
rect 675937 262578 676003 262581
rect 675937 262576 676292 262578
rect 675937 262520 675942 262576
rect 675998 262520 676292 262576
rect 675937 262518 676292 262520
rect 675937 262515 676003 262518
rect 658181 262442 658247 262445
rect 674230 262442 674236 262444
rect 658181 262440 674236 262442
rect 658181 262384 658186 262440
rect 658242 262384 674236 262440
rect 658181 262382 674236 262384
rect 658181 262379 658247 262382
rect 674230 262380 674236 262382
rect 674300 262442 674306 262444
rect 676070 262442 676076 262444
rect 674300 262382 676076 262442
rect 674300 262380 674306 262382
rect 676070 262380 676076 262382
rect 676140 262380 676146 262444
rect 676029 262170 676095 262173
rect 676029 262168 676292 262170
rect 676029 262112 676034 262168
rect 676090 262112 676292 262168
rect 676029 262110 676292 262112
rect 676029 262107 676095 262110
rect 676029 261762 676095 261765
rect 676029 261760 676292 261762
rect 676029 261704 676034 261760
rect 676090 261704 676292 261760
rect 676029 261702 676292 261704
rect 676029 261699 676095 261702
rect 676121 261218 676187 261221
rect 676262 261218 676322 261324
rect 676121 261216 676322 261218
rect 676121 261160 676126 261216
rect 676182 261160 676322 261216
rect 676121 261158 676322 261160
rect 676121 261155 676187 261158
rect 675937 260946 676003 260949
rect 675937 260944 676292 260946
rect 675937 260888 675942 260944
rect 675998 260888 676292 260944
rect 675937 260886 676292 260888
rect 675937 260883 676003 260886
rect 675569 260538 675635 260541
rect 675569 260536 676292 260538
rect 675569 260480 675574 260536
rect 675630 260480 676292 260536
rect 675569 260478 676292 260480
rect 675569 260475 675635 260478
rect 417785 260266 417851 260269
rect 412436 260264 417851 260266
rect 412436 260208 417790 260264
rect 417846 260208 417851 260264
rect 412436 260206 417851 260208
rect 417785 260203 417851 260206
rect 675569 260130 675635 260133
rect 675569 260128 676292 260130
rect 675569 260072 675574 260128
rect 675630 260072 676292 260128
rect 675569 260070 676292 260072
rect 675569 260067 675635 260070
rect 184933 259994 184999 259997
rect 184933 259992 191820 259994
rect 184933 259936 184938 259992
rect 184994 259936 191820 259992
rect 184933 259934 191820 259936
rect 184933 259931 184999 259934
rect 676121 259586 676187 259589
rect 676262 259586 676322 259692
rect 676121 259584 676322 259586
rect 676121 259528 676126 259584
rect 676182 259528 676322 259584
rect 676121 259526 676322 259528
rect 676121 259523 676187 259526
rect 676029 259314 676095 259317
rect 676029 259312 676292 259314
rect 676029 259256 676034 259312
rect 676090 259256 676292 259312
rect 676029 259254 676292 259256
rect 676029 259251 676095 259254
rect 676121 258770 676187 258773
rect 676262 258770 676322 258876
rect 676121 258768 676322 258770
rect 676121 258712 676126 258768
rect 676182 258712 676322 258768
rect 676121 258710 676322 258712
rect 676121 258707 676187 258710
rect 679022 258365 679082 258468
rect 41505 258362 41571 258365
rect 41462 258360 41571 258362
rect 41462 258304 41510 258360
rect 41566 258304 41571 258360
rect 41462 258299 41571 258304
rect 678973 258360 679082 258365
rect 678973 258304 678978 258360
rect 679034 258304 679082 258360
rect 678973 258302 679082 258304
rect 678973 258299 679039 258302
rect 41462 258060 41522 258299
rect 684542 257957 684602 258060
rect 418337 257954 418403 257957
rect 412436 257952 418403 257954
rect 412436 257896 418342 257952
rect 418398 257896 418403 257952
rect 412436 257894 418403 257896
rect 418337 257891 418403 257894
rect 678973 257954 679039 257957
rect 678973 257952 679082 257954
rect 678973 257896 678978 257952
rect 679034 257896 679082 257952
rect 678973 257891 679082 257896
rect 684493 257952 684602 257957
rect 684493 257896 684498 257952
rect 684554 257896 684602 257952
rect 684493 257894 684602 257896
rect 684493 257891 684559 257894
rect 41781 257682 41847 257685
rect 41492 257680 41847 257682
rect 41492 257624 41786 257680
rect 41842 257624 41847 257680
rect 679022 257652 679082 257891
rect 41492 257622 41847 257624
rect 41781 257619 41847 257622
rect 41505 257546 41571 257549
rect 41462 257544 41571 257546
rect 41462 257488 41510 257544
rect 41566 257488 41571 257544
rect 41462 257483 41571 257488
rect 684493 257546 684559 257549
rect 684493 257544 684602 257546
rect 684493 257488 684498 257544
rect 684554 257488 684602 257544
rect 684493 257483 684602 257488
rect 41462 257244 41522 257483
rect 684542 257244 684602 257483
rect 41781 256866 41847 256869
rect 42190 256866 42196 256868
rect 41492 256864 42196 256866
rect 41492 256808 41786 256864
rect 41842 256808 42196 256864
rect 41492 256806 42196 256808
rect 41781 256803 41847 256806
rect 42190 256804 42196 256806
rect 42260 256804 42266 256868
rect 41462 256324 41522 256428
rect 41454 256260 41460 256324
rect 41524 256260 41530 256324
rect 43529 256050 43595 256053
rect 41492 256048 43595 256050
rect 41492 255992 43534 256048
rect 43590 255992 43595 256048
rect 41492 255990 43595 255992
rect 43529 255987 43595 255990
rect 43437 255642 43503 255645
rect 41492 255640 43503 255642
rect 41492 255584 43442 255640
rect 43498 255584 43503 255640
rect 41492 255582 43503 255584
rect 43437 255579 43503 255582
rect 41454 255444 41460 255508
rect 41524 255444 41530 255508
rect 416773 255506 416839 255509
rect 412436 255504 416839 255506
rect 412436 255448 416778 255504
rect 416834 255448 416839 255504
rect 412436 255446 416839 255448
rect 41462 255234 41522 255444
rect 416773 255443 416839 255446
rect 45921 255234 45987 255237
rect 41462 255232 45987 255234
rect 41462 255204 45926 255232
rect 41492 255176 45926 255204
rect 45982 255176 45987 255232
rect 41492 255174 45987 255176
rect 45921 255171 45987 255174
rect 41638 255098 41644 255100
rect 41462 255038 41644 255098
rect 41462 254796 41522 255038
rect 41638 255036 41644 255038
rect 41708 255036 41714 255100
rect 42006 254418 42012 254420
rect 41492 254358 42012 254418
rect 42006 254356 42012 254358
rect 42076 254418 42082 254420
rect 45737 254418 45803 254421
rect 42076 254416 45803 254418
rect 42076 254360 45742 254416
rect 45798 254360 45803 254416
rect 42076 254358 45803 254360
rect 42076 254356 42082 254358
rect 45737 254355 45803 254358
rect 41822 254010 41828 254012
rect 41492 253950 41828 254010
rect 41822 253948 41828 253950
rect 41892 253948 41898 254012
rect 42701 253602 42767 253605
rect 41492 253600 42767 253602
rect 41492 253544 42706 253600
rect 42762 253544 42767 253600
rect 41492 253542 42767 253544
rect 42701 253539 42767 253542
rect 416773 253194 416839 253197
rect 412436 253192 416839 253194
rect 31710 253061 31770 253164
rect 412436 253136 416778 253192
rect 416834 253136 416839 253192
rect 412436 253134 416839 253136
rect 416773 253131 416839 253134
rect 31661 253056 31770 253061
rect 31661 253000 31666 253056
rect 31722 253000 31770 253056
rect 31661 252998 31770 253000
rect 31661 252995 31727 252998
rect 42006 252786 42012 252788
rect 41492 252726 42012 252786
rect 42006 252724 42012 252726
rect 42076 252724 42082 252788
rect 42885 252378 42951 252381
rect 41492 252376 42951 252378
rect 41492 252320 42890 252376
rect 42946 252320 42951 252376
rect 41492 252318 42951 252320
rect 42885 252315 42951 252318
rect 184933 251970 184999 251973
rect 184933 251968 191820 251970
rect 32998 251837 33058 251940
rect 184933 251912 184938 251968
rect 184994 251912 191820 251968
rect 184933 251910 191820 251912
rect 184933 251907 184999 251910
rect 32998 251832 33107 251837
rect 32998 251776 33046 251832
rect 33102 251776 33107 251832
rect 32998 251774 33107 251776
rect 33041 251771 33107 251774
rect 43713 251562 43779 251565
rect 41492 251560 43779 251562
rect 41492 251504 43718 251560
rect 43774 251504 43779 251560
rect 41492 251502 43779 251504
rect 43713 251499 43779 251502
rect 43805 251154 43871 251157
rect 41492 251152 43871 251154
rect 41492 251096 43810 251152
rect 43866 251096 43871 251152
rect 41492 251094 43871 251096
rect 43805 251091 43871 251094
rect 416773 250746 416839 250749
rect 412436 250744 416839 250746
rect 32814 250613 32874 250716
rect 412436 250688 416778 250744
rect 416834 250688 416839 250744
rect 412436 250686 416839 250688
rect 416773 250683 416839 250686
rect 32765 250608 32874 250613
rect 32765 250552 32770 250608
rect 32826 250552 32874 250608
rect 32765 250550 32874 250552
rect 32765 250547 32831 250550
rect 32814 250205 32874 250308
rect 32814 250200 32923 250205
rect 32814 250144 32862 250200
rect 32918 250144 32923 250200
rect 32814 250142 32923 250144
rect 32857 250139 32923 250142
rect 32998 249797 33058 249900
rect 32949 249792 33058 249797
rect 32949 249736 32954 249792
rect 33010 249736 33058 249792
rect 32949 249734 33058 249736
rect 32949 249731 33015 249734
rect 43253 249522 43319 249525
rect 41492 249520 43319 249522
rect 41492 249464 43258 249520
rect 43314 249464 43319 249520
rect 41492 249462 43319 249464
rect 43253 249459 43319 249462
rect 43345 249114 43411 249117
rect 41492 249112 43411 249114
rect 41492 249056 43350 249112
rect 43406 249056 43411 249112
rect 41492 249054 43411 249056
rect 43345 249051 43411 249054
rect 43069 248706 43135 248709
rect 41492 248704 43135 248706
rect 41492 248648 43074 248704
rect 43130 248648 43135 248704
rect 41492 248646 43135 248648
rect 43069 248643 43135 248646
rect 418061 248298 418127 248301
rect 412436 248296 418127 248298
rect 38334 248165 38394 248268
rect 412436 248240 418066 248296
rect 418122 248240 418127 248296
rect 412436 248238 418127 248240
rect 418061 248235 418127 248238
rect 38285 248160 38394 248165
rect 38285 248104 38290 248160
rect 38346 248104 38394 248160
rect 38285 248102 38394 248104
rect 38285 248099 38351 248102
rect 41462 247757 41522 247860
rect 41462 247752 41571 247757
rect 41462 247696 41510 247752
rect 41566 247696 41571 247752
rect 41462 247694 41571 247696
rect 41505 247691 41571 247694
rect 41462 247349 41522 247452
rect 41462 247344 41571 247349
rect 41462 247288 41510 247344
rect 41566 247288 41571 247344
rect 41462 247286 41571 247288
rect 41505 247283 41571 247286
rect 41462 246941 41522 247044
rect 41462 246936 41571 246941
rect 41462 246880 41510 246936
rect 41566 246880 41571 246936
rect 41462 246878 41571 246880
rect 41505 246875 41571 246878
rect 418429 245986 418495 245989
rect 412436 245984 418495 245986
rect 412436 245928 418434 245984
rect 418490 245928 418495 245984
rect 412436 245926 418495 245928
rect 418429 245923 418495 245926
rect 184933 244082 184999 244085
rect 184933 244080 191820 244082
rect 184933 244024 184938 244080
rect 184994 244024 191820 244080
rect 184933 244022 191820 244024
rect 184933 244019 184999 244022
rect 418153 243538 418219 243541
rect 412436 243536 418219 243538
rect 412436 243480 418158 243536
rect 418214 243480 418219 243536
rect 412436 243478 418219 243480
rect 418153 243475 418219 243478
rect 418521 241226 418587 241229
rect 412436 241224 418587 241226
rect 412436 241168 418526 241224
rect 418582 241168 418587 241224
rect 412436 241166 418587 241168
rect 418521 241163 418587 241166
rect 250161 237282 250227 237285
rect 265709 237282 265775 237285
rect 250161 237280 265775 237282
rect 250161 237224 250166 237280
rect 250222 237224 265714 237280
rect 265770 237224 265775 237280
rect 250161 237222 265775 237224
rect 250161 237219 250227 237222
rect 265709 237219 265775 237222
rect 153101 237146 153167 237149
rect 210049 237146 210115 237149
rect 153101 237144 210115 237146
rect 153101 237088 153106 237144
rect 153162 237088 210054 237144
rect 210110 237088 210115 237144
rect 153101 237086 210115 237088
rect 153101 237083 153167 237086
rect 210049 237083 210115 237086
rect 375833 237146 375899 237149
rect 486417 237146 486483 237149
rect 375833 237144 486483 237146
rect 375833 237088 375838 237144
rect 375894 237088 486422 237144
rect 486478 237088 486483 237144
rect 375833 237086 486483 237088
rect 375833 237083 375899 237086
rect 486417 237083 486483 237086
rect 106181 237010 106247 237013
rect 207565 237010 207631 237013
rect 106181 237008 207631 237010
rect 106181 236952 106186 237008
rect 106242 236952 207570 237008
rect 207626 236952 207631 237008
rect 106181 236950 207631 236952
rect 106181 236947 106247 236950
rect 207565 236947 207631 236950
rect 249885 237010 249951 237013
rect 268561 237010 268627 237013
rect 249885 237008 268627 237010
rect 249885 236952 249890 237008
rect 249946 236952 268566 237008
rect 268622 236952 268627 237008
rect 249885 236950 268627 236952
rect 249885 236947 249951 236950
rect 268561 236947 268627 236950
rect 378317 237010 378383 237013
rect 492305 237010 492371 237013
rect 378317 237008 492371 237010
rect 378317 236952 378322 237008
rect 378378 236952 492310 237008
rect 492366 236952 492371 237008
rect 378317 236950 492371 236952
rect 378317 236947 378383 236950
rect 492305 236947 492371 236950
rect 89621 236874 89687 236877
rect 196985 236874 197051 236877
rect 89621 236872 197051 236874
rect 89621 236816 89626 236872
rect 89682 236816 196990 236872
rect 197046 236816 197051 236872
rect 89621 236814 197051 236816
rect 89621 236811 89687 236814
rect 196985 236811 197051 236814
rect 252553 236874 252619 236877
rect 271413 236874 271479 236877
rect 252553 236872 271479 236874
rect 252553 236816 252558 236872
rect 252614 236816 271418 236872
rect 271474 236816 271479 236872
rect 252553 236814 271479 236816
rect 252553 236811 252619 236814
rect 271413 236811 271479 236814
rect 378685 236874 378751 236877
rect 492581 236874 492647 236877
rect 378685 236872 492647 236874
rect 378685 236816 378690 236872
rect 378746 236816 492586 236872
rect 492642 236816 492647 236872
rect 378685 236814 492647 236816
rect 378685 236811 378751 236814
rect 492581 236811 492647 236814
rect 97901 236738 97967 236741
rect 205817 236738 205883 236741
rect 97901 236736 205883 236738
rect 97901 236680 97906 236736
rect 97962 236680 205822 236736
rect 205878 236680 205883 236736
rect 97901 236678 205883 236680
rect 97901 236675 97967 236678
rect 205817 236675 205883 236678
rect 249701 236738 249767 236741
rect 269941 236738 270007 236741
rect 249701 236736 270007 236738
rect 249701 236680 249706 236736
rect 249762 236680 269946 236736
rect 270002 236680 270007 236736
rect 249701 236678 270007 236680
rect 249701 236675 249767 236678
rect 269941 236675 270007 236678
rect 381169 236738 381235 236741
rect 496997 236738 497063 236741
rect 381169 236736 497063 236738
rect 381169 236680 381174 236736
rect 381230 236680 497002 236736
rect 497058 236680 497063 236736
rect 381169 236678 497063 236680
rect 381169 236675 381235 236678
rect 496997 236675 497063 236678
rect 95141 236602 95207 236605
rect 206185 236602 206251 236605
rect 95141 236600 206251 236602
rect 95141 236544 95146 236600
rect 95202 236544 206190 236600
rect 206246 236544 206251 236600
rect 95141 236542 206251 236544
rect 95141 236539 95207 236542
rect 206185 236539 206251 236542
rect 238753 236602 238819 236605
rect 268193 236602 268259 236605
rect 238753 236600 268259 236602
rect 238753 236544 238758 236600
rect 238814 236544 268198 236600
rect 268254 236544 268259 236600
rect 238753 236542 268259 236544
rect 238753 236539 238819 236542
rect 268193 236539 268259 236542
rect 383653 236602 383719 236605
rect 502701 236602 502767 236605
rect 383653 236600 502767 236602
rect 383653 236544 383658 236600
rect 383714 236544 502706 236600
rect 502762 236544 502767 236600
rect 383653 236542 502767 236544
rect 383653 236539 383719 236542
rect 502701 236539 502767 236542
rect 81341 236466 81407 236469
rect 200481 236466 200547 236469
rect 81341 236464 200547 236466
rect 81341 236408 81346 236464
rect 81402 236408 200486 236464
rect 200542 236408 200547 236464
rect 81341 236406 200547 236408
rect 81341 236403 81407 236406
rect 200481 236403 200547 236406
rect 240041 236466 240107 236469
rect 271781 236466 271847 236469
rect 240041 236464 271847 236466
rect 240041 236408 240046 236464
rect 240102 236408 271786 236464
rect 271842 236408 271847 236464
rect 240041 236406 271847 236408
rect 240041 236403 240107 236406
rect 271781 236403 271847 236406
rect 381537 236466 381603 236469
rect 499941 236466 500007 236469
rect 381537 236464 500007 236466
rect 381537 236408 381542 236464
rect 381598 236408 499946 236464
rect 500002 236408 500007 236464
rect 381537 236406 500007 236408
rect 381537 236403 381603 236406
rect 499941 236403 500007 236406
rect 73061 236330 73127 236333
rect 194409 236330 194475 236333
rect 73061 236328 194475 236330
rect 73061 236272 73066 236328
rect 73122 236272 194414 236328
rect 194470 236272 194475 236328
rect 73061 236270 194475 236272
rect 73061 236267 73127 236270
rect 194409 236267 194475 236270
rect 234521 236330 234587 236333
rect 268929 236330 268995 236333
rect 234521 236328 268995 236330
rect 234521 236272 234526 236328
rect 234582 236272 268934 236328
rect 268990 236272 268995 236328
rect 234521 236270 268995 236272
rect 234521 236267 234587 236270
rect 268929 236267 268995 236270
rect 385861 236330 385927 236333
rect 507853 236330 507919 236333
rect 385861 236328 507919 236330
rect 385861 236272 385866 236328
rect 385922 236272 507858 236328
rect 507914 236272 507919 236328
rect 385861 236270 507919 236272
rect 385861 236267 385927 236270
rect 507853 236267 507919 236270
rect 75821 236194 75887 236197
rect 197629 236194 197695 236197
rect 75821 236192 197695 236194
rect 75821 236136 75826 236192
rect 75882 236136 197634 236192
rect 197690 236136 197695 236192
rect 75821 236134 197695 236136
rect 75821 236131 75887 236134
rect 197629 236131 197695 236134
rect 229001 236194 229067 236197
rect 267089 236194 267155 236197
rect 229001 236192 267155 236194
rect 229001 236136 229006 236192
rect 229062 236136 267094 236192
rect 267150 236136 267155 236192
rect 229001 236134 267155 236136
rect 229001 236131 229067 236134
rect 267089 236131 267155 236134
rect 387977 236194 388043 236197
rect 513741 236194 513807 236197
rect 387977 236192 513807 236194
rect 387977 236136 387982 236192
rect 388038 236136 513746 236192
rect 513802 236136 513807 236192
rect 387977 236134 513807 236136
rect 387977 236131 388043 236134
rect 513741 236131 513807 236134
rect 78581 236058 78647 236061
rect 202965 236058 203031 236061
rect 78581 236056 203031 236058
rect 78581 236000 78586 236056
rect 78642 236000 202970 236056
rect 203026 236000 203031 236056
rect 78581 235998 203031 236000
rect 78581 235995 78647 235998
rect 202965 235995 203031 235998
rect 226241 236058 226307 236061
rect 266077 236058 266143 236061
rect 226241 236056 266143 236058
rect 226241 236000 226246 236056
rect 226302 236000 266082 236056
rect 266138 236000 266143 236056
rect 226241 235998 266143 236000
rect 226241 235995 226307 235998
rect 266077 235995 266143 235998
rect 389081 236058 389147 236061
rect 517421 236058 517487 236061
rect 389081 236056 517487 236058
rect 389081 236000 389086 236056
rect 389142 236000 517426 236056
rect 517482 236000 517487 236056
rect 389081 235998 517487 236000
rect 389081 235995 389147 235998
rect 517421 235995 517487 235998
rect 62021 235922 62087 235925
rect 194777 235922 194843 235925
rect 62021 235920 194843 235922
rect 62021 235864 62026 235920
rect 62082 235864 194782 235920
rect 194838 235864 194843 235920
rect 62021 235862 194843 235864
rect 62021 235859 62087 235862
rect 194777 235859 194843 235862
rect 217685 235922 217751 235925
rect 262857 235922 262923 235925
rect 217685 235920 262923 235922
rect 217685 235864 217690 235920
rect 217746 235864 262862 235920
rect 262918 235864 262923 235920
rect 217685 235862 262923 235864
rect 217685 235859 217751 235862
rect 262857 235859 262923 235862
rect 391197 235922 391263 235925
rect 522941 235922 523007 235925
rect 391197 235920 523007 235922
rect 391197 235864 391202 235920
rect 391258 235864 522946 235920
rect 523002 235864 523007 235920
rect 391197 235862 523007 235864
rect 391197 235859 391263 235862
rect 522941 235859 523007 235862
rect 366541 228850 366607 228853
rect 465073 228850 465139 228853
rect 366541 228848 465139 228850
rect 366541 228792 366546 228848
rect 366602 228792 465078 228848
rect 465134 228792 465139 228848
rect 366541 228790 465139 228792
rect 366541 228787 366607 228790
rect 465073 228787 465139 228790
rect 368013 228714 368079 228717
rect 468385 228714 468451 228717
rect 368013 228712 468451 228714
rect 368013 228656 368018 228712
rect 368074 228656 468390 228712
rect 468446 228656 468451 228712
rect 368013 228654 468451 228656
rect 368013 228651 368079 228654
rect 468385 228651 468451 228654
rect 371233 228578 371299 228581
rect 472617 228578 472683 228581
rect 371233 228576 472683 228578
rect 371233 228520 371238 228576
rect 371294 228520 472622 228576
rect 472678 228520 472683 228576
rect 371233 228518 472683 228520
rect 371233 228515 371299 228518
rect 472617 228515 472683 228518
rect 369761 228442 369827 228445
rect 469213 228442 469279 228445
rect 369761 228440 469279 228442
rect 369761 228384 369766 228440
rect 369822 228384 469218 228440
rect 469274 228384 469279 228440
rect 369761 228382 469279 228384
rect 369761 228379 369827 228382
rect 469213 228379 469279 228382
rect 372613 228306 372679 228309
rect 476021 228306 476087 228309
rect 372613 228304 476087 228306
rect 372613 228248 372618 228304
rect 372674 228248 476026 228304
rect 476082 228248 476087 228304
rect 372613 228246 476087 228248
rect 372613 228243 372679 228246
rect 476021 228243 476087 228246
rect 370865 228170 370931 228173
rect 475101 228170 475167 228173
rect 370865 228168 475167 228170
rect 370865 228112 370870 228168
rect 370926 228112 475106 228168
rect 475162 228112 475167 228168
rect 370865 228110 475167 228112
rect 370865 228107 370931 228110
rect 475101 228107 475167 228110
rect 369393 228034 369459 228037
rect 471973 228034 472039 228037
rect 369393 228032 472039 228034
rect 369393 227976 369398 228032
rect 369454 227976 471978 228032
rect 472034 227976 472039 228032
rect 369393 227974 472039 227976
rect 369393 227971 369459 227974
rect 471973 227971 472039 227974
rect 374085 227898 374151 227901
rect 479333 227898 479399 227901
rect 374085 227896 479399 227898
rect 374085 227840 374090 227896
rect 374146 227840 479338 227896
rect 479394 227840 479399 227896
rect 374085 227838 479399 227840
rect 374085 227835 374151 227838
rect 479333 227835 479399 227838
rect 373717 227762 373783 227765
rect 481909 227762 481975 227765
rect 373717 227760 481975 227762
rect 373717 227704 373722 227760
rect 373778 227704 481914 227760
rect 481970 227704 481975 227760
rect 373717 227702 481975 227704
rect 373717 227699 373783 227702
rect 481909 227699 481975 227702
rect 372245 227626 372311 227629
rect 478505 227626 478571 227629
rect 372245 227624 478571 227626
rect 372245 227568 372250 227624
rect 372306 227568 478510 227624
rect 478566 227568 478571 227624
rect 372245 227566 478571 227568
rect 372245 227563 372311 227566
rect 478505 227563 478571 227566
rect 102041 226130 102107 226133
rect 212809 226130 212875 226133
rect 102041 226128 212875 226130
rect 102041 226072 102046 226128
rect 102102 226072 212814 226128
rect 212870 226072 212875 226128
rect 102041 226070 212875 226072
rect 102041 226067 102107 226070
rect 212809 226067 212875 226070
rect 360929 226130 360995 226133
rect 451549 226130 451615 226133
rect 360929 226128 451615 226130
rect 360929 226072 360934 226128
rect 360990 226072 451554 226128
rect 451610 226072 451615 226128
rect 360929 226070 451615 226072
rect 360929 226067 360995 226070
rect 451549 226067 451615 226070
rect 41965 225996 42031 225997
rect 41965 225992 42012 225996
rect 42076 225994 42082 225996
rect 98913 225994 98979 225997
rect 210877 225994 210943 225997
rect 41965 225936 41970 225992
rect 41965 225932 42012 225936
rect 42076 225934 42122 225994
rect 98913 225992 210943 225994
rect 98913 225936 98918 225992
rect 98974 225936 210882 225992
rect 210938 225936 210943 225992
rect 98913 225934 210943 225936
rect 42076 225932 42082 225934
rect 41965 225931 42031 225932
rect 98913 225931 98979 225934
rect 210877 225931 210943 225934
rect 364057 225994 364123 225997
rect 454953 225994 455019 225997
rect 364057 225992 455019 225994
rect 364057 225936 364062 225992
rect 364118 225936 454958 225992
rect 455014 225936 455019 225992
rect 364057 225934 455019 225936
rect 364057 225931 364123 225934
rect 454953 225931 455019 225934
rect 88885 225858 88951 225861
rect 206645 225858 206711 225861
rect 88885 225856 206711 225858
rect 88885 225800 88890 225856
rect 88946 225800 206650 225856
rect 206706 225800 206711 225856
rect 88885 225798 206711 225800
rect 88885 225795 88951 225798
rect 206645 225795 206711 225798
rect 367001 225858 367067 225861
rect 460013 225858 460079 225861
rect 367001 225856 460079 225858
rect 367001 225800 367006 225856
rect 367062 225800 460018 225856
rect 460074 225800 460079 225856
rect 367001 225798 460079 225800
rect 367001 225795 367067 225798
rect 460013 225795 460079 225798
rect 92197 225722 92263 225725
rect 208025 225722 208091 225725
rect 92197 225720 208091 225722
rect 92197 225664 92202 225720
rect 92258 225664 208030 225720
rect 208086 225664 208091 225720
rect 92197 225662 208091 225664
rect 92197 225659 92263 225662
rect 208025 225659 208091 225662
rect 363689 225722 363755 225725
rect 456609 225722 456675 225725
rect 363689 225720 456675 225722
rect 363689 225664 363694 225720
rect 363750 225664 456614 225720
rect 456670 225664 456675 225720
rect 363689 225662 456675 225664
rect 363689 225659 363755 225662
rect 456609 225659 456675 225662
rect 83825 225586 83891 225589
rect 204805 225586 204871 225589
rect 83825 225584 204871 225586
rect 83825 225528 83830 225584
rect 83886 225528 204810 225584
rect 204866 225528 204871 225584
rect 83825 225526 204871 225528
rect 83825 225523 83891 225526
rect 204805 225523 204871 225526
rect 366357 225586 366423 225589
rect 463693 225586 463759 225589
rect 366357 225584 463759 225586
rect 366357 225528 366362 225584
rect 366418 225528 463698 225584
rect 463754 225528 463759 225584
rect 366357 225526 463759 225528
rect 366357 225523 366423 225526
rect 463693 225523 463759 225526
rect 80421 225450 80487 225453
rect 203425 225450 203491 225453
rect 80421 225448 203491 225450
rect 80421 225392 80426 225448
rect 80482 225392 203430 225448
rect 203486 225392 203491 225448
rect 80421 225390 203491 225392
rect 80421 225387 80487 225390
rect 203425 225387 203491 225390
rect 369117 225450 369183 225453
rect 466729 225450 466795 225453
rect 369117 225448 466795 225450
rect 369117 225392 369122 225448
rect 369178 225392 466734 225448
rect 466790 225392 466795 225448
rect 369117 225390 466795 225392
rect 369117 225387 369183 225390
rect 466729 225387 466795 225390
rect 77109 225314 77175 225317
rect 202045 225314 202111 225317
rect 77109 225312 202111 225314
rect 77109 225256 77114 225312
rect 77170 225256 202050 225312
rect 202106 225256 202111 225312
rect 77109 225254 202111 225256
rect 77109 225251 77175 225254
rect 202045 225251 202111 225254
rect 371969 225314 372035 225317
rect 473445 225314 473511 225317
rect 371969 225312 473511 225314
rect 371969 225256 371974 225312
rect 372030 225256 473450 225312
rect 473506 225256 473511 225312
rect 371969 225254 473511 225256
rect 371969 225251 372035 225254
rect 473445 225251 473511 225254
rect 70393 225178 70459 225181
rect 199101 225178 199167 225181
rect 70393 225176 199167 225178
rect 70393 225120 70398 225176
rect 70454 225120 199106 225176
rect 199162 225120 199167 225176
rect 70393 225118 199167 225120
rect 70393 225115 70459 225118
rect 199101 225115 199167 225118
rect 369209 225178 369275 225181
rect 470133 225178 470199 225181
rect 369209 225176 470199 225178
rect 369209 225120 369214 225176
rect 369270 225120 470138 225176
rect 470194 225120 470199 225176
rect 369209 225118 470199 225120
rect 369209 225115 369275 225118
rect 470133 225115 470199 225118
rect 63401 225042 63467 225045
rect 196249 225042 196315 225045
rect 63401 225040 196315 225042
rect 63401 224984 63406 225040
rect 63462 224984 196254 225040
rect 196310 224984 196315 225040
rect 63401 224982 196315 224984
rect 63401 224979 63467 224982
rect 196249 224979 196315 224982
rect 372061 225042 372127 225045
rect 476849 225042 476915 225045
rect 372061 225040 476915 225042
rect 372061 224984 372066 225040
rect 372122 224984 476854 225040
rect 476910 224984 476915 225040
rect 372061 224982 476915 224984
rect 372061 224979 372127 224982
rect 476849 224979 476915 224982
rect 56869 224906 56935 224909
rect 193397 224906 193463 224909
rect 56869 224904 193463 224906
rect 56869 224848 56874 224904
rect 56930 224848 193402 224904
rect 193458 224848 193463 224904
rect 56869 224846 193463 224848
rect 56869 224843 56935 224846
rect 193397 224843 193463 224846
rect 374729 224906 374795 224909
rect 480253 224906 480319 224909
rect 374729 224904 480319 224906
rect 374729 224848 374734 224904
rect 374790 224848 480258 224904
rect 480314 224848 480319 224904
rect 374729 224846 480319 224848
rect 374729 224843 374795 224846
rect 480253 224843 480319 224846
rect 703997 224362 704063 224365
rect 708965 224362 709031 224365
rect 703997 224360 709031 224362
rect 703997 224304 704002 224360
rect 704058 224304 708970 224360
rect 709026 224304 709031 224360
rect 703997 224302 709031 224304
rect 703997 224299 704063 224302
rect 708965 224299 709031 224302
rect 704457 224226 704523 224229
rect 708505 224226 708571 224229
rect 704457 224224 708571 224226
rect 704457 224168 704462 224224
rect 704518 224168 708510 224224
rect 708566 224168 708571 224224
rect 704457 224166 708571 224168
rect 704457 224163 704523 224166
rect 708505 224163 708571 224166
rect 339309 223546 339375 223549
rect 396901 223546 396967 223549
rect 339309 223544 396967 223546
rect 339309 223488 339314 223544
rect 339370 223488 396906 223544
rect 396962 223488 396967 223544
rect 339309 223486 396967 223488
rect 339309 223483 339375 223486
rect 396901 223483 396967 223486
rect 676029 223546 676095 223549
rect 676029 223544 676292 223546
rect 676029 223488 676034 223544
rect 676090 223488 676292 223544
rect 676029 223486 676292 223488
rect 676029 223483 676095 223486
rect 121361 223410 121427 223413
rect 221549 223410 221615 223413
rect 121361 223408 221615 223410
rect 121361 223352 121366 223408
rect 121422 223352 221554 223408
rect 221610 223352 221615 223408
rect 121361 223350 221615 223352
rect 121361 223347 121427 223350
rect 221549 223347 221615 223350
rect 374637 223410 374703 223413
rect 483841 223410 483907 223413
rect 374637 223408 483907 223410
rect 374637 223352 374642 223408
rect 374698 223352 483846 223408
rect 483902 223352 483907 223408
rect 374637 223350 483907 223352
rect 374637 223347 374703 223350
rect 483841 223347 483907 223350
rect 111609 223274 111675 223277
rect 217317 223274 217383 223277
rect 111609 223272 217383 223274
rect 111609 223216 111614 223272
rect 111670 223216 217322 223272
rect 217378 223216 217383 223272
rect 111609 223214 217383 223216
rect 111609 223211 111675 223214
rect 217317 223211 217383 223214
rect 377581 223274 377647 223277
rect 489453 223274 489519 223277
rect 377581 223272 489519 223274
rect 377581 223216 377586 223272
rect 377642 223216 489458 223272
rect 489514 223216 489519 223272
rect 377581 223214 489519 223216
rect 377581 223211 377647 223214
rect 489453 223211 489519 223214
rect 104801 223138 104867 223141
rect 214465 223138 214531 223141
rect 104801 223136 214531 223138
rect 104801 223080 104806 223136
rect 104862 223080 214470 223136
rect 214526 223080 214531 223136
rect 104801 223078 214531 223080
rect 104801 223075 104867 223078
rect 214465 223075 214531 223078
rect 331029 223138 331095 223141
rect 376753 223138 376819 223141
rect 331029 223136 376819 223138
rect 331029 223080 331034 223136
rect 331090 223080 376758 223136
rect 376814 223080 376819 223136
rect 331029 223078 376819 223080
rect 331029 223075 331095 223078
rect 376753 223075 376819 223078
rect 377949 223138 378015 223141
rect 488625 223138 488691 223141
rect 377949 223136 488691 223138
rect 377949 223080 377954 223136
rect 378010 223080 488630 223136
rect 488686 223080 488691 223136
rect 377949 223078 488691 223080
rect 377949 223075 378015 223078
rect 488625 223075 488691 223078
rect 675845 223138 675911 223141
rect 675845 223136 676292 223138
rect 675845 223080 675850 223136
rect 675906 223080 676292 223136
rect 675845 223078 676292 223080
rect 675845 223075 675911 223078
rect 96429 223002 96495 223005
rect 211245 223002 211311 223005
rect 96429 223000 211311 223002
rect 96429 222944 96434 223000
rect 96490 222944 211250 223000
rect 211306 222944 211311 223000
rect 96429 222942 211311 222944
rect 96429 222939 96495 222942
rect 211245 222939 211311 222942
rect 331121 223002 331187 223005
rect 377581 223002 377647 223005
rect 331121 223000 377647 223002
rect 331121 222944 331126 223000
rect 331182 222944 377586 223000
rect 377642 222944 377647 223000
rect 331121 222942 377647 222944
rect 331121 222939 331187 222942
rect 377581 222939 377647 222942
rect 380709 223002 380775 223005
rect 495341 223002 495407 223005
rect 380709 223000 495407 223002
rect 380709 222944 380714 223000
rect 380770 222944 495346 223000
rect 495402 222944 495407 223000
rect 380709 222942 495407 222944
rect 380709 222939 380775 222942
rect 495341 222939 495407 222942
rect 79593 222866 79659 222869
rect 204345 222866 204411 222869
rect 79593 222864 204411 222866
rect 79593 222808 79598 222864
rect 79654 222808 204350 222864
rect 204406 222808 204411 222864
rect 79593 222806 204411 222808
rect 79593 222803 79659 222806
rect 204345 222803 204411 222806
rect 328085 222866 328151 222869
rect 374177 222866 374243 222869
rect 328085 222864 374243 222866
rect 328085 222808 328090 222864
rect 328146 222808 374182 222864
rect 374238 222808 374243 222864
rect 328085 222806 374243 222808
rect 328085 222803 328151 222806
rect 374177 222803 374243 222806
rect 380433 222866 380499 222869
rect 494053 222866 494119 222869
rect 380433 222864 494119 222866
rect 380433 222808 380438 222864
rect 380494 222808 494058 222864
rect 494114 222808 494119 222864
rect 380433 222806 494119 222808
rect 380433 222803 380499 222806
rect 494053 222803 494119 222806
rect 72877 222730 72943 222733
rect 201677 222730 201743 222733
rect 72877 222728 201743 222730
rect 72877 222672 72882 222728
rect 72938 222672 201682 222728
rect 201738 222672 201743 222728
rect 72877 222670 201743 222672
rect 72877 222667 72943 222670
rect 201677 222667 201743 222670
rect 330753 222730 330819 222733
rect 375373 222730 375439 222733
rect 330753 222728 375439 222730
rect 330753 222672 330758 222728
rect 330814 222672 375378 222728
rect 375434 222672 375439 222728
rect 330753 222670 375439 222672
rect 330753 222667 330819 222670
rect 375373 222667 375439 222670
rect 386229 222730 386295 222733
rect 507117 222730 507183 222733
rect 386229 222728 507183 222730
rect 386229 222672 386234 222728
rect 386290 222672 507122 222728
rect 507178 222672 507183 222728
rect 386229 222670 507183 222672
rect 386229 222667 386295 222670
rect 507117 222667 507183 222670
rect 675937 222730 676003 222733
rect 675937 222728 676292 222730
rect 675937 222672 675942 222728
rect 675998 222672 676292 222728
rect 675937 222670 676292 222672
rect 675937 222667 676003 222670
rect 74441 222594 74507 222597
rect 201861 222594 201927 222597
rect 74441 222592 201927 222594
rect 74441 222536 74446 222592
rect 74502 222536 201866 222592
rect 201922 222536 201927 222592
rect 74441 222534 201927 222536
rect 74441 222531 74507 222534
rect 201861 222531 201927 222534
rect 330937 222594 331003 222597
rect 381077 222594 381143 222597
rect 330937 222592 381143 222594
rect 330937 222536 330942 222592
rect 330998 222536 381082 222592
rect 381138 222536 381143 222592
rect 330937 222534 381143 222536
rect 330937 222531 331003 222534
rect 381077 222531 381143 222534
rect 382917 222594 382983 222597
rect 502609 222594 502675 222597
rect 382917 222592 502675 222594
rect 382917 222536 382922 222592
rect 382978 222536 502614 222592
rect 502670 222536 502675 222592
rect 382917 222534 502675 222536
rect 382917 222531 382983 222534
rect 502609 222531 502675 222534
rect 572621 222594 572687 222597
rect 574369 222594 574435 222597
rect 572621 222592 574435 222594
rect 572621 222536 572626 222592
rect 572682 222536 574374 222592
rect 574430 222536 574435 222592
rect 572621 222534 574435 222536
rect 572621 222531 572687 222534
rect 574369 222531 574435 222534
rect 67817 222458 67883 222461
rect 198733 222458 198799 222461
rect 67817 222456 198799 222458
rect 67817 222400 67822 222456
rect 67878 222400 198738 222456
rect 198794 222400 198799 222456
rect 67817 222398 198799 222400
rect 67817 222395 67883 222398
rect 198733 222395 198799 222398
rect 333605 222458 333671 222461
rect 384297 222458 384363 222461
rect 333605 222456 384363 222458
rect 333605 222400 333610 222456
rect 333666 222400 384302 222456
rect 384358 222400 384363 222456
rect 333605 222398 384363 222400
rect 333605 222395 333671 222398
rect 384297 222395 384363 222398
rect 388989 222458 389055 222461
rect 510613 222458 510679 222461
rect 519721 222458 519787 222461
rect 388989 222456 510679 222458
rect 388989 222400 388994 222456
rect 389050 222400 510618 222456
rect 510674 222400 510679 222456
rect 388989 222398 510679 222400
rect 388989 222395 389055 222398
rect 510613 222395 510679 222398
rect 516090 222456 519787 222458
rect 516090 222400 519726 222456
rect 519782 222400 519787 222456
rect 516090 222398 519787 222400
rect 66161 222322 66227 222325
rect 196157 222322 196223 222325
rect 66161 222320 196223 222322
rect 66161 222264 66166 222320
rect 66222 222264 196162 222320
rect 196218 222264 196223 222320
rect 66161 222262 196223 222264
rect 66161 222259 66227 222262
rect 196157 222259 196223 222262
rect 333697 222322 333763 222325
rect 387701 222322 387767 222325
rect 333697 222320 387767 222322
rect 333697 222264 333702 222320
rect 333758 222264 387706 222320
rect 387762 222264 387767 222320
rect 333697 222262 387767 222264
rect 333697 222259 333763 222262
rect 387701 222259 387767 222262
rect 391841 222322 391907 222325
rect 516090 222322 516150 222398
rect 519721 222395 519787 222398
rect 391841 222320 516150 222322
rect 391841 222264 391846 222320
rect 391902 222264 516150 222320
rect 391841 222262 516150 222264
rect 517421 222322 517487 222325
rect 517881 222322 517947 222325
rect 528645 222322 528711 222325
rect 517421 222320 528711 222322
rect 517421 222264 517426 222320
rect 517482 222264 517886 222320
rect 517942 222264 528650 222320
rect 528706 222264 528711 222320
rect 517421 222262 528711 222264
rect 391841 222259 391907 222262
rect 517421 222259 517487 222262
rect 517881 222259 517947 222262
rect 528645 222259 528711 222262
rect 675753 222322 675819 222325
rect 675753 222320 676292 222322
rect 675753 222264 675758 222320
rect 675814 222264 676292 222320
rect 675753 222262 676292 222264
rect 675753 222259 675819 222262
rect 61101 222186 61167 222189
rect 196525 222186 196591 222189
rect 61101 222184 196591 222186
rect 61101 222128 61106 222184
rect 61162 222128 196530 222184
rect 196586 222128 196591 222184
rect 61101 222126 196591 222128
rect 61101 222123 61167 222126
rect 196525 222123 196591 222126
rect 341609 222186 341675 222189
rect 400397 222186 400463 222189
rect 341609 222184 400463 222186
rect 341609 222128 341614 222184
rect 341670 222128 400402 222184
rect 400458 222128 400463 222184
rect 341609 222126 400463 222128
rect 341609 222123 341675 222126
rect 400397 222123 400463 222126
rect 411161 222186 411227 222189
rect 569309 222186 569375 222189
rect 411161 222184 569375 222186
rect 411161 222128 411166 222184
rect 411222 222128 569314 222184
rect 569370 222128 569375 222184
rect 411161 222126 569375 222128
rect 411161 222123 411227 222126
rect 569309 222123 569375 222126
rect 569861 222186 569927 222189
rect 573541 222186 573607 222189
rect 569861 222184 573607 222186
rect 569861 222128 569866 222184
rect 569922 222128 573546 222184
rect 573602 222128 573607 222184
rect 569861 222126 573607 222128
rect 569861 222123 569927 222126
rect 573541 222123 573607 222126
rect 336181 222050 336247 222053
rect 390185 222050 390251 222053
rect 336181 222048 390251 222050
rect 336181 221992 336186 222048
rect 336242 221992 390190 222048
rect 390246 221992 390251 222048
rect 336181 221990 390251 221992
rect 336181 221987 336247 221990
rect 390185 221987 390251 221990
rect 528461 222050 528527 222053
rect 628005 222050 628071 222053
rect 528461 222048 628071 222050
rect 528461 221992 528466 222048
rect 528522 221992 628010 222048
rect 628066 221992 628071 222048
rect 528461 221990 628071 221992
rect 528461 221987 528527 221990
rect 628005 221987 628071 221990
rect 522941 221914 523007 221917
rect 627085 221914 627151 221917
rect 522941 221912 627151 221914
rect 522941 221856 522946 221912
rect 523002 221856 627090 221912
rect 627146 221856 627151 221912
rect 522941 221854 627151 221856
rect 522941 221851 523007 221854
rect 627085 221851 627151 221854
rect 675569 221914 675635 221917
rect 675569 221912 676292 221914
rect 675569 221856 675574 221912
rect 675630 221856 676292 221912
rect 675569 221854 676292 221856
rect 675569 221851 675635 221854
rect 527909 221778 527975 221781
rect 528461 221778 528527 221781
rect 527909 221776 528527 221778
rect 527909 221720 527914 221776
rect 527970 221720 528466 221776
rect 528522 221720 528527 221776
rect 527909 221718 528527 221720
rect 527909 221715 527975 221718
rect 528461 221715 528527 221718
rect 528645 221778 528711 221781
rect 626165 221778 626231 221781
rect 528645 221776 626231 221778
rect 528645 221720 528650 221776
rect 528706 221720 626170 221776
rect 626226 221720 626231 221776
rect 528645 221718 626231 221720
rect 528645 221715 528711 221718
rect 626165 221715 626231 221718
rect 510613 221642 510679 221645
rect 512453 221642 512519 221645
rect 625245 221642 625311 221645
rect 510613 221640 625311 221642
rect 510613 221584 510618 221640
rect 510674 221584 512458 221640
rect 512514 221584 625250 221640
rect 625306 221584 625311 221640
rect 510613 221582 625311 221584
rect 510613 221579 510679 221582
rect 512453 221579 512519 221582
rect 625245 221579 625311 221582
rect 502609 221506 502675 221509
rect 623405 221506 623471 221509
rect 502609 221504 623471 221506
rect 502609 221448 502614 221504
rect 502670 221448 623410 221504
rect 623466 221448 623471 221504
rect 502609 221446 623471 221448
rect 502609 221443 502675 221446
rect 623405 221443 623471 221446
rect 675753 221506 675819 221509
rect 675753 221504 676292 221506
rect 675753 221448 675758 221504
rect 675814 221448 676292 221504
rect 675753 221446 676292 221448
rect 675753 221443 675819 221446
rect 507117 221370 507183 221373
rect 624325 221370 624391 221373
rect 507117 221368 624391 221370
rect 507117 221312 507122 221368
rect 507178 221312 624330 221368
rect 624386 221312 624391 221368
rect 507117 221310 624391 221312
rect 507117 221307 507183 221310
rect 624325 221307 624391 221310
rect 488625 221234 488691 221237
rect 621473 221234 621539 221237
rect 488625 221232 621539 221234
rect 488625 221176 488630 221232
rect 488686 221176 621478 221232
rect 621534 221176 621539 221232
rect 488625 221174 621539 221176
rect 488625 221171 488691 221174
rect 621473 221171 621539 221174
rect 494053 221098 494119 221101
rect 496445 221098 496511 221101
rect 637389 221098 637455 221101
rect 494053 221096 637455 221098
rect 494053 221040 494058 221096
rect 494114 221040 496450 221096
rect 496506 221040 637394 221096
rect 637450 221040 637455 221096
rect 494053 221038 637455 221040
rect 494053 221035 494119 221038
rect 496445 221035 496511 221038
rect 637389 221035 637455 221038
rect 675753 221098 675819 221101
rect 675753 221096 676292 221098
rect 675753 221040 675758 221096
rect 675814 221040 676292 221096
rect 675753 221038 676292 221040
rect 675753 221035 675819 221038
rect 492673 220962 492739 220965
rect 636929 220962 636995 220965
rect 492673 220960 636995 220962
rect 492673 220904 492678 220960
rect 492734 220904 636934 220960
rect 636990 220904 636995 220960
rect 492673 220902 636995 220904
rect 492673 220899 492739 220902
rect 636929 220899 636995 220902
rect 675661 220690 675727 220693
rect 675661 220688 676292 220690
rect 675661 220632 675666 220688
rect 675722 220632 676292 220688
rect 675661 220630 676292 220632
rect 675661 220627 675727 220630
rect 675937 220282 676003 220285
rect 675937 220280 676292 220282
rect 675937 220224 675942 220280
rect 675998 220224 676292 220280
rect 675937 220222 676292 220224
rect 675937 220219 676003 220222
rect 676070 219948 676076 220012
rect 676140 219948 676146 220012
rect 676078 219874 676138 219948
rect 676078 219814 676292 219874
rect 676029 219466 676095 219469
rect 676029 219464 676292 219466
rect 676029 219408 676034 219464
rect 676090 219408 676292 219464
rect 676029 219406 676292 219408
rect 676029 219403 676095 219406
rect 676029 219058 676095 219061
rect 676029 219056 676292 219058
rect 676029 219000 676034 219056
rect 676090 219000 676292 219056
rect 676029 218998 676292 219000
rect 676029 218995 676095 218998
rect 675937 218650 676003 218653
rect 675937 218648 676292 218650
rect 675937 218592 675942 218648
rect 675998 218592 676292 218648
rect 675937 218590 676292 218592
rect 675937 218587 676003 218590
rect 676029 218242 676095 218245
rect 676029 218240 676292 218242
rect 676029 218184 676034 218240
rect 676090 218184 676292 218240
rect 676029 218182 676292 218184
rect 676029 218179 676095 218182
rect 676029 217834 676095 217837
rect 676029 217832 676292 217834
rect 676029 217776 676034 217832
rect 676090 217776 676292 217832
rect 676029 217774 676292 217776
rect 676029 217771 676095 217774
rect 675937 217426 676003 217429
rect 675937 217424 676292 217426
rect 675937 217368 675942 217424
rect 675998 217368 676292 217424
rect 675937 217366 676292 217368
rect 675937 217363 676003 217366
rect 675661 217018 675727 217021
rect 675661 217016 676292 217018
rect 675661 216960 675666 217016
rect 675722 216960 676292 217016
rect 675661 216958 676292 216960
rect 675661 216955 675727 216958
rect 675753 216610 675819 216613
rect 675753 216608 676292 216610
rect 675753 216552 675758 216608
rect 675814 216552 676292 216608
rect 675753 216550 676292 216552
rect 675753 216547 675819 216550
rect 579705 216202 579771 216205
rect 576380 216200 579771 216202
rect 576380 216144 579710 216200
rect 579766 216144 579771 216200
rect 576380 216142 579771 216144
rect 579705 216139 579771 216142
rect 676029 216202 676095 216205
rect 676029 216200 676292 216202
rect 676029 216144 676034 216200
rect 676090 216144 676292 216200
rect 676029 216142 676292 216144
rect 676029 216139 676095 216142
rect 675937 215794 676003 215797
rect 675937 215792 676292 215794
rect 675937 215736 675942 215792
rect 675998 215736 676292 215792
rect 675937 215734 676292 215736
rect 675937 215731 676003 215734
rect 675845 215386 675911 215389
rect 675845 215384 676292 215386
rect 675845 215328 675850 215384
rect 675906 215328 676292 215384
rect 675845 215326 676292 215328
rect 675845 215323 675911 215326
rect 41505 215114 41571 215117
rect 41462 215112 41571 215114
rect 41462 215056 41510 215112
rect 41566 215056 41571 215112
rect 41462 215051 41571 215056
rect 41462 214948 41522 215051
rect 676029 214978 676095 214981
rect 676029 214976 676292 214978
rect 676029 214920 676034 214976
rect 676090 214920 676292 214976
rect 676029 214918 676292 214920
rect 676029 214915 676095 214918
rect 41413 214706 41479 214709
rect 582281 214706 582347 214709
rect 41413 214704 41522 214706
rect 41413 214648 41418 214704
rect 41474 214648 41522 214704
rect 41413 214643 41522 214648
rect 576380 214704 582347 214706
rect 576380 214648 582286 214704
rect 582342 214648 582347 214704
rect 576380 214646 582347 214648
rect 582281 214643 582347 214646
rect 41462 214540 41522 214643
rect 676029 214570 676095 214573
rect 676029 214568 676292 214570
rect 676029 214512 676034 214568
rect 676090 214512 676292 214568
rect 676029 214510 676292 214512
rect 676029 214507 676095 214510
rect 41597 214298 41663 214301
rect 41462 214296 41663 214298
rect 41462 214240 41602 214296
rect 41658 214240 41663 214296
rect 41462 214238 41663 214240
rect 41462 214132 41522 214238
rect 41597 214235 41663 214238
rect 675937 214162 676003 214165
rect 675937 214160 676292 214162
rect 675937 214104 675942 214160
rect 675998 214104 676292 214160
rect 675937 214102 676292 214104
rect 675937 214099 676003 214102
rect 41505 213890 41571 213893
rect 41462 213888 41571 213890
rect 41462 213832 41510 213888
rect 41566 213832 41571 213888
rect 41462 213827 41571 213832
rect 41462 213724 41522 213827
rect 675937 213754 676003 213757
rect 675937 213752 676292 213754
rect 675937 213696 675942 213752
rect 675998 213696 676292 213752
rect 675937 213694 676292 213696
rect 675937 213691 676003 213694
rect 42190 213346 42196 213348
rect 41492 213286 42196 213346
rect 42190 213284 42196 213286
rect 42260 213284 42266 213348
rect 675886 213284 675892 213348
rect 675956 213346 675962 213348
rect 675956 213286 676292 213346
rect 675956 213284 675962 213286
rect 580257 213210 580323 213213
rect 576380 213208 580323 213210
rect 576380 213152 580262 213208
rect 580318 213152 580323 213208
rect 576380 213150 580323 213152
rect 580257 213147 580323 213150
rect 41505 213074 41571 213077
rect 41462 213072 41571 213074
rect 41462 213016 41510 213072
rect 41566 213016 41571 213072
rect 41462 213011 41571 213016
rect 41462 212908 41522 213011
rect 675845 212938 675911 212941
rect 675845 212936 676292 212938
rect 675845 212880 675850 212936
rect 675906 212880 676292 212936
rect 675845 212878 676292 212880
rect 675845 212875 675911 212878
rect 46933 212530 46999 212533
rect 41492 212528 46999 212530
rect 41492 212472 46938 212528
rect 46994 212472 46999 212528
rect 41492 212470 46999 212472
rect 46933 212467 46999 212470
rect 675385 212530 675451 212533
rect 675886 212530 675892 212532
rect 675385 212528 675892 212530
rect 675385 212472 675390 212528
rect 675446 212472 675892 212528
rect 675385 212470 675892 212472
rect 675385 212467 675451 212470
rect 675886 212468 675892 212470
rect 675956 212530 675962 212532
rect 675956 212470 676292 212530
rect 675956 212468 675962 212470
rect 45645 212122 45711 212125
rect 41492 212120 45711 212122
rect 41492 212064 45650 212120
rect 45706 212064 45711 212120
rect 41492 212062 45711 212064
rect 45645 212059 45711 212062
rect 675845 212122 675911 212125
rect 675845 212120 676292 212122
rect 675845 212064 675850 212120
rect 675906 212064 676292 212120
rect 675845 212062 676292 212064
rect 675845 212059 675911 212062
rect 41638 211850 41644 211852
rect 41462 211790 41644 211850
rect 41462 211684 41522 211790
rect 41638 211788 41644 211790
rect 41708 211788 41714 211852
rect 581637 211714 581703 211717
rect 576380 211712 581703 211714
rect 576380 211656 581642 211712
rect 581698 211656 581703 211712
rect 576380 211654 581703 211656
rect 581637 211651 581703 211654
rect 45461 211306 45527 211309
rect 41492 211304 45527 211306
rect 41492 211248 45466 211304
rect 45522 211248 45527 211304
rect 41492 211246 45527 211248
rect 45461 211243 45527 211246
rect 41822 210898 41828 210900
rect 41492 210838 41828 210898
rect 41822 210836 41828 210838
rect 41892 210836 41898 210900
rect 42742 210490 42748 210492
rect 41492 210430 42748 210490
rect 42742 210428 42748 210430
rect 42812 210428 42818 210492
rect 580533 210218 580599 210221
rect 576380 210216 580599 210218
rect 576380 210160 580538 210216
rect 580594 210160 580599 210216
rect 576380 210158 580599 210160
rect 580533 210155 580599 210158
rect 32998 209813 33058 210052
rect 32949 209808 33058 209813
rect 32949 209752 32954 209808
rect 33010 209752 33058 209808
rect 32949 209750 33058 209752
rect 32949 209747 33015 209750
rect 41462 209402 41522 209644
rect 599761 209538 599827 209541
rect 599761 209536 606556 209538
rect 599761 209480 599766 209536
rect 599822 209480 606556 209536
rect 599761 209478 606556 209480
rect 599761 209475 599827 209478
rect 41638 209402 41644 209404
rect 41462 209342 41644 209402
rect 41638 209340 41644 209342
rect 41708 209340 41714 209404
rect 42374 209266 42380 209268
rect 41492 209206 42380 209266
rect 42374 209204 42380 209206
rect 42444 209204 42450 209268
rect 671061 209266 671127 209269
rect 666356 209264 671127 209266
rect 666356 209208 671066 209264
rect 671122 209208 671127 209264
rect 666356 209206 671127 209208
rect 671061 209203 671127 209206
rect 42558 208858 42564 208860
rect 41492 208798 42564 208858
rect 42558 208796 42564 208798
rect 42628 208796 42634 208860
rect 581453 208722 581519 208725
rect 576380 208720 581519 208722
rect 576380 208664 581458 208720
rect 581514 208664 581519 208720
rect 576380 208662 581519 208664
rect 581453 208659 581519 208662
rect 599945 208586 600011 208589
rect 599945 208584 606556 208586
rect 599945 208528 599950 208584
rect 600006 208528 606556 208584
rect 599945 208526 606556 208528
rect 599945 208523 600011 208526
rect 32998 208181 33058 208420
rect 32998 208176 33107 208181
rect 32998 208120 33046 208176
rect 33102 208120 33107 208176
rect 32998 208118 33107 208120
rect 33041 208115 33107 208118
rect 41822 208042 41828 208044
rect 41492 207982 41828 208042
rect 41822 207980 41828 207982
rect 41892 207980 41898 208044
rect 42190 207634 42196 207636
rect 41492 207574 42196 207634
rect 42190 207572 42196 207574
rect 42260 207572 42266 207636
rect 599853 207498 599919 207501
rect 599853 207496 606556 207498
rect 599853 207440 599858 207496
rect 599914 207440 606556 207496
rect 599853 207438 606556 207440
rect 599853 207435 599919 207438
rect 42006 207226 42012 207228
rect 41492 207166 42012 207226
rect 42006 207164 42012 207166
rect 42076 207164 42082 207228
rect 582281 207090 582347 207093
rect 576380 207088 582347 207090
rect 576380 207032 582286 207088
rect 582342 207032 582347 207088
rect 576380 207030 582347 207032
rect 582281 207027 582347 207030
rect 42885 206818 42951 206821
rect 41492 206816 42951 206818
rect 41492 206760 42890 206816
rect 42946 206760 42951 206816
rect 41492 206758 42951 206760
rect 42885 206755 42951 206758
rect 600037 206546 600103 206549
rect 600037 206544 606556 206546
rect 600037 206488 600042 206544
rect 600098 206488 606556 206544
rect 600037 206486 606556 206488
rect 600037 206483 600103 206486
rect 43069 206410 43135 206413
rect 41492 206408 43135 206410
rect 41492 206352 43074 206408
rect 43130 206352 43135 206408
rect 41492 206350 43135 206352
rect 43069 206347 43135 206350
rect 41462 205732 41522 205972
rect 671061 205866 671127 205869
rect 666356 205864 671127 205866
rect 666356 205808 671066 205864
rect 671122 205808 671127 205864
rect 666356 205806 671127 205808
rect 671061 205803 671127 205806
rect 41454 205668 41460 205732
rect 41524 205668 41530 205732
rect 42977 205594 43043 205597
rect 582281 205594 582347 205597
rect 41492 205592 43043 205594
rect 41492 205536 42982 205592
rect 43038 205536 43043 205592
rect 41492 205534 43043 205536
rect 576380 205592 582347 205594
rect 576380 205536 582286 205592
rect 582342 205536 582347 205592
rect 576380 205534 582347 205536
rect 42977 205531 43043 205534
rect 582281 205531 582347 205534
rect 599117 205458 599183 205461
rect 599117 205456 606556 205458
rect 599117 205400 599122 205456
rect 599178 205400 606556 205456
rect 599117 205398 606556 205400
rect 599117 205395 599183 205398
rect 42793 205186 42859 205189
rect 41492 205184 42859 205186
rect 41492 205128 42798 205184
rect 42854 205128 42859 205184
rect 41492 205126 42859 205128
rect 42793 205123 42859 205126
rect 31845 204914 31911 204917
rect 31845 204912 31954 204914
rect 31845 204856 31850 204912
rect 31906 204856 31954 204912
rect 31845 204851 31954 204856
rect 31894 204748 31954 204851
rect 600957 204506 601023 204509
rect 600957 204504 606556 204506
rect 600957 204448 600962 204504
rect 601018 204448 606556 204504
rect 600957 204446 606556 204448
rect 600957 204443 601023 204446
rect 48221 204370 48287 204373
rect 41492 204368 48287 204370
rect 41492 204312 48226 204368
rect 48282 204312 48287 204368
rect 41492 204310 48287 204312
rect 48221 204307 48287 204310
rect 670969 204234 671035 204237
rect 666356 204232 671035 204234
rect 666356 204176 670974 204232
rect 671030 204176 671035 204232
rect 666356 204174 671035 204176
rect 670969 204171 671035 204174
rect 31661 204098 31727 204101
rect 581821 204098 581887 204101
rect 31661 204096 31770 204098
rect 31661 204040 31666 204096
rect 31722 204040 31770 204096
rect 31661 204035 31770 204040
rect 576380 204096 581887 204098
rect 576380 204040 581826 204096
rect 581882 204040 581887 204096
rect 576380 204038 581887 204040
rect 581821 204035 581887 204038
rect 31710 203932 31770 204035
rect 601141 203418 601207 203421
rect 601141 203416 606556 203418
rect 601141 203360 601146 203416
rect 601202 203360 606556 203416
rect 601141 203358 606556 203360
rect 601141 203355 601207 203358
rect 581085 202602 581151 202605
rect 576380 202600 581151 202602
rect 576380 202544 581090 202600
rect 581146 202544 581151 202600
rect 576380 202542 581151 202544
rect 581085 202539 581151 202542
rect 599945 202466 600011 202469
rect 599945 202464 606556 202466
rect 599945 202408 599950 202464
rect 600006 202408 606556 202464
rect 599945 202406 606556 202408
rect 599945 202403 600011 202406
rect 599025 201378 599091 201381
rect 599025 201376 606556 201378
rect 599025 201320 599030 201376
rect 599086 201320 606556 201376
rect 599025 201318 606556 201320
rect 599025 201315 599091 201318
rect 581085 201106 581151 201109
rect 576380 201104 581151 201106
rect 576380 201048 581090 201104
rect 581146 201048 581151 201104
rect 576380 201046 581151 201048
rect 581085 201043 581151 201046
rect 670969 200834 671035 200837
rect 666356 200832 671035 200834
rect 666356 200776 670974 200832
rect 671030 200776 671035 200832
rect 666356 200774 671035 200776
rect 670969 200771 671035 200774
rect 599945 200426 600011 200429
rect 599945 200424 606556 200426
rect 599945 200368 599950 200424
rect 600006 200368 606556 200424
rect 599945 200366 606556 200368
rect 599945 200363 600011 200366
rect 582281 199610 582347 199613
rect 576380 199608 582347 199610
rect 576380 199552 582286 199608
rect 582342 199552 582347 199608
rect 576380 199550 582347 199552
rect 582281 199547 582347 199550
rect 599945 199338 600011 199341
rect 599945 199336 606556 199338
rect 599945 199280 599950 199336
rect 600006 199280 606556 199336
rect 599945 199278 606556 199280
rect 599945 199275 600011 199278
rect 670877 199066 670943 199069
rect 666356 199064 670943 199066
rect 666356 199008 670882 199064
rect 670938 199008 670943 199064
rect 666356 199006 670943 199008
rect 670877 199003 670943 199006
rect 599117 198386 599183 198389
rect 599117 198384 606556 198386
rect 599117 198328 599122 198384
rect 599178 198328 606556 198384
rect 599117 198326 606556 198328
rect 599117 198323 599183 198326
rect 581269 197978 581335 197981
rect 576380 197976 581335 197978
rect 576380 197920 581274 197976
rect 581330 197920 581335 197976
rect 576380 197918 581335 197920
rect 581269 197915 581335 197918
rect 599301 197298 599367 197301
rect 599301 197296 606556 197298
rect 599301 197240 599306 197296
rect 599362 197240 606556 197296
rect 599301 197238 606556 197240
rect 599301 197235 599367 197238
rect 580809 196482 580875 196485
rect 576380 196480 580875 196482
rect 576380 196424 580814 196480
rect 580870 196424 580875 196480
rect 576380 196422 580875 196424
rect 580809 196419 580875 196422
rect 599945 196346 600011 196349
rect 599945 196344 606556 196346
rect 599945 196288 599950 196344
rect 600006 196288 606556 196344
rect 599945 196286 606556 196288
rect 599945 196283 600011 196286
rect 670877 195666 670943 195669
rect 666356 195664 670943 195666
rect 666356 195608 670882 195664
rect 670938 195608 670943 195664
rect 666356 195606 670943 195608
rect 670877 195603 670943 195606
rect 599945 195258 600011 195261
rect 599945 195256 606556 195258
rect 599945 195200 599950 195256
rect 600006 195200 606556 195256
rect 599945 195198 606556 195200
rect 599945 195195 600011 195198
rect 582281 194986 582347 194989
rect 576380 194984 582347 194986
rect 576380 194928 582286 194984
rect 582342 194928 582347 194984
rect 576380 194926 582347 194928
rect 582281 194923 582347 194926
rect 599117 194306 599183 194309
rect 599117 194304 606556 194306
rect 599117 194248 599122 194304
rect 599178 194248 606556 194304
rect 599117 194246 606556 194248
rect 599117 194243 599183 194246
rect 670785 194034 670851 194037
rect 666356 194032 670851 194034
rect 666356 193976 670790 194032
rect 670846 193976 670851 194032
rect 666356 193974 670851 193976
rect 670785 193971 670851 193974
rect 582189 193490 582255 193493
rect 576380 193488 582255 193490
rect 576380 193432 582194 193488
rect 582250 193432 582255 193488
rect 576380 193430 582255 193432
rect 582189 193427 582255 193430
rect 599853 193218 599919 193221
rect 599853 193216 606556 193218
rect 599853 193160 599858 193216
rect 599914 193160 606556 193216
rect 599853 193158 606556 193160
rect 599853 193155 599919 193158
rect 599945 192266 600011 192269
rect 599945 192264 606556 192266
rect 599945 192208 599950 192264
rect 600006 192208 606556 192264
rect 599945 192206 606556 192208
rect 599945 192203 600011 192206
rect 582281 191994 582347 191997
rect 576380 191992 582347 191994
rect 576380 191936 582286 191992
rect 582342 191936 582347 191992
rect 576380 191934 582347 191936
rect 582281 191931 582347 191934
rect 599853 191178 599919 191181
rect 599853 191176 606556 191178
rect 599853 191120 599858 191176
rect 599914 191120 606556 191176
rect 599853 191118 606556 191120
rect 599853 191115 599919 191118
rect 670785 190634 670851 190637
rect 666356 190632 670851 190634
rect 666356 190576 670790 190632
rect 670846 190576 670851 190632
rect 666356 190574 670851 190576
rect 670785 190571 670851 190574
rect 581269 190498 581335 190501
rect 576380 190496 581335 190498
rect 576380 190440 581274 190496
rect 581330 190440 581335 190496
rect 576380 190438 581335 190440
rect 581269 190435 581335 190438
rect 42149 190226 42215 190229
rect 42558 190226 42564 190228
rect 42149 190224 42564 190226
rect 42149 190168 42154 190224
rect 42210 190168 42564 190224
rect 42149 190166 42564 190168
rect 42149 190163 42215 190166
rect 42558 190164 42564 190166
rect 42628 190164 42634 190228
rect 600957 190226 601023 190229
rect 600957 190224 606556 190226
rect 600957 190168 600962 190224
rect 601018 190168 606556 190224
rect 600957 190166 606556 190168
rect 600957 190163 601023 190166
rect 601601 189138 601667 189141
rect 601601 189136 606556 189138
rect 601601 189080 601606 189136
rect 601662 189080 606556 189136
rect 601601 189078 606556 189080
rect 601601 189075 601667 189078
rect 670693 189002 670759 189005
rect 666356 189000 670759 189002
rect 666356 188944 670698 189000
rect 670754 188944 670759 189000
rect 666356 188942 670759 188944
rect 670693 188939 670759 188942
rect 579705 188866 579771 188869
rect 576380 188864 579771 188866
rect 576380 188808 579710 188864
rect 579766 188808 579771 188864
rect 576380 188806 579771 188808
rect 579705 188803 579771 188806
rect 601509 188186 601575 188189
rect 601509 188184 606556 188186
rect 601509 188128 601514 188184
rect 601570 188128 606556 188184
rect 601509 188126 606556 188128
rect 601509 188123 601575 188126
rect 41454 187580 41460 187644
rect 41524 187642 41530 187644
rect 41873 187642 41939 187645
rect 41524 187640 41939 187642
rect 41524 187584 41878 187640
rect 41934 187584 41939 187640
rect 41524 187582 41939 187584
rect 41524 187580 41530 187582
rect 41873 187579 41939 187582
rect 582281 187370 582347 187373
rect 576380 187368 582347 187370
rect 576380 187312 582286 187368
rect 582342 187312 582347 187368
rect 576380 187310 582347 187312
rect 582281 187307 582347 187310
rect 41965 187100 42031 187101
rect 41965 187096 42012 187100
rect 42076 187098 42082 187100
rect 599945 187098 600011 187101
rect 41965 187040 41970 187096
rect 41965 187036 42012 187040
rect 42076 187038 42122 187098
rect 599945 187096 606556 187098
rect 599945 187040 599950 187096
rect 600006 187040 606556 187096
rect 599945 187038 606556 187040
rect 42076 187036 42082 187038
rect 41965 187035 42031 187036
rect 599945 187035 600011 187038
rect 42057 186418 42123 186421
rect 42190 186418 42196 186420
rect 42057 186416 42196 186418
rect 42057 186360 42062 186416
rect 42118 186360 42196 186416
rect 42057 186358 42196 186360
rect 42057 186355 42123 186358
rect 42190 186356 42196 186358
rect 42260 186356 42266 186420
rect 600037 186146 600103 186149
rect 600037 186144 606556 186146
rect 600037 186088 600042 186144
rect 600098 186088 606556 186144
rect 600037 186086 606556 186088
rect 600037 186083 600103 186086
rect 42149 185874 42215 185877
rect 42374 185874 42380 185876
rect 42149 185872 42380 185874
rect 42149 185816 42154 185872
rect 42210 185816 42380 185872
rect 42149 185814 42380 185816
rect 42149 185811 42215 185814
rect 42374 185812 42380 185814
rect 42444 185812 42450 185876
rect 582189 185874 582255 185877
rect 576380 185872 582255 185874
rect 576380 185816 582194 185872
rect 582250 185816 582255 185872
rect 576380 185814 582255 185816
rect 582189 185811 582255 185814
rect 670693 185602 670759 185605
rect 666356 185600 670759 185602
rect 666356 185544 670698 185600
rect 670754 185544 670759 185600
rect 666356 185542 670759 185544
rect 670693 185539 670759 185542
rect 599853 185058 599919 185061
rect 599853 185056 606556 185058
rect 599853 185000 599858 185056
rect 599914 185000 606556 185056
rect 599853 184998 606556 185000
rect 599853 184995 599919 184998
rect 580901 184378 580967 184381
rect 576380 184376 580967 184378
rect 576380 184320 580906 184376
rect 580962 184320 580967 184376
rect 576380 184318 580967 184320
rect 580901 184315 580967 184318
rect 42149 184242 42215 184245
rect 42742 184242 42748 184244
rect 42149 184240 42748 184242
rect 42149 184184 42154 184240
rect 42210 184184 42748 184240
rect 42149 184182 42748 184184
rect 42149 184179 42215 184182
rect 42742 184180 42748 184182
rect 42812 184180 42818 184244
rect 599761 184106 599827 184109
rect 599761 184104 606556 184106
rect 599761 184048 599766 184104
rect 599822 184048 606556 184104
rect 599761 184046 606556 184048
rect 599761 184043 599827 184046
rect 666737 183834 666803 183837
rect 672073 183834 672139 183837
rect 666356 183832 672139 183834
rect 666356 183776 666742 183832
rect 666798 183776 672078 183832
rect 672134 183776 672139 183832
rect 666356 183774 672139 183776
rect 666737 183771 666803 183774
rect 672073 183771 672139 183774
rect 41781 183700 41847 183701
rect 41781 183696 41828 183700
rect 41892 183698 41898 183700
rect 41781 183640 41786 183696
rect 41781 183636 41828 183640
rect 41892 183638 41938 183698
rect 41892 183636 41898 183638
rect 41781 183635 41847 183636
rect 599945 183018 600011 183021
rect 599945 183016 606556 183018
rect 599945 182960 599950 183016
rect 600006 182960 606556 183016
rect 599945 182958 606556 182960
rect 599945 182955 600011 182958
rect 580257 182882 580323 182885
rect 576380 182880 580323 182882
rect 576380 182824 580262 182880
rect 580318 182824 580323 182880
rect 576380 182822 580323 182824
rect 580257 182819 580323 182822
rect 41638 182684 41644 182748
rect 41708 182746 41714 182748
rect 41781 182746 41847 182749
rect 41708 182744 41847 182746
rect 41708 182688 41786 182744
rect 41842 182688 41847 182744
rect 41708 182686 41847 182688
rect 41708 182684 41714 182686
rect 41781 182683 41847 182686
rect 599853 182066 599919 182069
rect 599853 182064 606556 182066
rect 599853 182008 599858 182064
rect 599914 182008 606556 182064
rect 599853 182006 606556 182008
rect 599853 182003 599919 182006
rect 580533 181386 580599 181389
rect 576380 181384 580599 181386
rect 576380 181328 580538 181384
rect 580594 181328 580599 181384
rect 576380 181326 580599 181328
rect 580533 181323 580599 181326
rect 600129 180978 600195 180981
rect 600129 180976 606556 180978
rect 600129 180920 600134 180976
rect 600190 180920 606556 180976
rect 600129 180918 606556 180920
rect 600129 180915 600195 180918
rect 666737 180434 666803 180437
rect 666356 180432 666803 180434
rect 666356 180376 666742 180432
rect 666798 180376 666803 180432
rect 666356 180374 666803 180376
rect 666737 180371 666803 180374
rect 600037 180026 600103 180029
rect 600037 180024 606556 180026
rect 600037 179968 600042 180024
rect 600098 179968 606556 180024
rect 600037 179966 606556 179968
rect 600037 179963 600103 179966
rect 581821 179754 581887 179757
rect 576380 179752 581887 179754
rect 576380 179696 581826 179752
rect 581882 179696 581887 179752
rect 576380 179694 581887 179696
rect 581821 179691 581887 179694
rect 703905 179346 703971 179349
rect 709057 179346 709123 179349
rect 703905 179344 709123 179346
rect 703905 179288 703910 179344
rect 703966 179288 709062 179344
rect 709118 179288 709123 179344
rect 703905 179286 709123 179288
rect 703905 179283 703971 179286
rect 709057 179283 709123 179286
rect 599669 178938 599735 178941
rect 599669 178936 606556 178938
rect 599669 178880 599674 178936
rect 599730 178880 606556 178936
rect 599669 178878 606556 178880
rect 599669 178875 599735 178878
rect 666737 178802 666803 178805
rect 672165 178802 672231 178805
rect 666356 178800 672231 178802
rect 666356 178744 666742 178800
rect 666798 178744 672170 178800
rect 672226 178744 672231 178800
rect 666356 178742 672231 178744
rect 666737 178739 666803 178742
rect 672165 178739 672231 178742
rect 675753 178530 675819 178533
rect 675753 178528 676292 178530
rect 675753 178472 675758 178528
rect 675814 178472 676292 178528
rect 675753 178470 676292 178472
rect 675753 178467 675819 178470
rect 581085 178258 581151 178261
rect 576380 178256 581151 178258
rect 576380 178200 581090 178256
rect 581146 178200 581151 178256
rect 576380 178198 581151 178200
rect 581085 178195 581151 178198
rect 675937 178122 676003 178125
rect 675937 178120 676292 178122
rect 675937 178064 675942 178120
rect 675998 178064 676292 178120
rect 675937 178062 676292 178064
rect 675937 178059 676003 178062
rect 599761 177986 599827 177989
rect 599761 177984 606556 177986
rect 599761 177928 599766 177984
rect 599822 177928 606556 177984
rect 599761 177926 606556 177928
rect 599761 177923 599827 177926
rect 676029 177714 676095 177717
rect 676029 177712 676292 177714
rect 676029 177656 676034 177712
rect 676090 177656 676292 177712
rect 676029 177654 676292 177656
rect 676029 177651 676095 177654
rect 675845 177306 675911 177309
rect 675845 177304 676292 177306
rect 675845 177248 675850 177304
rect 675906 177248 676292 177304
rect 675845 177246 676292 177248
rect 675845 177243 675911 177246
rect 598933 176898 598999 176901
rect 675937 176898 676003 176901
rect 598933 176896 606556 176898
rect 598933 176840 598938 176896
rect 598994 176840 606556 176896
rect 598933 176838 606556 176840
rect 675937 176896 676292 176898
rect 675937 176840 675942 176896
rect 675998 176840 676292 176896
rect 675937 176838 676292 176840
rect 598933 176835 598999 176838
rect 675937 176835 676003 176838
rect 580717 176762 580783 176765
rect 576380 176760 580783 176762
rect 576380 176704 580722 176760
rect 580778 176704 580783 176760
rect 576380 176702 580783 176704
rect 580717 176699 580783 176702
rect 676029 176490 676095 176493
rect 676029 176488 676292 176490
rect 676029 176432 676034 176488
rect 676090 176432 676292 176488
rect 676029 176430 676292 176432
rect 676029 176427 676095 176430
rect 675937 176082 676003 176085
rect 675937 176080 676292 176082
rect 675937 176024 675942 176080
rect 675998 176024 676292 176080
rect 675937 176022 676292 176024
rect 675937 176019 676003 176022
rect 600221 175946 600287 175949
rect 600221 175944 606556 175946
rect 600221 175888 600226 175944
rect 600282 175888 606556 175944
rect 600221 175886 606556 175888
rect 600221 175883 600287 175886
rect 676029 175674 676095 175677
rect 676029 175672 676292 175674
rect 676029 175616 676034 175672
rect 676090 175616 676292 175672
rect 676029 175614 676292 175616
rect 676029 175611 676095 175614
rect 666737 175402 666803 175405
rect 666356 175400 666803 175402
rect 666356 175344 666742 175400
rect 666798 175344 666803 175400
rect 666356 175342 666803 175344
rect 666737 175339 666803 175342
rect 581453 175266 581519 175269
rect 576380 175264 581519 175266
rect 576380 175208 581458 175264
rect 581514 175208 581519 175264
rect 576380 175206 581519 175208
rect 581453 175203 581519 175206
rect 675937 175266 676003 175269
rect 675937 175264 676292 175266
rect 675937 175208 675942 175264
rect 675998 175208 676292 175264
rect 675937 175206 676292 175208
rect 675937 175203 676003 175206
rect 599945 174858 600011 174861
rect 676029 174858 676095 174861
rect 599945 174856 606556 174858
rect 599945 174800 599950 174856
rect 600006 174800 606556 174856
rect 599945 174798 606556 174800
rect 676029 174856 676292 174858
rect 676029 174800 676034 174856
rect 676090 174800 676292 174856
rect 676029 174798 676292 174800
rect 599945 174795 600011 174798
rect 676029 174795 676095 174798
rect 676029 174450 676095 174453
rect 676029 174448 676292 174450
rect 676029 174392 676034 174448
rect 676090 174392 676292 174448
rect 676029 174390 676292 174392
rect 676029 174387 676095 174390
rect 676029 174042 676095 174045
rect 676029 174040 676292 174042
rect 676029 173984 676034 174040
rect 676090 173984 676292 174040
rect 676029 173982 676292 173984
rect 676029 173979 676095 173982
rect 601417 173906 601483 173909
rect 601417 173904 606556 173906
rect 601417 173848 601422 173904
rect 601478 173848 606556 173904
rect 601417 173846 606556 173848
rect 601417 173843 601483 173846
rect 582281 173770 582347 173773
rect 576380 173768 582347 173770
rect 576380 173712 582286 173768
rect 582342 173712 582347 173768
rect 576380 173710 582347 173712
rect 582281 173707 582347 173710
rect 666737 173634 666803 173637
rect 671797 173634 671863 173637
rect 666356 173632 671863 173634
rect 666356 173576 666742 173632
rect 666798 173576 671802 173632
rect 671858 173576 671863 173632
rect 666356 173574 671863 173576
rect 666737 173571 666803 173574
rect 671797 173571 671863 173574
rect 675886 173572 675892 173636
rect 675956 173634 675962 173636
rect 675956 173574 676292 173634
rect 675956 173572 675962 173574
rect 675753 173226 675819 173229
rect 675753 173224 676292 173226
rect 675753 173168 675758 173224
rect 675814 173168 676292 173224
rect 675753 173166 676292 173168
rect 675753 173163 675819 173166
rect 599853 172818 599919 172821
rect 676029 172818 676095 172821
rect 599853 172816 606556 172818
rect 599853 172760 599858 172816
rect 599914 172760 606556 172816
rect 599853 172758 606556 172760
rect 676029 172816 676292 172818
rect 676029 172760 676034 172816
rect 676090 172760 676292 172816
rect 676029 172758 676292 172760
rect 599853 172755 599919 172758
rect 676029 172755 676095 172758
rect 675937 172410 676003 172413
rect 675937 172408 676292 172410
rect 675937 172352 675942 172408
rect 675998 172352 676292 172408
rect 675937 172350 676292 172352
rect 675937 172347 676003 172350
rect 579705 172274 579771 172277
rect 576380 172272 579771 172274
rect 576380 172216 579710 172272
rect 579766 172216 579771 172272
rect 576380 172214 579771 172216
rect 579705 172211 579771 172214
rect 676078 171942 676292 172002
rect 599945 171866 600011 171869
rect 676078 171868 676138 171942
rect 599945 171864 606556 171866
rect 599945 171808 599950 171864
rect 600006 171808 606556 171864
rect 599945 171806 606556 171808
rect 599945 171803 600011 171806
rect 676070 171804 676076 171868
rect 676140 171804 676146 171868
rect 676029 171594 676095 171597
rect 676029 171592 676292 171594
rect 676029 171536 676034 171592
rect 676090 171536 676292 171592
rect 676029 171534 676292 171536
rect 676029 171531 676095 171534
rect 675937 171186 676003 171189
rect 675937 171184 676292 171186
rect 675937 171128 675942 171184
rect 675998 171128 676292 171184
rect 675937 171126 676292 171128
rect 675937 171123 676003 171126
rect 598933 170778 598999 170781
rect 676029 170778 676095 170781
rect 598933 170776 606556 170778
rect 598933 170720 598938 170776
rect 598994 170720 606556 170776
rect 598933 170718 606556 170720
rect 676029 170776 676292 170778
rect 676029 170720 676034 170776
rect 676090 170720 676292 170776
rect 676029 170718 676292 170720
rect 598933 170715 598999 170718
rect 676029 170715 676095 170718
rect 580901 170642 580967 170645
rect 576380 170640 580967 170642
rect 576380 170584 580906 170640
rect 580962 170584 580967 170640
rect 576380 170582 580967 170584
rect 580901 170579 580967 170582
rect 675937 170370 676003 170373
rect 675937 170368 676292 170370
rect 675937 170312 675942 170368
rect 675998 170312 676292 170368
rect 675937 170310 676292 170312
rect 675937 170307 676003 170310
rect 666737 170234 666803 170237
rect 666356 170232 666803 170234
rect 666356 170176 666742 170232
rect 666798 170176 666803 170232
rect 666356 170174 666803 170176
rect 666737 170171 666803 170174
rect 675937 169962 676003 169965
rect 675937 169960 676292 169962
rect 675937 169904 675942 169960
rect 675998 169904 676292 169960
rect 675937 169902 676292 169904
rect 675937 169899 676003 169902
rect 599945 169826 600011 169829
rect 599945 169824 606556 169826
rect 599945 169768 599950 169824
rect 600006 169768 606556 169824
rect 599945 169766 606556 169768
rect 599945 169763 600011 169766
rect 676029 169554 676095 169557
rect 676029 169552 676292 169554
rect 676029 169496 676034 169552
rect 676090 169496 676292 169552
rect 676029 169494 676292 169496
rect 676029 169491 676095 169494
rect 580073 169146 580139 169149
rect 576380 169144 580139 169146
rect 576380 169088 580078 169144
rect 580134 169088 580139 169144
rect 576380 169086 580139 169088
rect 580073 169083 580139 169086
rect 675937 169146 676003 169149
rect 675937 169144 676292 169146
rect 675937 169088 675942 169144
rect 675998 169088 676292 169144
rect 675937 169086 676292 169088
rect 675937 169083 676003 169086
rect 599485 168738 599551 168741
rect 675845 168738 675911 168741
rect 599485 168736 606556 168738
rect 599485 168680 599490 168736
rect 599546 168680 606556 168736
rect 599485 168678 606556 168680
rect 675845 168736 676292 168738
rect 675845 168680 675850 168736
rect 675906 168680 676292 168736
rect 675845 168678 676292 168680
rect 599485 168675 599551 168678
rect 675845 168675 675911 168678
rect 666737 168602 666803 168605
rect 672349 168602 672415 168605
rect 666356 168600 672415 168602
rect 666356 168544 666742 168600
rect 666798 168544 672354 168600
rect 672410 168544 672415 168600
rect 666356 168542 672415 168544
rect 666737 168539 666803 168542
rect 672349 168539 672415 168542
rect 676029 168330 676095 168333
rect 676029 168328 676292 168330
rect 676029 168272 676034 168328
rect 676090 168272 676292 168328
rect 676029 168270 676292 168272
rect 676029 168267 676095 168270
rect 676029 167922 676095 167925
rect 676029 167920 676292 167922
rect 676029 167864 676034 167920
rect 676090 167864 676292 167920
rect 676029 167862 676292 167864
rect 676029 167859 676095 167862
rect 599853 167786 599919 167789
rect 599853 167784 606556 167786
rect 599853 167728 599858 167784
rect 599914 167728 606556 167784
rect 599853 167726 606556 167728
rect 599853 167723 599919 167726
rect 581085 167650 581151 167653
rect 576380 167648 581151 167650
rect 576380 167592 581090 167648
rect 581146 167592 581151 167648
rect 576380 167590 581151 167592
rect 581085 167587 581151 167590
rect 676029 167514 676095 167517
rect 676029 167512 676292 167514
rect 676029 167456 676034 167512
rect 676090 167456 676292 167512
rect 676029 167454 676292 167456
rect 676029 167451 676095 167454
rect 600037 166698 600103 166701
rect 600037 166696 606556 166698
rect 600037 166640 600042 166696
rect 600098 166640 606556 166696
rect 600037 166638 606556 166640
rect 600037 166635 600103 166638
rect 580165 166154 580231 166157
rect 576380 166152 580231 166154
rect 576380 166096 580170 166152
rect 580226 166096 580231 166152
rect 576380 166094 580231 166096
rect 580165 166091 580231 166094
rect 599945 165746 600011 165749
rect 599945 165744 606556 165746
rect 599945 165688 599950 165744
rect 600006 165688 606556 165744
rect 599945 165686 606556 165688
rect 599945 165683 600011 165686
rect 666737 165202 666803 165205
rect 666356 165200 666803 165202
rect 666356 165144 666742 165200
rect 666798 165144 666803 165200
rect 666356 165142 666803 165144
rect 666737 165139 666803 165142
rect 580809 164658 580875 164661
rect 576380 164656 580875 164658
rect 576380 164600 580814 164656
rect 580870 164600 580875 164656
rect 576380 164598 580875 164600
rect 580809 164595 580875 164598
rect 599853 164658 599919 164661
rect 599853 164656 606556 164658
rect 599853 164600 599858 164656
rect 599914 164600 606556 164656
rect 599853 164598 606556 164600
rect 599853 164595 599919 164598
rect 599945 163706 600011 163709
rect 599945 163704 606556 163706
rect 599945 163648 599950 163704
rect 600006 163648 606556 163704
rect 599945 163646 606556 163648
rect 599945 163643 600011 163646
rect 666737 163570 666803 163573
rect 672441 163570 672507 163573
rect 666356 163568 672507 163570
rect 666356 163512 666742 163568
rect 666798 163512 672446 163568
rect 672502 163512 672507 163568
rect 666356 163510 672507 163512
rect 666737 163507 666803 163510
rect 672441 163507 672507 163510
rect 581821 163162 581887 163165
rect 576380 163160 581887 163162
rect 576380 163104 581826 163160
rect 581882 163104 581887 163160
rect 576380 163102 581887 163104
rect 581821 163099 581887 163102
rect 600037 162618 600103 162621
rect 600037 162616 606556 162618
rect 600037 162560 600042 162616
rect 600098 162560 606556 162616
rect 600037 162558 606556 162560
rect 600037 162555 600103 162558
rect 599853 161666 599919 161669
rect 599853 161664 606556 161666
rect 599853 161608 599858 161664
rect 599914 161608 606556 161664
rect 599853 161606 606556 161608
rect 599853 161603 599919 161606
rect 579889 161530 579955 161533
rect 576380 161528 579955 161530
rect 576380 161472 579894 161528
rect 579950 161472 579955 161528
rect 576380 161470 579955 161472
rect 579889 161467 579955 161470
rect 599945 160578 600011 160581
rect 599945 160576 606556 160578
rect 599945 160520 599950 160576
rect 600006 160520 606556 160576
rect 599945 160518 606556 160520
rect 599945 160515 600011 160518
rect 666737 160170 666803 160173
rect 666356 160168 666803 160170
rect 666356 160112 666742 160168
rect 666798 160112 666803 160168
rect 666356 160110 666803 160112
rect 666737 160107 666803 160110
rect 582189 160034 582255 160037
rect 576380 160032 582255 160034
rect 576380 159976 582194 160032
rect 582250 159976 582255 160032
rect 576380 159974 582255 159976
rect 582189 159971 582255 159974
rect 600037 159626 600103 159629
rect 600037 159624 606556 159626
rect 600037 159568 600042 159624
rect 600098 159568 606556 159624
rect 600037 159566 606556 159568
rect 600037 159563 600103 159566
rect 579705 158538 579771 158541
rect 576380 158536 579771 158538
rect 576380 158480 579710 158536
rect 579766 158480 579771 158536
rect 576380 158478 579771 158480
rect 579705 158475 579771 158478
rect 599853 158538 599919 158541
rect 599853 158536 606556 158538
rect 599853 158480 599858 158536
rect 599914 158480 606556 158536
rect 599853 158478 606556 158480
rect 599853 158475 599919 158478
rect 666737 158402 666803 158405
rect 672533 158402 672599 158405
rect 666356 158400 672599 158402
rect 666356 158344 666742 158400
rect 666798 158344 672538 158400
rect 672594 158344 672599 158400
rect 666356 158342 672599 158344
rect 666737 158339 666803 158342
rect 672533 158339 672599 158342
rect 599945 157586 600011 157589
rect 599945 157584 606556 157586
rect 599945 157528 599950 157584
rect 600006 157528 606556 157584
rect 599945 157526 606556 157528
rect 599945 157523 600011 157526
rect 581913 157042 581979 157045
rect 576380 157040 581979 157042
rect 576380 156984 581918 157040
rect 581974 156984 581979 157040
rect 576380 156982 581979 156984
rect 581913 156979 581979 156982
rect 599853 156498 599919 156501
rect 599853 156496 606556 156498
rect 599853 156440 599858 156496
rect 599914 156440 606556 156496
rect 599853 156438 606556 156440
rect 599853 156435 599919 156438
rect 580257 155546 580323 155549
rect 576380 155544 580323 155546
rect 576380 155488 580262 155544
rect 580318 155488 580323 155544
rect 576380 155486 580323 155488
rect 580257 155483 580323 155486
rect 599945 155546 600011 155549
rect 599945 155544 606556 155546
rect 599945 155488 599950 155544
rect 600006 155488 606556 155544
rect 599945 155486 606556 155488
rect 599945 155483 600011 155486
rect 666737 155002 666803 155005
rect 666356 155000 666803 155002
rect 666356 154944 666742 155000
rect 666798 154944 666803 155000
rect 666356 154942 666803 154944
rect 666737 154939 666803 154942
rect 600037 154458 600103 154461
rect 600037 154456 606556 154458
rect 600037 154400 600042 154456
rect 600098 154400 606556 154456
rect 600037 154398 606556 154400
rect 600037 154395 600103 154398
rect 582281 154050 582347 154053
rect 576380 154048 582347 154050
rect 576380 153992 582286 154048
rect 582342 153992 582347 154048
rect 576380 153990 582347 153992
rect 582281 153987 582347 153990
rect 599853 153506 599919 153509
rect 599853 153504 606556 153506
rect 599853 153448 599858 153504
rect 599914 153448 606556 153504
rect 599853 153446 606556 153448
rect 599853 153443 599919 153446
rect 666737 153370 666803 153373
rect 672625 153370 672691 153373
rect 666356 153368 672691 153370
rect 666356 153312 666742 153368
rect 666798 153312 672630 153368
rect 672686 153312 672691 153368
rect 666356 153310 672691 153312
rect 666737 153307 666803 153310
rect 672625 153307 672691 153310
rect 580073 152418 580139 152421
rect 576380 152416 580139 152418
rect 576380 152360 580078 152416
rect 580134 152360 580139 152416
rect 576380 152358 580139 152360
rect 580073 152355 580139 152358
rect 599945 152418 600011 152421
rect 599945 152416 606556 152418
rect 599945 152360 599950 152416
rect 600006 152360 606556 152416
rect 599945 152358 606556 152360
rect 599945 152355 600011 152358
rect 598933 151466 598999 151469
rect 598933 151464 606556 151466
rect 598933 151408 598938 151464
rect 598994 151408 606556 151464
rect 598933 151406 606556 151408
rect 598933 151403 598999 151406
rect 581545 150922 581611 150925
rect 576380 150920 581611 150922
rect 576380 150864 581550 150920
rect 581606 150864 581611 150920
rect 576380 150862 581611 150864
rect 581545 150859 581611 150862
rect 599853 150378 599919 150381
rect 599853 150376 606556 150378
rect 599853 150320 599858 150376
rect 599914 150320 606556 150376
rect 599853 150318 606556 150320
rect 599853 150315 599919 150318
rect 666737 149970 666803 149973
rect 666356 149968 666803 149970
rect 666356 149912 666742 149968
rect 666798 149912 666803 149968
rect 666356 149910 666803 149912
rect 666737 149907 666803 149910
rect 581637 149426 581703 149429
rect 576380 149424 581703 149426
rect 576380 149368 581642 149424
rect 581698 149368 581703 149424
rect 576380 149366 581703 149368
rect 581637 149363 581703 149366
rect 599945 149426 600011 149429
rect 599945 149424 606556 149426
rect 599945 149368 599950 149424
rect 600006 149368 606556 149424
rect 599945 149366 606556 149368
rect 599945 149363 600011 149366
rect 675753 148474 675819 148477
rect 675886 148474 675892 148476
rect 675753 148472 675892 148474
rect 675753 148416 675758 148472
rect 675814 148416 675892 148472
rect 675753 148414 675892 148416
rect 675753 148411 675819 148414
rect 675886 148412 675892 148414
rect 675956 148412 675962 148476
rect 599853 148338 599919 148341
rect 599853 148336 606556 148338
rect 599853 148280 599858 148336
rect 599914 148280 606556 148336
rect 599853 148278 606556 148280
rect 599853 148275 599919 148278
rect 666645 148202 666711 148205
rect 672717 148202 672783 148205
rect 666356 148200 672783 148202
rect 666356 148144 666650 148200
rect 666706 148144 672722 148200
rect 672778 148144 672783 148200
rect 666356 148142 672783 148144
rect 666645 148139 666711 148142
rect 672717 148139 672783 148142
rect 581085 147930 581151 147933
rect 576380 147928 581151 147930
rect 576380 147872 581090 147928
rect 581146 147872 581151 147928
rect 576380 147870 581151 147872
rect 581085 147867 581151 147870
rect 599945 147386 600011 147389
rect 599945 147384 606556 147386
rect 599945 147328 599950 147384
rect 600006 147328 606556 147384
rect 599945 147326 606556 147328
rect 599945 147323 600011 147326
rect 581729 146434 581795 146437
rect 576380 146432 581795 146434
rect 576380 146376 581734 146432
rect 581790 146376 581795 146432
rect 576380 146374 581795 146376
rect 581729 146371 581795 146374
rect 599577 146298 599643 146301
rect 675753 146298 675819 146301
rect 676070 146298 676076 146300
rect 599577 146296 606556 146298
rect 599577 146240 599582 146296
rect 599638 146240 606556 146296
rect 599577 146238 606556 146240
rect 675753 146296 676076 146298
rect 675753 146240 675758 146296
rect 675814 146240 676076 146296
rect 675753 146238 676076 146240
rect 599577 146235 599643 146238
rect 675753 146235 675819 146238
rect 676070 146236 676076 146238
rect 676140 146236 676146 146300
rect 599945 145346 600011 145349
rect 599945 145344 606556 145346
rect 599945 145288 599950 145344
rect 600006 145288 606556 145344
rect 599945 145286 606556 145288
rect 599945 145283 600011 145286
rect 581177 144938 581243 144941
rect 666645 144938 666711 144941
rect 576380 144936 581243 144938
rect 576380 144880 581182 144936
rect 581238 144880 581243 144936
rect 576380 144878 581243 144880
rect 666356 144936 666711 144938
rect 666356 144880 666650 144936
rect 666706 144880 666711 144936
rect 666356 144878 666711 144880
rect 581177 144875 581243 144878
rect 666645 144875 666711 144878
rect 599669 144258 599735 144261
rect 599669 144256 606556 144258
rect 599669 144200 599674 144256
rect 599730 144200 606556 144256
rect 599669 144198 606556 144200
rect 599669 144195 599735 144198
rect 580717 143306 580783 143309
rect 576380 143304 580783 143306
rect 576380 143248 580722 143304
rect 580778 143248 580783 143304
rect 576380 143246 580783 143248
rect 580717 143243 580783 143246
rect 599853 143306 599919 143309
rect 599853 143304 606556 143306
rect 599853 143248 599858 143304
rect 599914 143248 606556 143304
rect 599853 143246 606556 143248
rect 599853 143243 599919 143246
rect 666645 143170 666711 143173
rect 672901 143170 672967 143173
rect 666356 143168 672967 143170
rect 666356 143112 666650 143168
rect 666706 143112 672906 143168
rect 672962 143112 672967 143168
rect 666356 143110 672967 143112
rect 666645 143107 666711 143110
rect 672901 143107 672967 143110
rect 599945 142218 600011 142221
rect 599945 142216 606556 142218
rect 599945 142160 599950 142216
rect 600006 142160 606556 142216
rect 599945 142158 606556 142160
rect 599945 142155 600011 142158
rect 580993 141810 581059 141813
rect 576380 141808 581059 141810
rect 576380 141752 580998 141808
rect 581054 141752 581059 141808
rect 576380 141750 581059 141752
rect 580993 141747 581059 141750
rect 599301 141266 599367 141269
rect 599301 141264 606556 141266
rect 599301 141208 599306 141264
rect 599362 141208 606556 141264
rect 599301 141206 606556 141208
rect 599301 141203 599367 141206
rect 582005 140314 582071 140317
rect 576380 140312 582071 140314
rect 576380 140256 582010 140312
rect 582066 140256 582071 140312
rect 576380 140254 582071 140256
rect 582005 140251 582071 140254
rect 600037 140178 600103 140181
rect 600037 140176 606556 140178
rect 600037 140120 600042 140176
rect 600098 140120 606556 140176
rect 600037 140118 606556 140120
rect 600037 140115 600103 140118
rect 666645 139770 666711 139773
rect 666356 139768 666711 139770
rect 666356 139712 666650 139768
rect 666706 139712 666711 139768
rect 666356 139710 666711 139712
rect 666645 139707 666711 139710
rect 599853 139226 599919 139229
rect 599853 139224 606556 139226
rect 599853 139168 599858 139224
rect 599914 139168 606556 139224
rect 599853 139166 606556 139168
rect 599853 139163 599919 139166
rect 580625 138818 580691 138821
rect 576380 138816 580691 138818
rect 576380 138760 580630 138816
rect 580686 138760 580691 138816
rect 576380 138758 580691 138760
rect 580625 138755 580691 138758
rect 599945 138138 600011 138141
rect 670693 138138 670759 138141
rect 672993 138138 673059 138141
rect 599945 138136 606556 138138
rect 599945 138080 599950 138136
rect 600006 138080 606556 138136
rect 599945 138078 606556 138080
rect 666356 138136 673059 138138
rect 666356 138080 670698 138136
rect 670754 138080 672998 138136
rect 673054 138080 673059 138136
rect 666356 138078 673059 138080
rect 599945 138075 600011 138078
rect 670693 138075 670759 138078
rect 672993 138075 673059 138078
rect 580901 137322 580967 137325
rect 576380 137320 580967 137322
rect 576380 137264 580906 137320
rect 580962 137264 580967 137320
rect 576380 137262 580967 137264
rect 580901 137259 580967 137262
rect 599853 137186 599919 137189
rect 599853 137184 606556 137186
rect 599853 137128 599858 137184
rect 599914 137128 606556 137184
rect 599853 137126 606556 137128
rect 599853 137123 599919 137126
rect 599945 136098 600011 136101
rect 599945 136096 606556 136098
rect 599945 136040 599950 136096
rect 600006 136040 606556 136096
rect 599945 136038 606556 136040
rect 599945 136035 600011 136038
rect 582097 135826 582163 135829
rect 576380 135824 582163 135826
rect 576380 135768 582102 135824
rect 582158 135768 582163 135824
rect 576380 135766 582163 135768
rect 582097 135763 582163 135766
rect 599853 135146 599919 135149
rect 599853 135144 606556 135146
rect 599853 135088 599858 135144
rect 599914 135088 606556 135144
rect 599853 135086 606556 135088
rect 599853 135083 599919 135086
rect 670693 134738 670759 134741
rect 666356 134736 670759 134738
rect 666356 134680 670698 134736
rect 670754 134680 670759 134736
rect 666356 134678 670759 134680
rect 670693 134675 670759 134678
rect 580809 134194 580875 134197
rect 576380 134192 580875 134194
rect 576380 134136 580814 134192
rect 580870 134136 580875 134192
rect 576380 134134 580875 134136
rect 580809 134131 580875 134134
rect 703813 134194 703879 134197
rect 709057 134194 709123 134197
rect 703813 134192 709123 134194
rect 703813 134136 703818 134192
rect 703874 134136 709062 134192
rect 709118 134136 709123 134192
rect 703813 134134 709123 134136
rect 703813 134131 703879 134134
rect 709057 134131 709123 134134
rect 599945 134058 600011 134061
rect 599945 134056 606556 134058
rect 599945 134000 599950 134056
rect 600006 134000 606556 134056
rect 599945 133998 606556 134000
rect 599945 133995 600011 133998
rect 599301 133106 599367 133109
rect 676121 133106 676187 133109
rect 676262 133106 676322 133348
rect 599301 133104 606556 133106
rect 599301 133048 599306 133104
rect 599362 133048 606556 133104
rect 599301 133046 606556 133048
rect 676121 133104 676322 133106
rect 676121 133048 676126 133104
rect 676182 133048 676322 133104
rect 676121 133046 676322 133048
rect 599301 133043 599367 133046
rect 676121 133043 676187 133046
rect 666645 132970 666711 132973
rect 673085 132970 673151 132973
rect 666356 132968 673151 132970
rect 666356 132912 666650 132968
rect 666706 132912 673090 132968
rect 673146 132912 673151 132968
rect 666356 132910 673151 132912
rect 666645 132907 666711 132910
rect 673085 132907 673151 132910
rect 676029 132970 676095 132973
rect 676029 132968 676292 132970
rect 676029 132912 676034 132968
rect 676090 132912 676292 132968
rect 676029 132910 676292 132912
rect 676029 132907 676095 132910
rect 582189 132698 582255 132701
rect 576380 132696 582255 132698
rect 576380 132640 582194 132696
rect 582250 132640 582255 132696
rect 576380 132638 582255 132640
rect 582189 132635 582255 132638
rect 676213 132698 676279 132701
rect 676213 132696 676322 132698
rect 676213 132640 676218 132696
rect 676274 132640 676322 132696
rect 676213 132635 676322 132640
rect 676262 132532 676322 132635
rect 676213 132290 676279 132293
rect 676213 132288 676322 132290
rect 676213 132232 676218 132288
rect 676274 132232 676322 132288
rect 676213 132227 676322 132232
rect 676262 132124 676322 132227
rect 598933 132018 598999 132021
rect 598933 132016 606556 132018
rect 598933 131960 598938 132016
rect 598994 131960 606556 132016
rect 598933 131958 606556 131960
rect 598933 131955 598999 131958
rect 676029 131746 676095 131749
rect 676029 131744 676292 131746
rect 676029 131688 676034 131744
rect 676090 131688 676292 131744
rect 676029 131686 676292 131688
rect 676029 131683 676095 131686
rect 676213 131474 676279 131477
rect 676213 131472 676322 131474
rect 676213 131416 676218 131472
rect 676274 131416 676322 131472
rect 676213 131411 676322 131416
rect 676262 131308 676322 131411
rect 581913 131202 581979 131205
rect 576380 131200 581979 131202
rect 576380 131144 581918 131200
rect 581974 131144 581979 131200
rect 576380 131142 581979 131144
rect 581913 131139 581979 131142
rect 599853 131066 599919 131069
rect 599853 131064 606556 131066
rect 599853 131008 599858 131064
rect 599914 131008 606556 131064
rect 599853 131006 606556 131008
rect 599853 131003 599919 131006
rect 676029 130930 676095 130933
rect 676029 130928 676292 130930
rect 676029 130872 676034 130928
rect 676090 130872 676292 130928
rect 676029 130870 676292 130872
rect 676029 130867 676095 130870
rect 676213 130658 676279 130661
rect 676213 130656 676322 130658
rect 676213 130600 676218 130656
rect 676274 130600 676322 130656
rect 676213 130595 676322 130600
rect 676262 130492 676322 130595
rect 676029 130114 676095 130117
rect 676029 130112 676292 130114
rect 676029 130056 676034 130112
rect 676090 130056 676292 130112
rect 676029 130054 676292 130056
rect 676029 130051 676095 130054
rect 599945 129978 600011 129981
rect 599945 129976 606556 129978
rect 599945 129920 599950 129976
rect 600006 129920 606556 129976
rect 599945 129918 606556 129920
rect 599945 129915 600011 129918
rect 581821 129706 581887 129709
rect 576380 129704 581887 129706
rect 576380 129648 581826 129704
rect 581882 129648 581887 129704
rect 576380 129646 581887 129648
rect 581821 129643 581887 129646
rect 676029 129706 676095 129709
rect 676029 129704 676292 129706
rect 676029 129648 676034 129704
rect 676090 129648 676292 129704
rect 676029 129646 676292 129648
rect 676029 129643 676095 129646
rect 666645 129570 666711 129573
rect 666356 129568 666711 129570
rect 666356 129512 666650 129568
rect 666706 129512 666711 129568
rect 666356 129510 666711 129512
rect 666645 129507 666711 129510
rect 676213 129434 676279 129437
rect 676213 129432 676322 129434
rect 676213 129376 676218 129432
rect 676274 129376 676322 129432
rect 676213 129371 676322 129376
rect 676262 129268 676322 129371
rect 599853 129026 599919 129029
rect 599853 129024 606556 129026
rect 599853 128968 599858 129024
rect 599914 128968 606556 129024
rect 599853 128966 606556 128968
rect 599853 128963 599919 128966
rect 676029 128890 676095 128893
rect 676029 128888 676292 128890
rect 676029 128832 676034 128888
rect 676090 128832 676292 128888
rect 676029 128830 676292 128832
rect 676029 128827 676095 128830
rect 582281 128210 582347 128213
rect 576380 128208 582347 128210
rect 576380 128152 582286 128208
rect 582342 128152 582347 128208
rect 576380 128150 582347 128152
rect 582281 128147 582347 128150
rect 676070 128148 676076 128212
rect 676140 128210 676146 128212
rect 676262 128210 676322 128452
rect 676140 128150 676322 128210
rect 676140 128148 676146 128150
rect 675753 128074 675819 128077
rect 675753 128072 676292 128074
rect 675753 128016 675758 128072
rect 675814 128016 676292 128072
rect 675753 128014 676292 128016
rect 675753 128011 675819 128014
rect 599945 127938 600011 127941
rect 666645 127938 666711 127941
rect 672809 127938 672875 127941
rect 599945 127936 606556 127938
rect 599945 127880 599950 127936
rect 600006 127880 606556 127936
rect 599945 127878 606556 127880
rect 666356 127936 672875 127938
rect 666356 127880 666650 127936
rect 666706 127880 672814 127936
rect 672870 127880 672875 127936
rect 666356 127878 672875 127880
rect 599945 127875 600011 127878
rect 666645 127875 666711 127878
rect 672809 127875 672875 127878
rect 676029 127666 676095 127669
rect 676029 127664 676292 127666
rect 676029 127608 676034 127664
rect 676090 127608 676292 127664
rect 676029 127606 676292 127608
rect 676029 127603 676095 127606
rect 675937 127258 676003 127261
rect 675937 127256 676292 127258
rect 675937 127200 675942 127256
rect 675998 127200 676292 127256
rect 675937 127198 676292 127200
rect 675937 127195 676003 127198
rect 600037 126986 600103 126989
rect 600037 126984 606556 126986
rect 600037 126928 600042 126984
rect 600098 126928 606556 126984
rect 600037 126926 606556 126928
rect 600037 126923 600103 126926
rect 675886 126788 675892 126852
rect 675956 126850 675962 126852
rect 675956 126790 676292 126850
rect 675956 126788 675962 126790
rect 581637 126714 581703 126717
rect 576380 126712 581703 126714
rect 576380 126656 581642 126712
rect 581698 126656 581703 126712
rect 576380 126654 581703 126656
rect 581637 126651 581703 126654
rect 676029 126442 676095 126445
rect 676029 126440 676292 126442
rect 676029 126384 676034 126440
rect 676090 126384 676292 126440
rect 676029 126382 676292 126384
rect 676029 126379 676095 126382
rect 675937 126034 676003 126037
rect 675937 126032 676292 126034
rect 675937 125976 675942 126032
rect 675998 125976 676292 126032
rect 675937 125974 676292 125976
rect 675937 125971 676003 125974
rect 599853 125898 599919 125901
rect 599853 125896 606556 125898
rect 599853 125840 599858 125896
rect 599914 125840 606556 125896
rect 599853 125838 606556 125840
rect 599853 125835 599919 125838
rect 676121 125354 676187 125357
rect 676262 125354 676322 125596
rect 676121 125352 676322 125354
rect 676121 125296 676126 125352
rect 676182 125296 676322 125352
rect 676121 125294 676322 125296
rect 676121 125291 676187 125294
rect 675845 125218 675911 125221
rect 675845 125216 676292 125218
rect 675845 125160 675850 125216
rect 675906 125160 676292 125216
rect 675845 125158 676292 125160
rect 675845 125155 675911 125158
rect 581453 125082 581519 125085
rect 576380 125080 581519 125082
rect 576380 125024 581458 125080
rect 581514 125024 581519 125080
rect 576380 125022 581519 125024
rect 581453 125019 581519 125022
rect 599945 124946 600011 124949
rect 599945 124944 606556 124946
rect 599945 124888 599950 124944
rect 600006 124888 606556 124944
rect 599945 124886 606556 124888
rect 599945 124883 600011 124886
rect 675845 124810 675911 124813
rect 675845 124808 676292 124810
rect 675845 124752 675850 124808
rect 675906 124752 676292 124808
rect 675845 124750 676292 124752
rect 675845 124747 675911 124750
rect 666645 124538 666711 124541
rect 666356 124536 666711 124538
rect 666356 124480 666650 124536
rect 666706 124480 666711 124536
rect 666356 124478 666711 124480
rect 666645 124475 666711 124478
rect 675937 124402 676003 124405
rect 675937 124400 676292 124402
rect 675937 124344 675942 124400
rect 675998 124344 676292 124400
rect 675937 124342 676292 124344
rect 675937 124339 676003 124342
rect 676029 123994 676095 123997
rect 676029 123992 676292 123994
rect 676029 123936 676034 123992
rect 676090 123936 676292 123992
rect 676029 123934 676292 123936
rect 676029 123931 676095 123934
rect 598933 123858 598999 123861
rect 598933 123856 606556 123858
rect 598933 123800 598938 123856
rect 598994 123800 606556 123856
rect 598933 123798 606556 123800
rect 598933 123795 598999 123798
rect 581269 123586 581335 123589
rect 576380 123584 581335 123586
rect 576380 123528 581274 123584
rect 581330 123528 581335 123584
rect 576380 123526 581335 123528
rect 581269 123523 581335 123526
rect 675937 123586 676003 123589
rect 675937 123584 676292 123586
rect 675937 123528 675942 123584
rect 675998 123528 676292 123584
rect 675937 123526 676292 123528
rect 675937 123523 676003 123526
rect 676029 123178 676095 123181
rect 676029 123176 676292 123178
rect 676029 123120 676034 123176
rect 676090 123120 676292 123176
rect 676029 123118 676292 123120
rect 676029 123115 676095 123118
rect 599853 122906 599919 122909
rect 666645 122906 666711 122909
rect 673177 122906 673243 122909
rect 599853 122904 606556 122906
rect 599853 122848 599858 122904
rect 599914 122848 606556 122904
rect 599853 122846 606556 122848
rect 666356 122904 673243 122906
rect 666356 122848 666650 122904
rect 666706 122848 673182 122904
rect 673238 122848 673243 122904
rect 666356 122846 673243 122848
rect 599853 122843 599919 122846
rect 666645 122843 666711 122846
rect 673177 122843 673243 122846
rect 676029 122770 676095 122773
rect 676029 122768 676292 122770
rect 676029 122712 676034 122768
rect 676090 122712 676292 122768
rect 676029 122710 676292 122712
rect 676029 122707 676095 122710
rect 676029 122362 676095 122365
rect 676029 122360 676292 122362
rect 676029 122304 676034 122360
rect 676090 122304 676292 122360
rect 676029 122302 676292 122304
rect 676029 122299 676095 122302
rect 579705 122090 579771 122093
rect 576380 122088 579771 122090
rect 576380 122032 579710 122088
rect 579766 122032 579771 122088
rect 576380 122030 579771 122032
rect 579705 122027 579771 122030
rect 599945 121818 600011 121821
rect 599945 121816 606556 121818
rect 599945 121760 599950 121816
rect 600006 121760 606556 121816
rect 599945 121758 606556 121760
rect 599945 121755 600011 121758
rect 600037 120866 600103 120869
rect 600037 120864 606556 120866
rect 600037 120808 600042 120864
rect 600098 120808 606556 120864
rect 600037 120806 606556 120808
rect 600037 120803 600103 120806
rect 581729 120594 581795 120597
rect 576380 120592 581795 120594
rect 576380 120536 581734 120592
rect 581790 120536 581795 120592
rect 576380 120534 581795 120536
rect 581729 120531 581795 120534
rect 599853 119778 599919 119781
rect 599853 119776 606556 119778
rect 599853 119720 599858 119776
rect 599914 119720 606556 119776
rect 599853 119718 606556 119720
rect 599853 119715 599919 119718
rect 666645 119506 666711 119509
rect 666356 119504 666711 119506
rect 666356 119448 666650 119504
rect 666706 119448 666711 119504
rect 666356 119446 666711 119448
rect 666645 119443 666711 119446
rect 579797 119098 579863 119101
rect 576380 119096 579863 119098
rect 576380 119040 579802 119096
rect 579858 119040 579863 119096
rect 576380 119038 579863 119040
rect 579797 119035 579863 119038
rect 599945 118826 600011 118829
rect 599945 118824 606556 118826
rect 599945 118768 599950 118824
rect 600006 118768 606556 118824
rect 599945 118766 606556 118768
rect 599945 118763 600011 118766
rect 599853 117738 599919 117741
rect 672349 117738 672415 117741
rect 599853 117736 606556 117738
rect 599853 117680 599858 117736
rect 599914 117680 606556 117736
rect 599853 117678 606556 117680
rect 666356 117736 672415 117738
rect 666356 117680 672354 117736
rect 672410 117680 672415 117736
rect 666356 117678 672415 117680
rect 599853 117675 599919 117678
rect 672349 117675 672415 117678
rect 581545 117602 581611 117605
rect 576380 117600 581611 117602
rect 576380 117544 581550 117600
rect 581606 117544 581611 117600
rect 576380 117542 581611 117544
rect 581545 117539 581611 117542
rect 599945 116786 600011 116789
rect 599945 116784 606556 116786
rect 599945 116728 599950 116784
rect 600006 116728 606556 116784
rect 599945 116726 606556 116728
rect 599945 116723 600011 116726
rect 672165 116106 672231 116109
rect 666356 116104 672231 116106
rect 666356 116048 672170 116104
rect 672226 116048 672231 116104
rect 666356 116046 672231 116048
rect 672165 116043 672231 116046
rect 581361 115970 581427 115973
rect 576380 115968 581427 115970
rect 576380 115912 581366 115968
rect 581422 115912 581427 115968
rect 576380 115910 581427 115912
rect 581361 115907 581427 115910
rect 599853 115698 599919 115701
rect 599853 115696 606556 115698
rect 599853 115640 599858 115696
rect 599914 115640 606556 115696
rect 599853 115638 606556 115640
rect 599853 115635 599919 115638
rect 599945 114746 600011 114749
rect 599945 114744 606556 114746
rect 599945 114688 599950 114744
rect 600006 114688 606556 114744
rect 599945 114686 606556 114688
rect 599945 114683 600011 114686
rect 581177 114474 581243 114477
rect 576380 114472 581243 114474
rect 576380 114416 581182 114472
rect 581238 114416 581243 114472
rect 576380 114414 581243 114416
rect 581177 114411 581243 114414
rect 672073 114338 672139 114341
rect 666356 114336 672139 114338
rect 666356 114280 672078 114336
rect 672134 114280 672139 114336
rect 666356 114278 672139 114280
rect 672073 114275 672139 114278
rect 593370 113598 606556 113658
rect 580942 113188 580948 113252
rect 581012 113250 581018 113252
rect 593370 113250 593430 113598
rect 581012 113190 593430 113250
rect 581012 113188 581018 113190
rect 579889 112978 579955 112981
rect 576380 112976 579955 112978
rect 576380 112920 579894 112976
rect 579950 112920 579955 112976
rect 576380 112918 579955 112920
rect 579889 112915 579955 112918
rect 599945 112706 600011 112709
rect 671429 112706 671495 112709
rect 599945 112704 606556 112706
rect 599945 112648 599950 112704
rect 600006 112648 606556 112704
rect 599945 112646 606556 112648
rect 666356 112704 671495 112706
rect 666356 112648 671434 112704
rect 671490 112648 671495 112704
rect 666356 112646 671495 112648
rect 599945 112643 600011 112646
rect 671429 112643 671495 112646
rect 599761 111618 599827 111621
rect 599761 111616 606556 111618
rect 599761 111560 599766 111616
rect 599822 111560 606556 111616
rect 599761 111558 606556 111560
rect 599761 111555 599827 111558
rect 580993 111482 581059 111485
rect 576380 111480 581059 111482
rect 576380 111424 580998 111480
rect 581054 111424 581059 111480
rect 576380 111422 581059 111424
rect 580993 111419 581059 111422
rect 672901 110938 672967 110941
rect 666356 110936 672967 110938
rect 666356 110880 672906 110936
rect 672962 110880 672967 110936
rect 666356 110878 672967 110880
rect 672901 110875 672967 110878
rect 600221 110666 600287 110669
rect 600221 110664 606556 110666
rect 600221 110608 600226 110664
rect 600282 110608 606556 110664
rect 600221 110606 606556 110608
rect 600221 110603 600287 110606
rect 581085 109986 581151 109989
rect 576380 109984 581151 109986
rect 576380 109928 581090 109984
rect 581146 109928 581151 109984
rect 576380 109926 581151 109928
rect 581085 109923 581151 109926
rect 599945 109578 600011 109581
rect 599945 109576 606556 109578
rect 599945 109520 599950 109576
rect 600006 109520 606556 109576
rect 599945 109518 606556 109520
rect 599945 109515 600011 109518
rect 672257 109306 672323 109309
rect 666356 109304 672323 109306
rect 666356 109248 672262 109304
rect 672318 109248 672323 109304
rect 666356 109246 672323 109248
rect 672257 109243 672323 109246
rect 600313 108626 600379 108629
rect 600313 108624 606556 108626
rect 600313 108568 600318 108624
rect 600374 108568 606556 108624
rect 600313 108566 606556 108568
rect 600313 108563 600379 108566
rect 580073 108490 580139 108493
rect 576380 108488 580139 108490
rect 576380 108432 580078 108488
rect 580134 108432 580139 108488
rect 576380 108430 580139 108432
rect 580073 108427 580139 108430
rect 599945 107538 600011 107541
rect 671153 107538 671219 107541
rect 599945 107536 606556 107538
rect 599945 107480 599950 107536
rect 600006 107480 606556 107536
rect 599945 107478 606556 107480
rect 666356 107536 671219 107538
rect 666356 107480 671158 107536
rect 671214 107480 671219 107536
rect 666356 107478 671219 107480
rect 599945 107475 600011 107478
rect 671153 107475 671219 107478
rect 580165 106858 580231 106861
rect 576380 106856 580231 106858
rect 576380 106800 580170 106856
rect 580226 106800 580231 106856
rect 576380 106798 580231 106800
rect 580165 106795 580231 106798
rect 600405 106586 600471 106589
rect 600405 106584 606556 106586
rect 600405 106528 600410 106584
rect 600466 106528 606556 106584
rect 600405 106526 606556 106528
rect 600405 106523 600471 106526
rect 672441 105906 672507 105909
rect 666356 105904 672507 105906
rect 666356 105848 672446 105904
rect 672502 105848 672507 105904
rect 666356 105846 672507 105848
rect 672441 105843 672507 105846
rect 600589 105498 600655 105501
rect 600589 105496 606556 105498
rect 600589 105440 600594 105496
rect 600650 105440 606556 105496
rect 600589 105438 606556 105440
rect 600589 105435 600655 105438
rect 579981 105362 580047 105365
rect 576380 105360 580047 105362
rect 576380 105304 579986 105360
rect 580042 105304 580047 105360
rect 576380 105302 580047 105304
rect 579981 105299 580047 105302
rect 600681 104546 600747 104549
rect 600681 104544 606556 104546
rect 600681 104488 600686 104544
rect 600742 104488 606556 104544
rect 600681 104486 606556 104488
rect 600681 104483 600747 104486
rect 670785 104138 670851 104141
rect 666356 104136 670851 104138
rect 666356 104080 670790 104136
rect 670846 104080 670851 104136
rect 666356 104078 670851 104080
rect 670785 104075 670851 104078
rect 580257 103866 580323 103869
rect 576380 103864 580323 103866
rect 576380 103808 580262 103864
rect 580318 103808 580323 103864
rect 576380 103806 580323 103808
rect 580257 103803 580323 103806
rect 600497 103458 600563 103461
rect 600497 103456 606556 103458
rect 600497 103400 600502 103456
rect 600558 103400 606556 103456
rect 600497 103398 606556 103400
rect 600497 103395 600563 103398
rect 675753 103322 675819 103325
rect 676070 103322 676076 103324
rect 675753 103320 676076 103322
rect 675753 103264 675758 103320
rect 675814 103264 676076 103320
rect 675753 103262 676076 103264
rect 675753 103259 675819 103262
rect 676070 103260 676076 103262
rect 676140 103260 676146 103324
rect 600865 102506 600931 102509
rect 671981 102506 672047 102509
rect 600865 102504 606556 102506
rect 600865 102448 600870 102504
rect 600926 102448 606556 102504
rect 600865 102446 606556 102448
rect 666356 102504 672047 102506
rect 666356 102448 671986 102504
rect 672042 102448 672047 102504
rect 666356 102446 672047 102448
rect 600865 102443 600931 102446
rect 671981 102443 672047 102446
rect 580901 102370 580967 102373
rect 576380 102368 580967 102370
rect 576380 102312 580906 102368
rect 580962 102312 580967 102368
rect 576380 102310 580967 102312
rect 580901 102307 580967 102310
rect 600773 101418 600839 101421
rect 675753 101418 675819 101421
rect 675886 101418 675892 101420
rect 600773 101416 606556 101418
rect 600773 101360 600778 101416
rect 600834 101360 606556 101416
rect 600773 101358 606556 101360
rect 675753 101416 675892 101418
rect 675753 101360 675758 101416
rect 675814 101360 675892 101416
rect 675753 101358 675892 101360
rect 600773 101355 600839 101358
rect 675753 101355 675819 101358
rect 675886 101356 675892 101358
rect 675956 101356 675962 101420
rect 580441 100874 580507 100877
rect 670877 100874 670943 100877
rect 576380 100872 580507 100874
rect 576380 100816 580446 100872
rect 580502 100816 580507 100872
rect 576380 100814 580507 100816
rect 666356 100872 670943 100874
rect 666356 100816 670882 100872
rect 670938 100816 670943 100872
rect 666356 100814 670943 100816
rect 580441 100811 580507 100814
rect 670877 100811 670943 100814
rect 599945 100466 600011 100469
rect 599945 100464 606556 100466
rect 599945 100408 599950 100464
rect 600006 100408 606556 100464
rect 599945 100406 606556 100408
rect 599945 100403 600011 100406
rect 580533 99378 580599 99381
rect 576380 99376 580599 99378
rect 576380 99320 580538 99376
rect 580594 99320 580599 99376
rect 576380 99318 580599 99320
rect 580533 99315 580599 99318
rect 580349 97746 580415 97749
rect 576380 97744 580415 97746
rect 576380 97688 580354 97744
rect 580410 97688 580415 97744
rect 576380 97686 580415 97688
rect 580349 97683 580415 97686
rect 580717 96250 580783 96253
rect 576380 96248 580783 96250
rect 576380 96192 580722 96248
rect 580778 96192 580783 96248
rect 576380 96190 580783 96192
rect 580717 96187 580783 96190
rect 628281 95978 628347 95981
rect 628238 95976 628347 95978
rect 628238 95920 628286 95976
rect 628342 95920 628347 95976
rect 628238 95915 628347 95920
rect 628238 95404 628298 95915
rect 640517 95706 640583 95709
rect 640517 95704 642466 95706
rect 640517 95648 640522 95704
rect 640578 95648 642466 95704
rect 640517 95646 642466 95648
rect 640517 95643 640583 95646
rect 582189 94754 582255 94757
rect 576380 94752 582255 94754
rect 576380 94696 582194 94752
rect 582250 94696 582255 94752
rect 576380 94694 582255 94696
rect 582189 94691 582255 94694
rect 642406 94588 642466 95646
rect 662086 95508 662092 95572
rect 662156 95570 662162 95572
rect 662229 95570 662295 95573
rect 662156 95568 662295 95570
rect 662156 95512 662234 95568
rect 662290 95512 662295 95568
rect 662156 95510 662295 95512
rect 662156 95508 662162 95510
rect 662229 95507 662295 95510
rect 657353 94754 657419 94757
rect 657310 94752 657419 94754
rect 657310 94696 657358 94752
rect 657414 94696 657419 94752
rect 657310 94691 657419 94696
rect 627913 94482 627979 94485
rect 627913 94480 628268 94482
rect 627913 94424 627918 94480
rect 627974 94424 628268 94480
rect 627913 94422 628268 94424
rect 627913 94419 627979 94422
rect 657310 94180 657370 94691
rect 663241 93802 663307 93805
rect 663198 93800 663307 93802
rect 663198 93744 663246 93800
rect 663302 93744 663307 93800
rect 663198 93739 663307 93744
rect 627269 93530 627335 93533
rect 627269 93528 628268 93530
rect 627269 93472 627274 93528
rect 627330 93472 628268 93528
rect 627269 93470 628268 93472
rect 627269 93467 627335 93470
rect 655329 93394 655395 93397
rect 655329 93392 656788 93394
rect 655329 93336 655334 93392
rect 655390 93336 656788 93392
rect 663198 93364 663258 93739
rect 655329 93334 656788 93336
rect 655329 93331 655395 93334
rect 580809 93258 580875 93261
rect 576380 93256 580875 93258
rect 576380 93200 580814 93256
rect 580870 93200 580875 93256
rect 576380 93198 580875 93200
rect 580809 93195 580875 93198
rect 663333 93122 663399 93125
rect 663333 93120 663442 93122
rect 663333 93064 663338 93120
rect 663394 93064 663442 93120
rect 663333 93059 663442 93064
rect 642725 92714 642791 92717
rect 642725 92712 642834 92714
rect 642725 92656 642730 92712
rect 642786 92656 642834 92712
rect 642725 92651 642834 92656
rect 626441 92578 626507 92581
rect 626441 92576 628268 92578
rect 626441 92520 626446 92576
rect 626502 92520 628268 92576
rect 626441 92518 628268 92520
rect 626441 92515 626507 92518
rect 642774 92140 642834 92651
rect 653213 92578 653279 92581
rect 653213 92576 656788 92578
rect 653213 92520 653218 92576
rect 653274 92520 656788 92576
rect 663382 92548 663442 93059
rect 653213 92518 656788 92520
rect 653213 92515 653279 92518
rect 663425 92306 663491 92309
rect 663382 92304 663491 92306
rect 663382 92248 663430 92304
rect 663486 92248 663491 92304
rect 663382 92243 663491 92248
rect 580625 91762 580691 91765
rect 576380 91760 580691 91762
rect 576380 91704 580630 91760
rect 580686 91704 580691 91760
rect 663382 91732 663442 92243
rect 576380 91702 580691 91704
rect 580625 91699 580691 91702
rect 625889 91626 625955 91629
rect 625889 91624 628268 91626
rect 625889 91568 625894 91624
rect 625950 91568 628268 91624
rect 625889 91566 628268 91568
rect 625889 91563 625955 91566
rect 654041 91490 654107 91493
rect 654041 91488 656788 91490
rect 654041 91432 654046 91488
rect 654102 91432 656788 91488
rect 654041 91430 656788 91432
rect 654041 91427 654107 91430
rect 663241 91082 663307 91085
rect 663198 91080 663307 91082
rect 663198 91024 663246 91080
rect 663302 91024 663307 91080
rect 663198 91019 663307 91024
rect 623773 90674 623839 90677
rect 653489 90674 653555 90677
rect 623773 90672 628268 90674
rect 623773 90616 623778 90672
rect 623834 90616 628268 90672
rect 623773 90614 628268 90616
rect 653489 90672 656788 90674
rect 653489 90616 653494 90672
rect 653550 90616 656788 90672
rect 663198 90644 663258 91019
rect 653489 90614 656788 90616
rect 623773 90611 623839 90614
rect 653489 90611 653555 90614
rect 656985 90402 657051 90405
rect 663701 90402 663767 90405
rect 656942 90400 657051 90402
rect 656942 90344 656990 90400
rect 657046 90344 657051 90400
rect 656942 90339 657051 90344
rect 663566 90400 663767 90402
rect 663566 90344 663706 90400
rect 663762 90344 663767 90400
rect 663566 90342 663767 90344
rect 582005 90266 582071 90269
rect 576380 90264 582071 90266
rect 576380 90208 582010 90264
rect 582066 90208 582071 90264
rect 576380 90206 582071 90208
rect 582005 90203 582071 90206
rect 656942 89828 657002 90339
rect 663566 89828 663626 90342
rect 663701 90339 663767 90342
rect 623957 89722 624023 89725
rect 645945 89722 646011 89725
rect 623957 89720 628268 89722
rect 623957 89664 623962 89720
rect 624018 89664 628268 89720
rect 623957 89662 628268 89664
rect 642988 89720 646011 89722
rect 642988 89664 645950 89720
rect 646006 89664 646011 89720
rect 642988 89662 646011 89664
rect 623957 89659 624023 89662
rect 645945 89659 646011 89662
rect 663517 89586 663583 89589
rect 663517 89584 663626 89586
rect 663517 89528 663522 89584
rect 663578 89528 663626 89584
rect 663517 89523 663626 89528
rect 663566 89012 663626 89523
rect 623221 88906 623287 88909
rect 623221 88904 628268 88906
rect 623221 88848 623226 88904
rect 623282 88848 628268 88904
rect 623221 88846 628268 88848
rect 623221 88843 623287 88846
rect 662137 88772 662203 88773
rect 662086 88708 662092 88772
rect 662156 88770 662203 88772
rect 662156 88768 662248 88770
rect 662198 88712 662248 88768
rect 662156 88710 662248 88712
rect 662156 88708 662203 88710
rect 662137 88707 662203 88708
rect 582281 88634 582347 88637
rect 576380 88632 582347 88634
rect 576380 88576 582286 88632
rect 582342 88576 582347 88632
rect 576380 88574 582347 88576
rect 582281 88571 582347 88574
rect 622485 87954 622551 87957
rect 622485 87952 628268 87954
rect 622485 87896 622490 87952
rect 622546 87896 628268 87952
rect 622485 87894 628268 87896
rect 622485 87891 622551 87894
rect 582097 87138 582163 87141
rect 646037 87138 646103 87141
rect 576380 87136 582163 87138
rect 576380 87080 582102 87136
rect 582158 87080 582163 87136
rect 576380 87078 582163 87080
rect 642988 87136 646103 87138
rect 642988 87080 646042 87136
rect 646098 87080 646103 87136
rect 642988 87078 646103 87080
rect 582097 87075 582163 87078
rect 646037 87075 646103 87078
rect 622301 87002 622367 87005
rect 622301 87000 628268 87002
rect 622301 86944 622306 87000
rect 622362 86944 628268 87000
rect 622301 86942 628268 86944
rect 622301 86939 622367 86942
rect 623405 86050 623471 86053
rect 623405 86048 628268 86050
rect 623405 85992 623410 86048
rect 623466 85992 628268 86048
rect 623405 85990 628268 85992
rect 623405 85987 623471 85990
rect 581913 85642 581979 85645
rect 576380 85640 581979 85642
rect 576380 85584 581918 85640
rect 581974 85584 581979 85640
rect 576380 85582 581979 85584
rect 581913 85579 581979 85582
rect 623313 85098 623379 85101
rect 623313 85096 628268 85098
rect 623313 85040 623318 85096
rect 623374 85040 628268 85096
rect 623313 85038 628268 85040
rect 623313 85035 623379 85038
rect 646129 84690 646195 84693
rect 642988 84688 646195 84690
rect 642988 84632 646134 84688
rect 646190 84632 646195 84688
rect 642988 84630 646195 84632
rect 646129 84627 646195 84630
rect 581821 84146 581887 84149
rect 576380 84144 581887 84146
rect 576380 84088 581826 84144
rect 581882 84088 581887 84144
rect 576380 84086 581887 84088
rect 581821 84083 581887 84086
rect 621933 84146 621999 84149
rect 621933 84144 628268 84146
rect 621933 84088 621938 84144
rect 621994 84088 628268 84144
rect 621933 84086 628268 84088
rect 621933 84083 621999 84086
rect 623129 83194 623195 83197
rect 623129 83192 628268 83194
rect 623129 83136 623134 83192
rect 623190 83136 628268 83192
rect 623129 83134 628268 83136
rect 623129 83131 623195 83134
rect 579613 82650 579679 82653
rect 576380 82648 579679 82650
rect 576380 82592 579618 82648
rect 579674 82592 579679 82648
rect 576380 82590 579679 82592
rect 579613 82587 579679 82590
rect 622301 82242 622367 82245
rect 645853 82242 645919 82245
rect 622301 82240 628268 82242
rect 622301 82184 622306 82240
rect 622362 82184 628268 82240
rect 622301 82182 628268 82184
rect 642988 82240 645919 82242
rect 642988 82184 645858 82240
rect 645914 82184 645919 82240
rect 642988 82182 645919 82184
rect 622301 82179 622367 82182
rect 645853 82179 645919 82182
rect 622485 81426 622551 81429
rect 622485 81424 628268 81426
rect 622485 81368 622490 81424
rect 622546 81368 628268 81424
rect 622485 81366 628268 81368
rect 622485 81363 622551 81366
rect 581637 81154 581703 81157
rect 576380 81152 581703 81154
rect 576380 81096 581642 81152
rect 581698 81096 581703 81152
rect 576380 81094 581703 81096
rect 581637 81091 581703 81094
rect 581729 79522 581795 79525
rect 576380 79520 581795 79522
rect 576380 79464 581734 79520
rect 581790 79464 581795 79520
rect 576380 79462 581795 79464
rect 581729 79459 581795 79462
rect 581269 78026 581335 78029
rect 576380 78024 581335 78026
rect 576380 77968 581274 78024
rect 581330 77968 581335 78024
rect 576380 77966 581335 77968
rect 581269 77963 581335 77966
rect 581545 76530 581611 76533
rect 576380 76528 581611 76530
rect 576380 76472 581550 76528
rect 581606 76472 581611 76528
rect 576380 76470 581611 76472
rect 581545 76467 581611 76470
rect 581361 75034 581427 75037
rect 576380 75032 581427 75034
rect 576380 74976 581366 75032
rect 581422 74976 581427 75032
rect 576380 74974 581427 74976
rect 581361 74971 581427 74974
rect 580942 73538 580948 73540
rect 576380 73478 580948 73538
rect 580942 73476 580948 73478
rect 581012 73476 581018 73540
rect 581453 72042 581519 72045
rect 576380 72040 581519 72042
rect 576380 71984 581458 72040
rect 581514 71984 581519 72040
rect 576380 71982 581519 71984
rect 581453 71979 581519 71982
rect 581177 70410 581243 70413
rect 576380 70408 581243 70410
rect 576380 70352 581182 70408
rect 581238 70352 581243 70408
rect 576380 70350 581243 70352
rect 581177 70347 581243 70350
rect 582281 68914 582347 68917
rect 576380 68912 582347 68914
rect 576380 68856 582286 68912
rect 582342 68856 582347 68912
rect 576380 68854 582347 68856
rect 582281 68851 582347 68854
rect 581085 67418 581151 67421
rect 576380 67416 581151 67418
rect 576380 67360 581090 67416
rect 581146 67360 581151 67416
rect 576380 67358 581151 67360
rect 581085 67355 581151 67358
rect 580717 65922 580783 65925
rect 576380 65920 580783 65922
rect 576380 65864 580722 65920
rect 580778 65864 580783 65920
rect 576380 65862 580783 65864
rect 580717 65859 580783 65862
rect 580809 64426 580875 64429
rect 576380 64424 580875 64426
rect 576380 64368 580814 64424
rect 580870 64368 580875 64424
rect 576380 64366 580875 64368
rect 580809 64363 580875 64366
rect 582005 62930 582071 62933
rect 576380 62928 582071 62930
rect 576380 62872 582010 62928
rect 582066 62872 582071 62928
rect 576380 62870 582071 62872
rect 582005 62867 582071 62870
rect 582189 61298 582255 61301
rect 576380 61296 582255 61298
rect 576380 61240 582194 61296
rect 582250 61240 582255 61296
rect 576380 61238 582255 61240
rect 582189 61235 582255 61238
rect 579613 59802 579679 59805
rect 576380 59800 579679 59802
rect 576380 59744 579618 59800
rect 579674 59744 579679 59800
rect 576380 59742 579679 59744
rect 579613 59739 579679 59742
rect 579613 58306 579679 58309
rect 576380 58304 579679 58306
rect 576380 58248 579618 58304
rect 579674 58248 579679 58304
rect 576380 58246 579679 58248
rect 579613 58243 579679 58246
rect 581913 56810 581979 56813
rect 576380 56808 581979 56810
rect 576380 56752 581918 56808
rect 581974 56752 581979 56808
rect 576380 56750 581979 56752
rect 581913 56747 581979 56750
rect 582097 55314 582163 55317
rect 576380 55312 582163 55314
rect 576380 55256 582102 55312
rect 582158 55256 582163 55312
rect 576380 55254 582163 55256
rect 582097 55251 582163 55254
rect 580901 53818 580967 53821
rect 576380 53816 580967 53818
rect 576380 53760 580906 53816
rect 580962 53760 580967 53816
rect 576380 53758 580967 53760
rect 580901 53755 580967 53758
rect 646313 45114 646379 45117
rect 641394 45112 646379 45114
rect 641394 45056 646318 45112
rect 646374 45056 646379 45112
rect 641394 45054 646379 45056
rect 641394 44482 641454 45054
rect 646313 45051 646379 45054
rect 641302 43621 641362 43761
rect 641253 43616 641362 43621
rect 641253 43560 641258 43616
rect 641314 43560 641362 43616
rect 641253 43558 641362 43560
rect 641253 43555 641319 43558
rect 641161 42938 641227 42941
rect 641302 42938 641362 43396
rect 641161 42936 641362 42938
rect 641161 42880 641166 42936
rect 641222 42880 641362 42936
rect 641161 42878 641362 42880
rect 641161 42875 641227 42878
rect 194409 42258 194475 42261
rect 641253 42258 641319 42261
rect 194409 42256 641319 42258
rect 194409 42200 194414 42256
rect 194470 42200 641258 42256
rect 641314 42200 641319 42256
rect 194409 42198 641319 42200
rect 194409 42195 194475 42198
rect 641253 42195 641319 42198
rect 518525 42122 518591 42125
rect 521653 42122 521719 42125
rect 518525 42120 521719 42122
rect 518525 42064 518530 42120
rect 518586 42064 521658 42120
rect 521714 42064 521719 42120
rect 518525 42062 521719 42064
rect 518525 42059 518591 42062
rect 521653 42059 521719 42062
rect 415485 41986 415551 41989
rect 524045 41986 524111 41989
rect 415485 41984 524111 41986
rect 415485 41928 415490 41984
rect 415546 41928 524050 41984
rect 524106 41928 524111 41984
rect 415485 41926 524111 41928
rect 415485 41923 415551 41926
rect 524045 41923 524111 41926
rect 529657 41986 529723 41989
rect 535453 41986 535519 41989
rect 529657 41984 535519 41986
rect 529657 41928 529662 41984
rect 529718 41928 535458 41984
rect 535514 41928 535519 41984
rect 529657 41926 535519 41928
rect 529657 41923 529723 41926
rect 535453 41923 535519 41926
rect 187601 41850 187667 41853
rect 307293 41850 307359 41853
rect 362033 41850 362099 41853
rect 470317 41850 470383 41853
rect 594701 41850 594767 41853
rect 187601 41848 187710 41850
rect 187601 41792 187606 41848
rect 187662 41792 187710 41848
rect 187601 41787 187710 41792
rect 307293 41848 322950 41850
rect 307293 41792 307298 41848
rect 307354 41792 322950 41848
rect 307293 41790 322950 41792
rect 307293 41787 307359 41790
rect 187650 41306 187710 41787
rect 322890 41578 322950 41790
rect 362033 41848 380910 41850
rect 362033 41792 362038 41848
rect 362094 41792 380910 41848
rect 362033 41790 380910 41792
rect 362033 41787 362099 41790
rect 380850 41714 380910 41790
rect 470317 41848 594767 41850
rect 470317 41792 470322 41848
rect 470378 41792 594706 41848
rect 594762 41792 594767 41848
rect 470317 41790 594767 41792
rect 470317 41787 470383 41790
rect 594701 41787 594767 41790
rect 590745 41714 590811 41717
rect 380850 41712 590811 41714
rect 380850 41656 590750 41712
rect 590806 41656 590811 41712
rect 380850 41654 590811 41656
rect 590745 41651 590811 41654
rect 565813 41578 565879 41581
rect 322890 41576 565879 41578
rect 322890 41520 565818 41576
rect 565874 41520 565879 41576
rect 322890 41518 565879 41520
rect 565813 41515 565879 41518
rect 209773 41306 209839 41309
rect 212441 41306 212507 41309
rect 187650 41304 212507 41306
rect 187650 41248 209778 41304
rect 209834 41248 212446 41304
rect 212502 41248 212507 41304
rect 187650 41246 212507 41248
rect 209773 41243 209839 41246
rect 212441 41243 212507 41246
rect 218053 41306 218119 41309
rect 642633 41306 642699 41309
rect 218053 41304 642699 41306
rect 218053 41248 218058 41304
rect 218114 41248 642638 41304
rect 642694 41248 642699 41304
rect 218053 41246 642699 41248
rect 218053 41243 218119 41246
rect 642633 41243 642699 41246
rect 230841 16690 230907 16693
rect 225676 16688 230907 16690
rect 225676 16632 230846 16688
rect 230902 16632 230907 16688
rect 225676 16630 230907 16632
rect 230841 16627 230907 16630
rect 231025 15194 231091 15197
rect 225676 15192 231091 15194
rect 225676 15136 231030 15192
rect 231086 15136 231091 15192
rect 225676 15134 231091 15136
rect 231025 15131 231091 15134
rect 230749 13698 230815 13701
rect 225676 13696 230815 13698
rect 225676 13640 230754 13696
rect 230810 13640 230815 13696
rect 225676 13638 230815 13640
rect 230749 13635 230815 13638
rect 230933 12202 230999 12205
rect 225676 12200 230999 12202
rect 225676 12144 230938 12200
rect 230994 12144 230999 12200
rect 225676 12142 230999 12144
rect 230933 12139 230999 12142
rect 230473 10706 230539 10709
rect 225676 10704 230539 10706
rect 225676 10648 230478 10704
rect 230534 10648 230539 10704
rect 225676 10646 230539 10648
rect 230473 10643 230539 10646
rect 230657 9210 230723 9213
rect 225676 9208 230723 9210
rect 225676 9152 230662 9208
rect 230718 9152 230723 9208
rect 225676 9150 230723 9152
rect 230657 9147 230723 9150
rect 230565 7714 230631 7717
rect 225676 7712 230631 7714
rect 225676 7656 230570 7712
rect 230626 7656 230631 7712
rect 225676 7654 230631 7656
rect 230565 7651 230631 7654
rect 230381 6218 230447 6221
rect 225676 6216 230447 6218
rect 225676 6160 230386 6216
rect 230442 6160 230447 6216
rect 225676 6158 230447 6160
rect 230381 6155 230447 6158
<< via3 >>
rect 87828 996372 87892 996436
rect 87828 995616 87892 995620
rect 87828 995560 87842 995616
rect 87842 995560 87892 995616
rect 87828 995556 87892 995560
rect 187740 997188 187804 997252
rect 187740 995692 187804 995756
rect 476436 996372 476500 996436
rect 526116 996372 526180 996436
rect 476436 995480 476500 995484
rect 476436 995424 476486 995480
rect 476486 995424 476500 995480
rect 476436 995420 476500 995424
rect 526116 995480 526180 995484
rect 526116 995424 526166 995480
rect 526166 995424 526180 995480
rect 526116 995420 526180 995424
rect 674788 985764 674852 985828
rect 674972 985628 675036 985692
rect 44036 985492 44100 985556
rect 43484 985356 43548 985420
rect 43668 983316 43732 983380
rect 43300 983180 43364 983244
rect 43852 983044 43916 983108
rect 43116 982908 43180 982972
rect 41460 968764 41524 968828
rect 41644 965092 41708 965156
rect 41828 963384 41892 963388
rect 41828 963328 41842 963384
rect 41842 963328 41892 963384
rect 41828 963324 41892 963328
rect 41828 949452 41892 949516
rect 673868 938300 673932 938364
rect 676812 937212 676876 937276
rect 674788 937076 674852 937140
rect 41828 936940 41892 937004
rect 674972 936260 675036 936324
rect 42012 935308 42076 935372
rect 43116 927148 43180 927212
rect 42564 921980 42628 922044
rect 43484 921980 43548 922044
rect 676076 877236 676140 877300
rect 675708 876616 675772 876620
rect 675708 876560 675722 876616
rect 675722 876560 675772 876616
rect 675708 876556 675772 876560
rect 675340 875936 675404 875940
rect 675340 875880 675390 875936
rect 675390 875880 675404 875936
rect 675340 875876 675404 875880
rect 675524 874032 675588 874036
rect 675524 873976 675538 874032
rect 675538 873976 675588 874032
rect 675524 873972 675588 873976
rect 675892 872204 675956 872268
rect 41828 814132 41892 814196
rect 676260 797676 676324 797740
rect 676444 791964 676508 792028
rect 674972 787748 675036 787812
rect 674604 787340 674668 787404
rect 675156 786796 675220 786860
rect 674788 784076 674852 784140
rect 674420 783804 674484 783868
rect 674236 777412 674300 777476
rect 39988 773060 40052 773124
rect 676812 772652 676876 772716
rect 39988 771428 40052 771492
rect 674236 770264 674300 770268
rect 674236 770208 674250 770264
rect 674250 770208 674300 770264
rect 674236 770204 674300 770208
rect 673868 760276 673932 760340
rect 42012 757072 42076 757076
rect 42012 757016 42026 757072
rect 42026 757016 42076 757072
rect 42012 757012 42076 757016
rect 675340 757012 675404 757076
rect 676076 756332 676140 756396
rect 675524 755788 675588 755852
rect 675708 754564 675772 754628
rect 42012 754080 42076 754084
rect 42012 754024 42062 754080
rect 42062 754024 42076 754080
rect 42012 754020 42076 754024
rect 675892 752524 675956 752588
rect 676444 752252 676508 752316
rect 676260 751844 676324 751908
rect 676628 744092 676692 744156
rect 676260 743956 676324 744020
rect 675892 742868 675956 742932
rect 676076 742460 676140 742524
rect 674236 741644 674300 741708
rect 675340 739800 675404 739804
rect 675340 739744 675390 739800
rect 675390 739744 675404 739800
rect 675340 739740 675404 739744
rect 673868 739060 673932 739124
rect 675708 738576 675772 738580
rect 675708 738520 675722 738576
rect 675722 738520 675772 738576
rect 675708 738516 675772 738520
rect 676444 737972 676508 738036
rect 39988 731036 40052 731100
rect 44036 728452 44100 728516
rect 675156 711996 675220 712060
rect 674972 711180 675036 711244
rect 676260 710534 676324 710598
rect 676628 710594 676692 710598
rect 676628 710538 676642 710594
rect 676642 710538 676692 710594
rect 676628 710534 676692 710538
rect 674604 709548 674668 709612
rect 674788 709140 674852 709204
rect 674420 708732 674484 708796
rect 676260 699756 676324 699820
rect 676812 699620 676876 699684
rect 676996 699484 677060 699548
rect 675524 698184 675588 698188
rect 675524 698128 675538 698184
rect 675538 698128 675588 698184
rect 675524 698124 675588 698128
rect 673684 697308 673748 697372
rect 674420 696628 674484 696692
rect 674604 694724 674668 694788
rect 673500 694316 673564 694380
rect 674052 693500 674116 693564
rect 677180 692956 677244 693020
rect 676628 690100 676692 690164
rect 41276 686700 41340 686764
rect 39988 684252 40052 684316
rect 41644 684252 41708 684316
rect 44036 683980 44100 684044
rect 30604 677316 30668 677380
rect 30604 676908 30668 676972
rect 677548 666980 677612 667044
rect 674236 666844 674300 666908
rect 675892 666028 675956 666092
rect 675340 665620 675404 665684
rect 676076 664532 676140 664596
rect 673868 663988 673932 664052
rect 675708 663580 675772 663644
rect 676260 662900 676324 662964
rect 676444 662492 676508 662556
rect 676996 662084 677060 662148
rect 676812 661676 676876 661740
rect 674972 652836 675036 652900
rect 674788 652156 674852 652220
rect 675156 651612 675220 651676
rect 675340 648952 675404 648956
rect 675340 648896 675390 648952
rect 675390 648896 675404 648952
rect 675340 648892 675404 648896
rect 675892 648620 675956 648684
rect 39988 643452 40052 643516
rect 673868 623052 673932 623116
rect 677364 622780 677428 622844
rect 674420 621828 674484 621892
rect 673868 621556 673932 621620
rect 675524 621012 675588 621076
rect 674604 620604 674668 620668
rect 673684 619380 673748 619444
rect 673500 618972 673564 619036
rect 674052 618564 674116 618628
rect 677180 617476 677244 617540
rect 676628 617068 676692 617132
rect 676444 608908 676508 608972
rect 676628 608772 676692 608836
rect 675708 607608 675772 607612
rect 675708 607552 675722 607608
rect 675722 607552 675772 607608
rect 675708 607548 675772 607552
rect 676076 607276 676140 607340
rect 674604 606460 674668 606524
rect 674420 604692 674484 604756
rect 675524 604344 675588 604348
rect 675524 604288 675538 604344
rect 675538 604288 675588 604344
rect 675524 604284 675588 604288
rect 674236 603468 674300 603532
rect 676260 602924 676324 602988
rect 43852 600476 43916 600540
rect 40172 598572 40236 598636
rect 43668 598028 43732 598092
rect 40172 596124 40236 596188
rect 673868 578172 673932 578236
rect 675156 576540 675220 576604
rect 674972 575724 675036 575788
rect 674788 574092 674852 574156
rect 675340 573684 675404 573748
rect 675892 573276 675956 573340
rect 676628 571916 676692 571980
rect 676444 571508 676508 571572
rect 676812 564436 676876 564500
rect 675340 562396 675404 562460
rect 675892 561988 675956 562052
rect 675156 561172 675220 561236
rect 674972 558724 675036 558788
rect 676444 558316 676508 558380
rect 676628 557500 676692 557564
rect 41644 557092 41708 557156
rect 43852 556004 43916 556068
rect 39988 555460 40052 555524
rect 40172 555460 40236 555524
rect 41828 554780 41892 554844
rect 41828 540908 41892 540972
rect 41644 540772 41708 540836
rect 674604 531796 674668 531860
rect 675708 530776 675772 530840
rect 674420 530572 674484 530636
rect 676076 529348 676140 529412
rect 675524 528940 675588 529004
rect 674236 528532 674300 528596
rect 676260 527308 676324 527372
rect 676812 526900 676876 526964
rect 673500 489228 673564 489292
rect 673868 488412 673932 488476
rect 675156 487596 675220 487660
rect 675340 486780 675404 486844
rect 675892 485148 675956 485212
rect 674972 484740 675036 484804
rect 676076 484468 676140 484532
rect 676076 483380 676140 483444
rect 43852 428844 43916 428908
rect 41828 427892 41892 427956
rect 39988 427790 40052 427854
rect 41828 427212 41892 427276
rect 673868 400964 673932 401028
rect 42932 386276 42996 386340
rect 39988 384644 40052 384708
rect 40172 384644 40236 384708
rect 42748 383964 42812 384028
rect 40356 383828 40420 383892
rect 42748 383420 42812 383484
rect 40172 383012 40236 383076
rect 41460 382196 41524 382260
rect 674052 357444 674116 357508
rect 674420 355812 674484 355876
rect 41460 355676 41524 355740
rect 674236 354996 674300 355060
rect 676076 353636 676140 353700
rect 675892 352140 675956 352204
rect 42932 351868 42996 351932
rect 675708 350508 675772 350572
rect 40172 341396 40236 341460
rect 42748 340444 42812 340508
rect 42564 339356 42628 339420
rect 41828 339220 41892 339284
rect 41644 337316 41708 337380
rect 42196 337180 42260 337244
rect 42012 336772 42076 336836
rect 675708 330576 675772 330580
rect 675708 330520 675722 330576
rect 675722 330520 675772 330576
rect 675708 330516 675772 330520
rect 41460 329836 41524 329900
rect 42380 329700 42444 329764
rect 676076 328340 676140 328404
rect 675892 326844 675956 326908
rect 41460 319908 41524 319972
rect 42012 316976 42076 316980
rect 42012 316920 42026 316976
rect 42026 316920 42076 316976
rect 42012 316916 42076 316920
rect 40356 316100 40420 316164
rect 42196 316024 42260 316028
rect 42196 315968 42210 316024
rect 42210 315968 42260 316024
rect 42196 315964 42260 315968
rect 42380 315420 42444 315484
rect 42564 313788 42628 313852
rect 41644 313108 41708 313172
rect 41828 312352 41892 312356
rect 41828 312296 41842 312352
rect 41842 312296 41892 312352
rect 41828 312292 41892 312296
rect 675892 306308 675956 306372
rect 41828 300052 41892 300116
rect 41828 298420 41892 298484
rect 42012 297604 42076 297668
rect 42012 295156 42076 295220
rect 675892 292164 675956 292228
rect 42196 285908 42260 285972
rect 42380 285772 42444 285836
rect 42564 285636 42628 285700
rect 44036 278428 44100 278492
rect 674420 278292 674484 278356
rect 674052 278156 674116 278220
rect 674236 278020 674300 278084
rect 673868 277884 673932 277948
rect 673684 277748 673748 277812
rect 673500 277612 673564 277676
rect 42012 272368 42076 272372
rect 42012 272312 42026 272368
rect 42026 272312 42076 272368
rect 42012 272308 42076 272312
rect 42380 270404 42444 270468
rect 42196 270056 42260 270060
rect 42196 270000 42210 270056
rect 42210 270000 42260 270056
rect 42196 269996 42260 270000
rect 42564 269180 42628 269244
rect 674236 264556 674300 264620
rect 674236 262380 674300 262444
rect 676076 262380 676140 262444
rect 42196 256804 42260 256868
rect 41460 256260 41524 256324
rect 41460 255444 41524 255508
rect 41644 255036 41708 255100
rect 42012 254356 42076 254420
rect 41828 253948 41892 254012
rect 42012 252724 42076 252788
rect 42012 225992 42076 225996
rect 42012 225936 42026 225992
rect 42026 225936 42076 225992
rect 42012 225932 42076 225936
rect 676076 219948 676140 220012
rect 42196 213284 42260 213348
rect 675892 213284 675956 213348
rect 675892 212468 675956 212532
rect 41644 211788 41708 211852
rect 41828 210836 41892 210900
rect 42748 210428 42812 210492
rect 41644 209340 41708 209404
rect 42380 209204 42444 209268
rect 42564 208796 42628 208860
rect 41828 207980 41892 208044
rect 42196 207572 42260 207636
rect 42012 207164 42076 207228
rect 41460 205668 41524 205732
rect 42564 190164 42628 190228
rect 41460 187580 41524 187644
rect 42012 187096 42076 187100
rect 42012 187040 42026 187096
rect 42026 187040 42076 187096
rect 42012 187036 42076 187040
rect 42196 186356 42260 186420
rect 42380 185812 42444 185876
rect 42748 184180 42812 184244
rect 41828 183696 41892 183700
rect 41828 183640 41842 183696
rect 41842 183640 41892 183696
rect 41828 183636 41892 183640
rect 41644 182684 41708 182748
rect 675892 173572 675956 173636
rect 676076 171804 676140 171868
rect 675892 148412 675956 148476
rect 676076 146236 676140 146300
rect 676076 128148 676140 128212
rect 675892 126788 675956 126852
rect 580948 113188 581012 113252
rect 676076 103260 676140 103324
rect 675892 101356 675956 101420
rect 662092 95508 662156 95572
rect 662092 88768 662156 88772
rect 662092 88712 662142 88768
rect 662142 88712 662156 88768
rect 662092 88708 662156 88712
rect 580948 73476 581012 73540
<< metal4 >>
rect 187739 997252 187805 997253
rect 187739 997188 187740 997252
rect 187804 997188 187805 997252
rect 187739 997187 187805 997188
rect 87827 996436 87893 996437
rect 87827 996372 87828 996436
rect 87892 996372 87893 996436
rect 87827 996371 87893 996372
rect 87830 995621 87890 996371
rect 187742 995757 187802 997187
rect 476435 996436 476501 996437
rect 476435 996372 476436 996436
rect 476500 996372 476501 996436
rect 476435 996371 476501 996372
rect 526115 996436 526181 996437
rect 526115 996372 526116 996436
rect 526180 996372 526181 996436
rect 526115 996371 526181 996372
rect 187739 995756 187805 995757
rect 187739 995692 187740 995756
rect 187804 995692 187805 995756
rect 187739 995691 187805 995692
rect 87827 995620 87893 995621
rect 87827 995556 87828 995620
rect 87892 995556 87893 995620
rect 87827 995555 87893 995556
rect 476438 995485 476498 996371
rect 526118 995485 526178 996371
rect 476435 995484 476501 995485
rect 476435 995420 476436 995484
rect 476500 995420 476501 995484
rect 476435 995419 476501 995420
rect 526115 995484 526181 995485
rect 526115 995420 526116 995484
rect 526180 995420 526181 995484
rect 526115 995419 526181 995420
rect 674787 985828 674853 985829
rect 674787 985764 674788 985828
rect 674852 985764 674853 985828
rect 674787 985763 674853 985764
rect 44035 985556 44101 985557
rect 44035 985492 44036 985556
rect 44100 985492 44101 985556
rect 44035 985491 44101 985492
rect 43483 985420 43549 985421
rect 43483 985356 43484 985420
rect 43548 985356 43549 985420
rect 43483 985355 43549 985356
rect 43299 983244 43365 983245
rect 43299 983180 43300 983244
rect 43364 983180 43365 983244
rect 43299 983179 43365 983180
rect 43115 982972 43181 982973
rect 43115 982908 43116 982972
rect 43180 982908 43181 982972
rect 43115 982907 43181 982908
rect 41459 968828 41525 968829
rect 41459 968764 41460 968828
rect 41524 968764 41525 968828
rect 41459 968763 41525 968764
rect 41462 937410 41522 968763
rect 41643 965156 41709 965157
rect 41643 965092 41644 965156
rect 41708 965092 41709 965156
rect 41643 965091 41709 965092
rect 41646 938090 41706 965091
rect 41827 963388 41893 963389
rect 41827 963324 41828 963388
rect 41892 963324 41893 963388
rect 41827 963323 41893 963324
rect 41830 949517 41890 963323
rect 41827 949516 41893 949517
rect 41827 949452 41828 949516
rect 41892 949452 41893 949516
rect 41827 949451 41893 949452
rect 41646 938030 42074 938090
rect 41462 937350 41890 937410
rect 41830 937005 41890 937350
rect 41827 937004 41893 937005
rect 41827 936940 41828 937004
rect 41892 936940 41893 937004
rect 41827 936939 41893 936940
rect 42014 935373 42074 938030
rect 42011 935372 42077 935373
rect 42011 935308 42012 935372
rect 42076 935308 42077 935372
rect 42011 935307 42077 935308
rect 43118 927213 43178 982907
rect 43115 927212 43181 927213
rect 43115 927148 43116 927212
rect 43180 927148 43181 927212
rect 43115 927147 43181 927148
rect 43302 922450 43362 983179
rect 42566 922390 43362 922450
rect 42566 922045 42626 922390
rect 43486 922045 43546 985355
rect 43667 983380 43733 983381
rect 43667 983316 43668 983380
rect 43732 983316 43733 983380
rect 43667 983315 43733 983316
rect 42563 922044 42629 922045
rect 42563 921980 42564 922044
rect 42628 921980 42629 922044
rect 42563 921979 42629 921980
rect 43483 922044 43549 922045
rect 43483 921980 43484 922044
rect 43548 921980 43549 922044
rect 43483 921979 43549 921980
rect 39990 814270 41890 814330
rect 39990 773125 40050 814270
rect 41830 814197 41890 814270
rect 41827 814196 41893 814197
rect 41827 814132 41828 814196
rect 41892 814132 41893 814196
rect 41827 814131 41893 814132
rect 39987 773124 40053 773125
rect 39987 773060 39988 773124
rect 40052 773060 40053 773124
rect 39987 773059 40053 773060
rect 39987 771492 40053 771493
rect 39987 771428 39988 771492
rect 40052 771428 40053 771492
rect 39987 771427 40053 771428
rect 39990 731101 40050 771427
rect 42011 757076 42077 757077
rect 42011 757012 42012 757076
rect 42076 757012 42077 757076
rect 42011 757011 42077 757012
rect 42014 754085 42074 757011
rect 42011 754084 42077 754085
rect 42011 754020 42012 754084
rect 42076 754020 42077 754084
rect 42011 754019 42077 754020
rect 39987 731100 40053 731101
rect 39987 731036 39988 731100
rect 40052 731036 40053 731100
rect 39987 731035 40053 731036
rect 41275 686764 41341 686765
rect 41275 686700 41276 686764
rect 41340 686700 41341 686764
rect 41275 686699 41341 686700
rect 41278 684450 41338 686699
rect 41278 684390 41706 684450
rect 41646 684317 41706 684390
rect 39987 684316 40053 684317
rect 39987 684252 39988 684316
rect 40052 684252 40053 684316
rect 39987 684251 40053 684252
rect 41643 684316 41709 684317
rect 41643 684252 41644 684316
rect 41708 684252 41709 684316
rect 41643 684251 41709 684252
rect 30603 677380 30669 677381
rect 30603 677316 30604 677380
rect 30668 677316 30669 677380
rect 30603 677315 30669 677316
rect 30606 676973 30666 677315
rect 30603 676972 30669 676973
rect 30603 676908 30604 676972
rect 30668 676908 30669 676972
rect 30603 676907 30669 676908
rect 39990 643517 40050 684251
rect 39987 643516 40053 643517
rect 39987 643452 39988 643516
rect 40052 643452 40053 643516
rect 39987 643451 40053 643452
rect 40171 598636 40237 598637
rect 40171 598572 40172 598636
rect 40236 598572 40237 598636
rect 40171 598571 40237 598572
rect 40174 596189 40234 598571
rect 43670 598093 43730 983315
rect 43851 983108 43917 983109
rect 43851 983044 43852 983108
rect 43916 983044 43917 983108
rect 43851 983043 43917 983044
rect 43854 600541 43914 983043
rect 44038 728517 44098 985491
rect 673867 938364 673933 938365
rect 673867 938300 673868 938364
rect 673932 938300 673933 938364
rect 673867 938299 673933 938300
rect 673870 760341 673930 938299
rect 674790 937141 674850 985763
rect 674971 985692 675037 985693
rect 674971 985628 674972 985692
rect 675036 985628 675037 985692
rect 674971 985627 675037 985628
rect 674787 937140 674853 937141
rect 674787 937076 674788 937140
rect 674852 937076 674853 937140
rect 674787 937075 674853 937076
rect 674974 936325 675034 985627
rect 676811 937276 676877 937277
rect 676811 937212 676812 937276
rect 676876 937212 676877 937276
rect 676811 937211 676877 937212
rect 674971 936324 675037 936325
rect 674971 936260 674972 936324
rect 675036 936260 675037 936324
rect 674971 936259 675037 936260
rect 676075 877300 676141 877301
rect 676075 877236 676076 877300
rect 676140 877236 676141 877300
rect 676075 877235 676141 877236
rect 675707 876620 675773 876621
rect 675707 876556 675708 876620
rect 675772 876556 675773 876620
rect 675707 876555 675773 876556
rect 675339 875940 675405 875941
rect 675339 875876 675340 875940
rect 675404 875876 675405 875940
rect 675339 875875 675405 875876
rect 674971 787812 675037 787813
rect 674971 787748 674972 787812
rect 675036 787748 675037 787812
rect 674971 787747 675037 787748
rect 674603 787404 674669 787405
rect 674603 787340 674604 787404
rect 674668 787340 674669 787404
rect 674603 787339 674669 787340
rect 674419 783868 674485 783869
rect 674419 783804 674420 783868
rect 674484 783804 674485 783868
rect 674419 783803 674485 783804
rect 674235 777476 674301 777477
rect 674235 777412 674236 777476
rect 674300 777412 674301 777476
rect 674235 777411 674301 777412
rect 674238 770269 674298 777411
rect 674235 770268 674301 770269
rect 674235 770204 674236 770268
rect 674300 770204 674301 770268
rect 674235 770203 674301 770204
rect 673867 760340 673933 760341
rect 673867 760276 673868 760340
rect 673932 760276 673933 760340
rect 673867 760275 673933 760276
rect 674235 741708 674301 741709
rect 674235 741644 674236 741708
rect 674300 741644 674301 741708
rect 674235 741643 674301 741644
rect 673867 739124 673933 739125
rect 673867 739060 673868 739124
rect 673932 739060 673933 739124
rect 673867 739059 673933 739060
rect 44035 728516 44101 728517
rect 44035 728452 44036 728516
rect 44100 728452 44101 728516
rect 44035 728451 44101 728452
rect 673683 697372 673749 697373
rect 673683 697308 673684 697372
rect 673748 697308 673749 697372
rect 673683 697307 673749 697308
rect 673499 694380 673565 694381
rect 673499 694316 673500 694380
rect 673564 694316 673565 694380
rect 673499 694315 673565 694316
rect 44035 684044 44101 684045
rect 44035 683980 44036 684044
rect 44100 683980 44101 684044
rect 44035 683979 44101 683980
rect 43851 600540 43917 600541
rect 43851 600476 43852 600540
rect 43916 600476 43917 600540
rect 43851 600475 43917 600476
rect 43667 598092 43733 598093
rect 43667 598028 43668 598092
rect 43732 598028 43733 598092
rect 43667 598027 43733 598028
rect 40171 596188 40237 596189
rect 40171 596124 40172 596188
rect 40236 596124 40237 596188
rect 40171 596123 40237 596124
rect 40174 555525 40234 596123
rect 41643 557156 41709 557157
rect 41643 557092 41644 557156
rect 41708 557092 41709 557156
rect 41643 557091 41709 557092
rect 39987 555524 40053 555525
rect 39987 555460 39988 555524
rect 40052 555460 40053 555524
rect 39987 555459 40053 555460
rect 40171 555524 40237 555525
rect 40171 555460 40172 555524
rect 40236 555460 40237 555524
rect 40171 555459 40237 555460
rect 39990 428090 40050 555459
rect 41646 540837 41706 557091
rect 43851 556068 43917 556069
rect 43851 556004 43852 556068
rect 43916 556004 43917 556068
rect 43851 556003 43917 556004
rect 41827 554844 41893 554845
rect 41827 554780 41828 554844
rect 41892 554780 41893 554844
rect 41827 554779 41893 554780
rect 41830 540973 41890 554779
rect 41827 540972 41893 540973
rect 41827 540908 41828 540972
rect 41892 540908 41893 540972
rect 41827 540907 41893 540908
rect 41643 540836 41709 540837
rect 41643 540772 41644 540836
rect 41708 540772 41709 540836
rect 41643 540771 41709 540772
rect 43854 428909 43914 556003
rect 43851 428908 43917 428909
rect 43851 428844 43852 428908
rect 43916 428844 43917 428908
rect 43851 428843 43917 428844
rect 39990 428030 41890 428090
rect 41830 427957 41890 428030
rect 41827 427956 41893 427957
rect 41827 427892 41828 427956
rect 41892 427892 41893 427956
rect 41827 427891 41893 427892
rect 39987 427854 40053 427855
rect 39987 427790 39988 427854
rect 40052 427790 40053 427854
rect 39987 427789 40053 427790
rect 39990 425070 40050 427789
rect 41827 427276 41893 427277
rect 41827 427212 41828 427276
rect 41892 427212 41893 427276
rect 41827 427211 41893 427212
rect 41830 425070 41890 427211
rect 39990 425010 40234 425070
rect 40174 411270 40234 425010
rect 39990 411210 40234 411270
rect 40358 425010 41890 425070
rect 39990 384709 40050 411210
rect 39987 384708 40053 384709
rect 39987 384644 39988 384708
rect 40052 384644 40053 384708
rect 39987 384643 40053 384644
rect 40171 384708 40237 384709
rect 40171 384644 40172 384708
rect 40236 384644 40237 384708
rect 40171 384643 40237 384644
rect 39990 322950 40050 384643
rect 40174 383077 40234 384643
rect 40358 383893 40418 425010
rect 42931 386340 42997 386341
rect 42931 386276 42932 386340
rect 42996 386276 42997 386340
rect 42931 386275 42997 386276
rect 42747 384028 42813 384029
rect 42747 383964 42748 384028
rect 42812 383964 42813 384028
rect 42747 383963 42813 383964
rect 40355 383892 40421 383893
rect 40355 383828 40356 383892
rect 40420 383828 40421 383892
rect 40355 383827 40421 383828
rect 42750 383485 42810 383963
rect 42747 383484 42813 383485
rect 42747 383420 42748 383484
rect 42812 383420 42813 383484
rect 42747 383419 42813 383420
rect 40171 383076 40237 383077
rect 40171 383012 40172 383076
rect 40236 383012 40237 383076
rect 40171 383011 40237 383012
rect 40174 341461 40234 383011
rect 41459 382260 41525 382261
rect 41459 382196 41460 382260
rect 41524 382196 41525 382260
rect 41459 382195 41525 382196
rect 41462 355741 41522 382195
rect 41459 355740 41525 355741
rect 41459 355676 41460 355740
rect 41524 355676 41525 355740
rect 41459 355675 41525 355676
rect 40171 341460 40237 341461
rect 40171 341396 40172 341460
rect 40236 341396 40237 341460
rect 40171 341395 40237 341396
rect 42750 340509 42810 383419
rect 42934 351933 42994 386275
rect 42931 351932 42997 351933
rect 42931 351868 42932 351932
rect 42996 351868 42997 351932
rect 42931 351867 42997 351868
rect 42747 340508 42813 340509
rect 42747 340444 42748 340508
rect 42812 340444 42813 340508
rect 42747 340443 42813 340444
rect 42563 339420 42629 339421
rect 42563 339356 42564 339420
rect 42628 339356 42629 339420
rect 42563 339355 42629 339356
rect 41827 339284 41893 339285
rect 41827 339220 41828 339284
rect 41892 339220 41893 339284
rect 41827 339219 41893 339220
rect 41643 337380 41709 337381
rect 41643 337316 41644 337380
rect 41708 337316 41709 337380
rect 41643 337315 41709 337316
rect 41459 329900 41525 329901
rect 41459 329836 41460 329900
rect 41524 329836 41525 329900
rect 41459 329835 41525 329836
rect 39990 322890 40418 322950
rect 40358 316165 40418 322890
rect 41462 319973 41522 329835
rect 41459 319972 41525 319973
rect 41459 319908 41460 319972
rect 41524 319908 41525 319972
rect 41459 319907 41525 319908
rect 40355 316164 40421 316165
rect 40355 316100 40356 316164
rect 40420 316100 40421 316164
rect 40355 316099 40421 316100
rect 41646 313173 41706 337315
rect 41643 313172 41709 313173
rect 41643 313108 41644 313172
rect 41708 313108 41709 313172
rect 41643 313107 41709 313108
rect 41830 312357 41890 339219
rect 42195 337244 42261 337245
rect 42195 337180 42196 337244
rect 42260 337180 42261 337244
rect 42195 337179 42261 337180
rect 42011 336836 42077 336837
rect 42011 336772 42012 336836
rect 42076 336772 42077 336836
rect 42011 336771 42077 336772
rect 42014 316981 42074 336771
rect 42011 316980 42077 316981
rect 42011 316916 42012 316980
rect 42076 316916 42077 316980
rect 42011 316915 42077 316916
rect 42198 316029 42258 337179
rect 42379 329764 42445 329765
rect 42379 329700 42380 329764
rect 42444 329700 42445 329764
rect 42379 329699 42445 329700
rect 42195 316028 42261 316029
rect 42195 315964 42196 316028
rect 42260 315964 42261 316028
rect 42195 315963 42261 315964
rect 42382 315485 42442 329699
rect 42379 315484 42445 315485
rect 42379 315420 42380 315484
rect 42444 315420 42445 315484
rect 42379 315419 42445 315420
rect 42566 313853 42626 339355
rect 42563 313852 42629 313853
rect 42563 313788 42564 313852
rect 42628 313788 42629 313852
rect 42563 313787 42629 313788
rect 41827 312356 41893 312357
rect 41827 312292 41828 312356
rect 41892 312292 41893 312356
rect 41827 312291 41893 312292
rect 41827 300116 41893 300117
rect 41827 300052 41828 300116
rect 41892 300052 41893 300116
rect 41827 300051 41893 300052
rect 41830 298890 41890 300051
rect 41462 298830 41890 298890
rect 41462 256325 41522 298830
rect 41827 298484 41893 298485
rect 41827 298420 41828 298484
rect 41892 298420 41893 298484
rect 41827 298419 41893 298420
rect 41830 296170 41890 298419
rect 42011 297668 42077 297669
rect 42011 297604 42012 297668
rect 42076 297604 42077 297668
rect 42011 297603 42077 297604
rect 41646 296110 41890 296170
rect 41459 256324 41525 256325
rect 41459 256260 41460 256324
rect 41524 256260 41525 256324
rect 41459 256259 41525 256260
rect 41459 255508 41525 255509
rect 41459 255444 41460 255508
rect 41524 255444 41525 255508
rect 41459 255443 41525 255444
rect 41462 245670 41522 255443
rect 41646 255101 41706 296110
rect 42014 295490 42074 297603
rect 41830 295430 42074 295490
rect 41643 255100 41709 255101
rect 41643 255036 41644 255100
rect 41708 255036 41709 255100
rect 41643 255035 41709 255036
rect 41830 254013 41890 295430
rect 42011 295220 42077 295221
rect 42011 295156 42012 295220
rect 42076 295156 42077 295220
rect 42011 295155 42077 295156
rect 42014 272373 42074 295155
rect 42195 285972 42261 285973
rect 42195 285908 42196 285972
rect 42260 285908 42261 285972
rect 42195 285907 42261 285908
rect 42011 272372 42077 272373
rect 42011 272308 42012 272372
rect 42076 272308 42077 272372
rect 42011 272307 42077 272308
rect 42198 270061 42258 285907
rect 42379 285836 42445 285837
rect 42379 285772 42380 285836
rect 42444 285772 42445 285836
rect 42379 285771 42445 285772
rect 42382 270469 42442 285771
rect 42563 285700 42629 285701
rect 42563 285636 42564 285700
rect 42628 285636 42629 285700
rect 42563 285635 42629 285636
rect 42379 270468 42445 270469
rect 42379 270404 42380 270468
rect 42444 270404 42445 270468
rect 42379 270403 42445 270404
rect 42195 270060 42261 270061
rect 42195 269996 42196 270060
rect 42260 269996 42261 270060
rect 42195 269995 42261 269996
rect 42566 269245 42626 285635
rect 44038 278493 44098 683979
rect 673502 619037 673562 694315
rect 673686 619445 673746 697307
rect 673870 664053 673930 739059
rect 674051 693564 674117 693565
rect 674051 693500 674052 693564
rect 674116 693500 674117 693564
rect 674051 693499 674117 693500
rect 673867 664052 673933 664053
rect 673867 663988 673868 664052
rect 673932 663988 673933 664052
rect 673867 663987 673933 663988
rect 673867 623116 673933 623117
rect 673867 623052 673868 623116
rect 673932 623052 673933 623116
rect 673867 623051 673933 623052
rect 673870 621621 673930 623051
rect 673867 621620 673933 621621
rect 673867 621556 673868 621620
rect 673932 621556 673933 621620
rect 673867 621555 673933 621556
rect 673683 619444 673749 619445
rect 673683 619380 673684 619444
rect 673748 619380 673749 619444
rect 673683 619379 673749 619380
rect 673499 619036 673565 619037
rect 673499 618972 673500 619036
rect 673564 618972 673565 619036
rect 673499 618971 673565 618972
rect 673870 578237 673930 621555
rect 674054 618629 674114 693499
rect 674238 666909 674298 741643
rect 674422 708797 674482 783803
rect 674606 709613 674666 787339
rect 674787 784140 674853 784141
rect 674787 784076 674788 784140
rect 674852 784076 674853 784140
rect 674787 784075 674853 784076
rect 674603 709612 674669 709613
rect 674603 709548 674604 709612
rect 674668 709548 674669 709612
rect 674603 709547 674669 709548
rect 674790 709205 674850 784075
rect 674974 711245 675034 787747
rect 675155 786860 675221 786861
rect 675155 786796 675156 786860
rect 675220 786796 675221 786860
rect 675155 786795 675221 786796
rect 675158 712061 675218 786795
rect 675342 757077 675402 875875
rect 675523 874036 675589 874037
rect 675523 873972 675524 874036
rect 675588 873972 675589 874036
rect 675523 873971 675589 873972
rect 675339 757076 675405 757077
rect 675339 757012 675340 757076
rect 675404 757012 675405 757076
rect 675339 757011 675405 757012
rect 675526 755853 675586 873971
rect 675523 755852 675589 755853
rect 675523 755788 675524 755852
rect 675588 755788 675589 755852
rect 675523 755787 675589 755788
rect 675710 754629 675770 876555
rect 675891 872268 675957 872269
rect 675891 872204 675892 872268
rect 675956 872204 675957 872268
rect 675891 872203 675957 872204
rect 675707 754628 675773 754629
rect 675707 754564 675708 754628
rect 675772 754564 675773 754628
rect 675707 754563 675773 754564
rect 675894 752589 675954 872203
rect 676078 756397 676138 877235
rect 676259 797740 676325 797741
rect 676259 797676 676260 797740
rect 676324 797676 676325 797740
rect 676259 797675 676325 797676
rect 676075 756396 676141 756397
rect 676075 756332 676076 756396
rect 676140 756332 676141 756396
rect 676075 756331 676141 756332
rect 675891 752588 675957 752589
rect 675891 752524 675892 752588
rect 675956 752524 675957 752588
rect 675891 752523 675957 752524
rect 676262 751909 676322 797675
rect 676443 792028 676509 792029
rect 676443 791964 676444 792028
rect 676508 791964 676509 792028
rect 676443 791963 676509 791964
rect 676446 752317 676506 791963
rect 676814 772717 676874 937211
rect 676811 772716 676877 772717
rect 676811 772652 676812 772716
rect 676876 772652 676877 772716
rect 676811 772651 676877 772652
rect 676443 752316 676509 752317
rect 676443 752252 676444 752316
rect 676508 752252 676509 752316
rect 676443 752251 676509 752252
rect 676259 751908 676325 751909
rect 676259 751844 676260 751908
rect 676324 751844 676325 751908
rect 676259 751843 676325 751844
rect 676627 744156 676693 744157
rect 676627 744092 676628 744156
rect 676692 744092 676693 744156
rect 676627 744091 676693 744092
rect 676259 744020 676325 744021
rect 676259 743956 676260 744020
rect 676324 743956 676325 744020
rect 676259 743955 676325 743956
rect 675891 742932 675957 742933
rect 675891 742868 675892 742932
rect 675956 742868 675957 742932
rect 675891 742867 675957 742868
rect 675339 739804 675405 739805
rect 675339 739740 675340 739804
rect 675404 739740 675405 739804
rect 675339 739739 675405 739740
rect 675155 712060 675221 712061
rect 675155 711996 675156 712060
rect 675220 711996 675221 712060
rect 675155 711995 675221 711996
rect 674971 711244 675037 711245
rect 674971 711180 674972 711244
rect 675036 711180 675037 711244
rect 674971 711179 675037 711180
rect 674787 709204 674853 709205
rect 674787 709140 674788 709204
rect 674852 709140 674853 709204
rect 674787 709139 674853 709140
rect 674419 708796 674485 708797
rect 674419 708732 674420 708796
rect 674484 708732 674485 708796
rect 674419 708731 674485 708732
rect 674419 696692 674485 696693
rect 674419 696628 674420 696692
rect 674484 696628 674485 696692
rect 674419 696627 674485 696628
rect 674235 666908 674301 666909
rect 674235 666844 674236 666908
rect 674300 666844 674301 666908
rect 674235 666843 674301 666844
rect 674422 621893 674482 696627
rect 674603 694788 674669 694789
rect 674603 694724 674604 694788
rect 674668 694724 674669 694788
rect 674603 694723 674669 694724
rect 674419 621892 674485 621893
rect 674419 621828 674420 621892
rect 674484 621828 674485 621892
rect 674419 621827 674485 621828
rect 674606 620669 674666 694723
rect 675342 665685 675402 739739
rect 675707 738580 675773 738581
rect 675707 738516 675708 738580
rect 675772 738516 675773 738580
rect 675707 738515 675773 738516
rect 675523 698188 675589 698189
rect 675523 698124 675524 698188
rect 675588 698124 675589 698188
rect 675523 698123 675589 698124
rect 675339 665684 675405 665685
rect 675339 665620 675340 665684
rect 675404 665620 675405 665684
rect 675339 665619 675405 665620
rect 674971 652900 675037 652901
rect 674971 652836 674972 652900
rect 675036 652836 675037 652900
rect 674971 652835 675037 652836
rect 674787 652220 674853 652221
rect 674787 652156 674788 652220
rect 674852 652156 674853 652220
rect 674787 652155 674853 652156
rect 674603 620668 674669 620669
rect 674603 620604 674604 620668
rect 674668 620604 674669 620668
rect 674603 620603 674669 620604
rect 674051 618628 674117 618629
rect 674051 618564 674052 618628
rect 674116 618564 674117 618628
rect 674051 618563 674117 618564
rect 674603 606524 674669 606525
rect 674603 606460 674604 606524
rect 674668 606460 674669 606524
rect 674603 606459 674669 606460
rect 674419 604756 674485 604757
rect 674419 604692 674420 604756
rect 674484 604692 674485 604756
rect 674419 604691 674485 604692
rect 674235 603532 674301 603533
rect 674235 603468 674236 603532
rect 674300 603468 674301 603532
rect 674235 603467 674301 603468
rect 673867 578236 673933 578237
rect 673867 578172 673868 578236
rect 673932 578172 673933 578236
rect 673867 578171 673933 578172
rect 674238 528597 674298 603467
rect 674422 530637 674482 604691
rect 674606 531861 674666 606459
rect 674790 574157 674850 652155
rect 674974 575789 675034 652835
rect 675155 651676 675221 651677
rect 675155 651612 675156 651676
rect 675220 651612 675221 651676
rect 675155 651611 675221 651612
rect 675158 576605 675218 651611
rect 675339 648956 675405 648957
rect 675339 648892 675340 648956
rect 675404 648892 675405 648956
rect 675339 648891 675405 648892
rect 675155 576604 675221 576605
rect 675155 576540 675156 576604
rect 675220 576540 675221 576604
rect 675155 576539 675221 576540
rect 674971 575788 675037 575789
rect 674971 575724 674972 575788
rect 675036 575724 675037 575788
rect 674971 575723 675037 575724
rect 674787 574156 674853 574157
rect 674787 574092 674788 574156
rect 674852 574092 674853 574156
rect 674787 574091 674853 574092
rect 675342 573749 675402 648891
rect 675526 621077 675586 698123
rect 675710 663645 675770 738515
rect 675894 666093 675954 742867
rect 676075 742524 676141 742525
rect 676075 742460 676076 742524
rect 676140 742460 676141 742524
rect 676075 742459 676141 742460
rect 675891 666092 675957 666093
rect 675891 666028 675892 666092
rect 675956 666028 675957 666092
rect 675891 666027 675957 666028
rect 676078 664597 676138 742459
rect 676262 710599 676322 743955
rect 676443 738036 676509 738037
rect 676443 737972 676444 738036
rect 676508 737972 676509 738036
rect 676443 737971 676509 737972
rect 676259 710598 676325 710599
rect 676259 710534 676260 710598
rect 676324 710534 676325 710598
rect 676259 710533 676325 710534
rect 676259 699820 676325 699821
rect 676259 699756 676260 699820
rect 676324 699756 676325 699820
rect 676259 699755 676325 699756
rect 676075 664596 676141 664597
rect 676075 664532 676076 664596
rect 676140 664532 676141 664596
rect 676075 664531 676141 664532
rect 675707 663644 675773 663645
rect 675707 663580 675708 663644
rect 675772 663580 675773 663644
rect 675707 663579 675773 663580
rect 676262 662965 676322 699755
rect 676259 662964 676325 662965
rect 676259 662900 676260 662964
rect 676324 662900 676325 662964
rect 676259 662899 676325 662900
rect 676446 662557 676506 737971
rect 676630 710599 676690 744091
rect 676627 710598 676693 710599
rect 676627 710534 676628 710598
rect 676692 710534 676693 710598
rect 676627 710533 676693 710534
rect 676811 699684 676877 699685
rect 676811 699620 676812 699684
rect 676876 699620 676877 699684
rect 676811 699619 676877 699620
rect 676627 690164 676693 690165
rect 676627 690100 676628 690164
rect 676692 690100 676693 690164
rect 676627 690099 676693 690100
rect 676443 662556 676509 662557
rect 676443 662492 676444 662556
rect 676508 662492 676509 662556
rect 676443 662491 676509 662492
rect 675891 648684 675957 648685
rect 675891 648620 675892 648684
rect 675956 648620 675957 648684
rect 675891 648619 675957 648620
rect 675523 621076 675589 621077
rect 675523 621012 675524 621076
rect 675588 621012 675589 621076
rect 675523 621011 675589 621012
rect 675707 607612 675773 607613
rect 675707 607548 675708 607612
rect 675772 607548 675773 607612
rect 675707 607547 675773 607548
rect 675523 604348 675589 604349
rect 675523 604284 675524 604348
rect 675588 604284 675589 604348
rect 675523 604283 675589 604284
rect 675339 573748 675405 573749
rect 675339 573684 675340 573748
rect 675404 573684 675405 573748
rect 675339 573683 675405 573684
rect 675339 562460 675405 562461
rect 675339 562396 675340 562460
rect 675404 562396 675405 562460
rect 675339 562395 675405 562396
rect 675155 561236 675221 561237
rect 675155 561172 675156 561236
rect 675220 561172 675221 561236
rect 675155 561171 675221 561172
rect 674971 558788 675037 558789
rect 674971 558724 674972 558788
rect 675036 558724 675037 558788
rect 674971 558723 675037 558724
rect 674603 531860 674669 531861
rect 674603 531796 674604 531860
rect 674668 531796 674669 531860
rect 674603 531795 674669 531796
rect 674419 530636 674485 530637
rect 674419 530572 674420 530636
rect 674484 530572 674485 530636
rect 674419 530571 674485 530572
rect 674235 528596 674301 528597
rect 674235 528532 674236 528596
rect 674300 528532 674301 528596
rect 674235 528531 674301 528532
rect 673499 489292 673565 489293
rect 673499 489228 673500 489292
rect 673564 489228 673565 489292
rect 673499 489227 673565 489228
rect 673502 488550 673562 489227
rect 673502 488490 673746 488550
rect 673686 458190 673746 488490
rect 673867 488476 673933 488477
rect 673867 488412 673868 488476
rect 673932 488412 673933 488476
rect 673867 488411 673933 488412
rect 673502 458130 673746 458190
rect 44035 278492 44101 278493
rect 44035 278428 44036 278492
rect 44100 278428 44101 278492
rect 44035 278427 44101 278428
rect 673502 277677 673562 458130
rect 673870 438870 673930 488411
rect 674974 484805 675034 558723
rect 675158 487661 675218 561171
rect 675155 487660 675221 487661
rect 675155 487596 675156 487660
rect 675220 487596 675221 487660
rect 675155 487595 675221 487596
rect 675342 486845 675402 562395
rect 675526 529005 675586 604283
rect 675710 530841 675770 607547
rect 675894 573341 675954 648619
rect 676630 617133 676690 690099
rect 676814 661741 676874 699619
rect 676995 699548 677061 699549
rect 676995 699484 676996 699548
rect 677060 699484 677061 699548
rect 676995 699483 677061 699484
rect 676998 662149 677058 699483
rect 677179 693020 677245 693021
rect 677179 692956 677180 693020
rect 677244 692956 677245 693020
rect 677179 692955 677245 692956
rect 677182 676230 677242 692955
rect 677182 676170 677426 676230
rect 676995 662148 677061 662149
rect 676995 662084 676996 662148
rect 677060 662084 677061 662148
rect 676995 662083 677061 662084
rect 676811 661740 676877 661741
rect 676811 661676 676812 661740
rect 676876 661676 676877 661740
rect 676811 661675 676877 661676
rect 677366 656910 677426 676170
rect 677547 667044 677613 667045
rect 677547 666980 677548 667044
rect 677612 666980 677613 667044
rect 677547 666979 677613 666980
rect 677182 656850 677426 656910
rect 677182 617541 677242 656850
rect 677550 632070 677610 666979
rect 677366 632010 677610 632070
rect 677366 622845 677426 632010
rect 677363 622844 677429 622845
rect 677363 622780 677364 622844
rect 677428 622780 677429 622844
rect 677363 622779 677429 622780
rect 677179 617540 677245 617541
rect 677179 617476 677180 617540
rect 677244 617476 677245 617540
rect 677179 617475 677245 617476
rect 676627 617132 676693 617133
rect 676627 617068 676628 617132
rect 676692 617068 676693 617132
rect 676627 617067 676693 617068
rect 676443 608972 676509 608973
rect 676443 608908 676444 608972
rect 676508 608908 676509 608972
rect 676443 608907 676509 608908
rect 676075 607340 676141 607341
rect 676075 607276 676076 607340
rect 676140 607276 676141 607340
rect 676075 607275 676141 607276
rect 675891 573340 675957 573341
rect 675891 573276 675892 573340
rect 675956 573276 675957 573340
rect 675891 573275 675957 573276
rect 675891 562052 675957 562053
rect 675891 561988 675892 562052
rect 675956 561988 675957 562052
rect 675891 561987 675957 561988
rect 675707 530840 675773 530841
rect 675707 530776 675708 530840
rect 675772 530776 675773 530840
rect 675707 530775 675773 530776
rect 675523 529004 675589 529005
rect 675523 528940 675524 529004
rect 675588 528940 675589 529004
rect 675523 528939 675589 528940
rect 675339 486844 675405 486845
rect 675339 486780 675340 486844
rect 675404 486780 675405 486844
rect 675339 486779 675405 486780
rect 675894 485213 675954 561987
rect 676078 529413 676138 607275
rect 676259 602988 676325 602989
rect 676259 602924 676260 602988
rect 676324 602924 676325 602988
rect 676259 602923 676325 602924
rect 676075 529412 676141 529413
rect 676075 529348 676076 529412
rect 676140 529348 676141 529412
rect 676075 529347 676141 529348
rect 676262 527373 676322 602923
rect 676446 571573 676506 608907
rect 676627 608836 676693 608837
rect 676627 608772 676628 608836
rect 676692 608772 676693 608836
rect 676627 608771 676693 608772
rect 676630 571981 676690 608771
rect 676627 571980 676693 571981
rect 676627 571916 676628 571980
rect 676692 571916 676693 571980
rect 676627 571915 676693 571916
rect 676443 571572 676509 571573
rect 676443 571508 676444 571572
rect 676508 571508 676509 571572
rect 676443 571507 676509 571508
rect 676811 564500 676877 564501
rect 676811 564436 676812 564500
rect 676876 564436 676877 564500
rect 676811 564435 676877 564436
rect 676443 558380 676509 558381
rect 676443 558316 676444 558380
rect 676508 558316 676509 558380
rect 676443 558315 676509 558316
rect 676259 527372 676325 527373
rect 676259 527308 676260 527372
rect 676324 527308 676325 527372
rect 676259 527307 676325 527308
rect 675891 485212 675957 485213
rect 675891 485148 675892 485212
rect 675956 485148 675957 485212
rect 675891 485147 675957 485148
rect 674971 484804 675037 484805
rect 674971 484740 674972 484804
rect 675036 484740 675037 484804
rect 674971 484739 675037 484740
rect 676075 484532 676141 484533
rect 676075 484468 676076 484532
rect 676140 484530 676141 484532
rect 676446 484530 676506 558315
rect 676627 557564 676693 557565
rect 676627 557500 676628 557564
rect 676692 557500 676693 557564
rect 676627 557499 676693 557500
rect 676140 484470 676506 484530
rect 676140 484468 676141 484470
rect 676075 484467 676141 484468
rect 676075 483444 676141 483445
rect 676075 483380 676076 483444
rect 676140 483380 676141 483444
rect 676630 483442 676690 557499
rect 676814 526965 676874 564435
rect 676811 526964 676877 526965
rect 676811 526900 676812 526964
rect 676876 526900 676877 526964
rect 676811 526899 676877 526900
rect 676075 483379 676141 483380
rect 676262 483382 676690 483442
rect 676078 483170 676138 483379
rect 676262 483170 676322 483382
rect 676078 483110 676322 483170
rect 673686 438810 673930 438870
rect 673686 277813 673746 438810
rect 673867 401028 673933 401029
rect 673867 400964 673868 401028
rect 673932 400964 673933 401028
rect 673867 400963 673933 400964
rect 673870 277949 673930 400963
rect 674051 357508 674117 357509
rect 674051 357444 674052 357508
rect 674116 357444 674117 357508
rect 674051 357443 674117 357444
rect 674054 278221 674114 357443
rect 674419 355876 674485 355877
rect 674419 355812 674420 355876
rect 674484 355812 674485 355876
rect 674419 355811 674485 355812
rect 674235 355060 674301 355061
rect 674235 354996 674236 355060
rect 674300 354996 674301 355060
rect 674235 354995 674301 354996
rect 674051 278220 674117 278221
rect 674051 278156 674052 278220
rect 674116 278156 674117 278220
rect 674051 278155 674117 278156
rect 674238 278085 674298 354995
rect 674422 278357 674482 355811
rect 676075 353700 676141 353701
rect 676075 353636 676076 353700
rect 676140 353636 676141 353700
rect 676075 353635 676141 353636
rect 675891 352204 675957 352205
rect 675891 352140 675892 352204
rect 675956 352140 675957 352204
rect 675891 352139 675957 352140
rect 675707 350572 675773 350573
rect 675707 350508 675708 350572
rect 675772 350508 675773 350572
rect 675707 350507 675773 350508
rect 675710 330581 675770 350507
rect 675707 330580 675773 330581
rect 675707 330516 675708 330580
rect 675772 330516 675773 330580
rect 675707 330515 675773 330516
rect 675894 326909 675954 352139
rect 676078 328405 676138 353635
rect 676075 328404 676141 328405
rect 676075 328340 676076 328404
rect 676140 328340 676141 328404
rect 676075 328339 676141 328340
rect 675891 326908 675957 326909
rect 675891 326844 675892 326908
rect 675956 326844 675957 326908
rect 675891 326843 675957 326844
rect 675891 306372 675957 306373
rect 675891 306308 675892 306372
rect 675956 306308 675957 306372
rect 675891 306307 675957 306308
rect 675894 292229 675954 306307
rect 675891 292228 675957 292229
rect 675891 292164 675892 292228
rect 675956 292164 675957 292228
rect 675891 292163 675957 292164
rect 674419 278356 674485 278357
rect 674419 278292 674420 278356
rect 674484 278292 674485 278356
rect 674419 278291 674485 278292
rect 674235 278084 674301 278085
rect 674235 278020 674236 278084
rect 674300 278020 674301 278084
rect 674235 278019 674301 278020
rect 673867 277948 673933 277949
rect 673867 277884 673868 277948
rect 673932 277884 673933 277948
rect 673867 277883 673933 277884
rect 673683 277812 673749 277813
rect 673683 277748 673684 277812
rect 673748 277748 673749 277812
rect 673683 277747 673749 277748
rect 673499 277676 673565 277677
rect 673499 277612 673500 277676
rect 673564 277612 673565 277676
rect 673499 277611 673565 277612
rect 42563 269244 42629 269245
rect 42563 269180 42564 269244
rect 42628 269180 42629 269244
rect 42563 269179 42629 269180
rect 674235 264620 674301 264621
rect 674235 264556 674236 264620
rect 674300 264556 674301 264620
rect 674235 264555 674301 264556
rect 674238 262445 674298 264555
rect 674235 262444 674301 262445
rect 674235 262380 674236 262444
rect 674300 262380 674301 262444
rect 674235 262379 674301 262380
rect 676075 262444 676141 262445
rect 676075 262380 676076 262444
rect 676140 262380 676141 262444
rect 676075 262379 676141 262380
rect 42195 256868 42261 256869
rect 42195 256804 42196 256868
rect 42260 256804 42261 256868
rect 42195 256803 42261 256804
rect 42011 254420 42077 254421
rect 42011 254356 42012 254420
rect 42076 254356 42077 254420
rect 42011 254355 42077 254356
rect 41827 254012 41893 254013
rect 41827 253948 41828 254012
rect 41892 253948 41893 254012
rect 41827 253947 41893 253948
rect 42014 253330 42074 254355
rect 41830 253270 42074 253330
rect 41462 245610 41706 245670
rect 41646 211853 41706 245610
rect 41643 211852 41709 211853
rect 41643 211788 41644 211852
rect 41708 211788 41709 211852
rect 41643 211787 41709 211788
rect 41830 210901 41890 253270
rect 42011 252788 42077 252789
rect 42011 252724 42012 252788
rect 42076 252724 42077 252788
rect 42011 252723 42077 252724
rect 42014 225997 42074 252723
rect 42011 225996 42077 225997
rect 42011 225932 42012 225996
rect 42076 225932 42077 225996
rect 42011 225931 42077 225932
rect 42198 213349 42258 256803
rect 676078 220013 676138 262379
rect 676075 220012 676141 220013
rect 676075 219948 676076 220012
rect 676140 219948 676141 220012
rect 676075 219947 676141 219948
rect 42195 213348 42261 213349
rect 42195 213284 42196 213348
rect 42260 213284 42261 213348
rect 42195 213283 42261 213284
rect 675891 213348 675957 213349
rect 675891 213284 675892 213348
rect 675956 213284 675957 213348
rect 675891 213283 675957 213284
rect 675894 212533 675954 213283
rect 675891 212532 675957 212533
rect 675891 212468 675892 212532
rect 675956 212468 675957 212532
rect 675891 212467 675957 212468
rect 41827 210900 41893 210901
rect 41827 210836 41828 210900
rect 41892 210836 41893 210900
rect 41827 210835 41893 210836
rect 42747 210492 42813 210493
rect 42747 210428 42748 210492
rect 42812 210428 42813 210492
rect 42747 210427 42813 210428
rect 41643 209404 41709 209405
rect 41643 209340 41644 209404
rect 41708 209340 41709 209404
rect 41643 209339 41709 209340
rect 41459 205732 41525 205733
rect 41459 205668 41460 205732
rect 41524 205668 41525 205732
rect 41459 205667 41525 205668
rect 41462 187645 41522 205667
rect 41459 187644 41525 187645
rect 41459 187580 41460 187644
rect 41524 187580 41525 187644
rect 41459 187579 41525 187580
rect 41646 182749 41706 209339
rect 42379 209268 42445 209269
rect 42379 209204 42380 209268
rect 42444 209204 42445 209268
rect 42379 209203 42445 209204
rect 41827 208044 41893 208045
rect 41827 207980 41828 208044
rect 41892 207980 41893 208044
rect 41827 207979 41893 207980
rect 41830 183701 41890 207979
rect 42195 207636 42261 207637
rect 42195 207572 42196 207636
rect 42260 207572 42261 207636
rect 42195 207571 42261 207572
rect 42011 207228 42077 207229
rect 42011 207164 42012 207228
rect 42076 207164 42077 207228
rect 42011 207163 42077 207164
rect 42014 187101 42074 207163
rect 42011 187100 42077 187101
rect 42011 187036 42012 187100
rect 42076 187036 42077 187100
rect 42011 187035 42077 187036
rect 42198 186421 42258 207571
rect 42195 186420 42261 186421
rect 42195 186356 42196 186420
rect 42260 186356 42261 186420
rect 42195 186355 42261 186356
rect 42382 185877 42442 209203
rect 42563 208860 42629 208861
rect 42563 208796 42564 208860
rect 42628 208796 42629 208860
rect 42563 208795 42629 208796
rect 42566 190229 42626 208795
rect 42563 190228 42629 190229
rect 42563 190164 42564 190228
rect 42628 190164 42629 190228
rect 42563 190163 42629 190164
rect 42379 185876 42445 185877
rect 42379 185812 42380 185876
rect 42444 185812 42445 185876
rect 42379 185811 42445 185812
rect 42750 184245 42810 210427
rect 42747 184244 42813 184245
rect 42747 184180 42748 184244
rect 42812 184180 42813 184244
rect 42747 184179 42813 184180
rect 41827 183700 41893 183701
rect 41827 183636 41828 183700
rect 41892 183636 41893 183700
rect 41827 183635 41893 183636
rect 41643 182748 41709 182749
rect 41643 182684 41644 182748
rect 41708 182684 41709 182748
rect 41643 182683 41709 182684
rect 675891 173636 675957 173637
rect 675891 173572 675892 173636
rect 675956 173572 675957 173636
rect 675891 173571 675957 173572
rect 675894 148477 675954 173571
rect 676075 171868 676141 171869
rect 676075 171804 676076 171868
rect 676140 171804 676141 171868
rect 676075 171803 676141 171804
rect 675891 148476 675957 148477
rect 675891 148412 675892 148476
rect 675956 148412 675957 148476
rect 675891 148411 675957 148412
rect 676078 146301 676138 171803
rect 676075 146300 676141 146301
rect 676075 146236 676076 146300
rect 676140 146236 676141 146300
rect 676075 146235 676141 146236
rect 676075 128212 676141 128213
rect 676075 128148 676076 128212
rect 676140 128148 676141 128212
rect 676075 128147 676141 128148
rect 675891 126852 675957 126853
rect 675891 126788 675892 126852
rect 675956 126788 675957 126852
rect 675891 126787 675957 126788
rect 580947 113252 581013 113253
rect 580947 113188 580948 113252
rect 581012 113188 581013 113252
rect 580947 113187 581013 113188
rect 580950 73541 581010 113187
rect 675894 101421 675954 126787
rect 676078 103325 676138 128147
rect 676075 103324 676141 103325
rect 676075 103260 676076 103324
rect 676140 103260 676141 103324
rect 676075 103259 676141 103260
rect 675891 101420 675957 101421
rect 675891 101356 675892 101420
rect 675956 101356 675957 101420
rect 675891 101355 675957 101356
rect 662091 95572 662157 95573
rect 662091 95508 662092 95572
rect 662156 95508 662157 95572
rect 662091 95507 662157 95508
rect 662094 88773 662154 95507
rect 662091 88772 662157 88773
rect 662091 88708 662092 88772
rect 662156 88708 662157 88772
rect 662091 88707 662157 88708
rect 580947 73540 581013 73541
rect 580947 73476 580948 73540
rect 581012 73476 581013 73540
rect 580947 73475 581013 73476
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030788
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030788
rect 628240 1018512 640760 1031002
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876160
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18975 123778
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use user_id_programming  user_id_value
timestamp 1637275745
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1637275745
transform 1 0 52034 0 1 53002
box 382 -400 524400 164400
use xres_buf  rstb_level
timestamp 1637275745
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use simple_por  por
timestamp 1637275745
transform 1 0 630146 0 -1 51282
box 25 11 11344 8291
use digital_pll  pll
timestamp 1637275745
transform 1 0 628146 0 1 80944
box 0 0 15000 15000
use housekeeping  housekeeping
timestamp 1637275745
transform 1 0 606434 0 1 100002
box 0 0 60047 110190
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1637275745
transform -1 0 710203 0 1 121000
box 750 416 34000 13000
use gpio_defaults_block  gpio_01_defaults\[0\]
timestamp 1637275745
transform 1 0 703487 0 1 134000
box -38 0 6018 2224
use caravel_clocking  clocking
timestamp 1637275745
transform 1 0 205746 0 1 5488
box -38 -48 20000 12000
use gpio_defaults_block  gpio_37_defaults
timestamp 1637275745
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1637275745
transform 1 0 7631 0 1 202600
box 750 416 34000 13000
use gpio_defaults_block  gpio_01_defaults\[1\]
timestamp 1637275745
transform 1 0 703487 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1637275745
transform -1 0 710203 0 1 166200
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1637275745
transform -1 0 710203 0 1 211200
box 750 416 34000 13000
use gpio_defaults_block  gpio_36_defaults
timestamp 1637275745
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1637275745
transform 1 0 7631 0 1 245800
box 750 416 34000 13000
use mgmt_protect  mgmt_buffers
timestamp 1637275745
transform 1 0 192180 0 1 240036
box -400 -400 220400 24400
use gpio_defaults_block  gpio_234_defaults\[0\]
timestamp 1637275745
transform 1 0 703487 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_234_defaults\[1\]
timestamp 1637275745
transform 1 0 703487 0 1 269400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1637275745
transform -1 0 710203 0 1 256400
box 750 416 34000 13000
use gpio_defaults_block  gpio_35_defaults
timestamp 1637275745
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1637275745
transform 1 0 7631 0 1 289000
box 750 416 34000 13000
use gpio_defaults_block  gpio_234_defaults\[2\]
timestamp 1637275745
transform 1 0 703487 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1637275745
transform -1 0 710203 0 1 301400
box 750 416 34000 13000
use gpio_defaults_block  gpio_32_defaults
timestamp 1637275745
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_33_defaults
timestamp 1637275745
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_34_defaults
timestamp 1637275745
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1637275745
transform 1 0 7631 0 1 418600
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1637275745
transform 1 0 7631 0 1 375400
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1637275745
transform 1 0 7631 0 1 332200
box 750 416 34000 13000
use gpio_defaults_block  gpio_5_defaults
timestamp 1637275745
transform 1 0 703487 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_6_defaults
timestamp 1637275745
transform 1 0 703487 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_7_defaults
timestamp 1637275745
transform 1 0 703487 0 1 492800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1637275745
transform -1 0 710203 0 1 346400
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1637275745
transform -1 0 710203 0 1 391600
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1637275745
transform -1 0 710203 0 1 479800
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1637275745
transform 1 0 7631 0 1 546200
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1637275745
transform 1 0 7631 0 1 589400
box 750 416 34000 13000
use gpio_defaults_block  gpio_31_defaults
timestamp 1637275745
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_30_defaults
timestamp 1637275745
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1637275745
transform -1 0 710203 0 1 568800
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1637275745
transform -1 0 710203 0 1 523800
box 750 416 34000 13000
use gpio_defaults_block  gpio_9_defaults
timestamp 1637275745
transform 1 0 703487 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_8_defaults
timestamp 1637275745
transform 1 0 703487 0 1 536800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1637275745
transform 1 0 7631 0 1 675800
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1637275745
transform 1 0 7631 0 1 632600
box 750 416 34000 13000
use gpio_defaults_block  gpio_29_defaults
timestamp 1637275745
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_28_defaults
timestamp 1637275745
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1637275745
transform -1 0 710203 0 1 659000
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1637275745
transform -1 0 710203 0 1 614000
box 750 416 34000 13000
use gpio_defaults_block  gpio_11_defaults
timestamp 1637275745
transform 1 0 703487 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_10_defaults
timestamp 1637275745
transform 1 0 703487 0 1 627000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1637275745
transform 1 0 7631 0 1 719000
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1637275745
transform 1 0 7631 0 1 762200
box 750 416 34000 13000
use gpio_defaults_block  gpio_27_defaults
timestamp 1637275745
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_26_defaults
timestamp 1637275745
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1637275745
transform -1 0 710203 0 1 749200
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1637275745
transform -1 0 710203 0 1 704200
box 750 416 34000 13000
use gpio_defaults_block  gpio_13_defaults
timestamp 1637275745
transform 1 0 703487 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_12_defaults
timestamp 1637275745
transform 1 0 703487 0 1 717200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1637275745
transform 1 0 7631 0 1 805400
box 750 416 34000 13000
use gpio_defaults_block  gpio_25_defaults
timestamp 1637275745
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1637275745
transform 1 0 7631 0 1 931200
box 750 416 34000 13000
use gpio_defaults_block  gpio_24_defaults
timestamp 1637275745
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1637275745
transform -1 0 710203 0 1 927600
box 750 416 34000 13000
use gpio_defaults_block  gpio_14_defaults
timestamp 1637275745
transform 1 0 703487 0 1 940600
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1637275745
transform 0 1 97200 -1 0 1030077
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1637275745
transform 0 1 148600 -1 0 1030077
box 750 416 34000 13000
use gpio_defaults_block  gpio_23_defaults
timestamp 1637275745
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_22_defaults
timestamp 1637275745
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1637275745
transform 0 1 200000 -1 0 1030077
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1637275745
transform 0 1 251400 -1 0 1030077
box 750 416 34000 13000
use gpio_defaults_block  gpio_21_defaults
timestamp 1637275745
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1637275745
transform 0 1 303000 -1 0 1030077
box 750 416 34000 13000
use gpio_defaults_block  gpio_20_defaults
timestamp 1637275745
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_19_defaults
timestamp 1637275745
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1637275745
transform 0 1 420800 -1 0 1030077
box 750 416 34000 13000
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1637275745
transform 0 1 353400 -1 0 1030077
box 750 416 34000 13000
use gpio_defaults_block  gpio_18_defaults
timestamp 1637275745
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_17_defaults
timestamp 1637275745
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1637275745
transform 0 1 497800 -1 0 1030077
box 750 416 34000 13000
use gpio_defaults_block  gpio_16_defaults
timestamp 1637275745
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1637275745
transform 0 1 549200 -1 0 1030077
box 750 416 34000 13000
use gpio_defaults_block  gpio_15_defaults
timestamp 1637275745
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use user_project_wrapper  mprj
timestamp 1637275745
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use chip_io  padframe
timestamp 1637275745
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144149 18309 6 resetb
port 44 nsew signal input
rlabel metal5 s 6167 70054 19619 80934 6 vccd
port 45 nsew signal bidirectional
rlabel metal5 s 697980 909666 711432 920546 6 vccd1
port 46 nsew signal bidirectional
rlabel metal5 s 6167 914054 19619 924934 6 vccd2
port 47 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18975 6 vdda
port 48 nsew signal bidirectional
rlabel metal5 s 698624 819822 710788 831990 6 vdda1
port 49 nsew signal bidirectional
rlabel metal5 s 698624 505222 710788 517390 6 vdda1_2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 484410 18975 496578 6 vdda2
port 51 nsew signal bidirectional
rlabel metal5 s 6811 111610 18975 123778 6 vddio
port 52 nsew signal bidirectional
rlabel metal5 s 6811 871210 18975 883378 6 vddio_2
port 53 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18975 6 vssa
port 54 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030788 6 vssa1
port 55 nsew signal bidirectional
rlabel metal5 s 698624 417022 710788 429190 6 vssa1_2
port 56 nsew signal bidirectional
rlabel metal5 s 6811 829010 18975 841178 6 vssa2
port 57 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19619 6 vssd
port 58 nsew signal bidirectional
rlabel metal5 s 697980 461866 711432 472746 6 vssd1
port 59 nsew signal bidirectional
rlabel metal5 s 6167 442854 19619 453734 6 vssd2
port 60 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18975 6 vssio
port 61 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030788 6 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
