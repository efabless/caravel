VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_logic_high
  CLASS BLOCK ;
  FOREIGN gpio_logic_high ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.000 BY 22.000 ;
  PIN gpio_logic1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 2.000 ;
    END
  END gpio_logic1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.660 2.480 2.260 19.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 8.260 2.480 9.860 19.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.860 2.480 17.460 19.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.220 2.920 21.400 4.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.220 10.520 21.400 12.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.220 18.120 21.400 19.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 4.260 2.480 5.860 19.280 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.860 2.480 13.460 19.280 ;
    END
    PORT
      LAYER met2 ;
        RECT 19.460 2.480 21.060 19.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.220 6.520 21.400 8.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.220 14.120 21.400 15.720 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 0.460 2.635 21.160 19.125 ;
      LAYER met1 ;
        RECT 0.460 2.480 21.160 19.280 ;
      LAYER met2 ;
        RECT 10.680 2.280 10.940 17.670 ;
  END
END gpio_logic_high
END LIBRARY

