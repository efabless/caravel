* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for mprj2_logic_high abstract view
.subckt mprj2_logic_high HI vccd2 vssd2
.ends

* Black-box entry subcircuit for mprj_logic_high abstract view
.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46]
+ HI[47] HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57]
+ HI[58] HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68]
+ HI[69] HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79]
+ HI[7] HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8]
+ HI[90] HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1
+ vssd1
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv vccd vssd vdda1 vssa1 vdda2 vssa2 mprj2_vdd_logic1 mprj_vdd_logic1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd vccd1_uq1 vccd2_uq0 vdda1_uq0 vdda2_uq0 vssd vssd2_uq0
+ vssa1_uq0 vssa2_uq0 vssd1_uq1
XFILLER_3_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1828_A wire1828/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1902 wire1903/X vssd vssd vccd vccd _615_/B sky130_fd_sc_hd__buf_6
XFILLER_28_1583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1913 wire1914/X vssd vssd vccd vccd wire1913/X sky130_fd_sc_hd__buf_6
XFILLER_28_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1666 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1924 wire1924/A vssd vssd vccd vccd wire1924/X sky130_fd_sc_hd__buf_6
Xwire1935 wire1936/X vssd vssd vccd vccd wire1935/X sky130_fd_sc_hd__buf_6
XFILLER_3_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1946 wire1947/X vssd vssd vccd vccd wire1946/X sky130_fd_sc_hd__buf_6
XTAP_3202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1957 wire1958/X vssd vssd vccd vccd _595_/B sky130_fd_sc_hd__buf_6
XFILLER_19_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1968 wire1968/A vssd vssd vccd vccd wire1968/X sky130_fd_sc_hd__buf_6
XFILLER_18_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1979 wire1980/X vssd vssd vccd vccd _584_/B sky130_fd_sc_hd__buf_6
XTAP_3235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input127_A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2044_A wire2044/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_501_ _501_/A _501_/B vssd vssd vccd vccd _501_/X sky130_fd_sc_hd__and2_4
XANTENNA_202 _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_213 _230_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_224 _205_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_246 _539_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 _480_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_432_ _560_/A _432_/B _432_/C vssd vssd vccd vccd _432_/X sky130_fd_sc_hd__and3b_4
XFILLER_26_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_268 _544_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_279 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_363_ _363_/A _363_/B vssd vssd vccd vccd _363_/X sky130_fd_sc_hd__and2_2
XTAP_1888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input92_A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_294_ _294_/A _294_/B vssd vssd vccd vccd _294_/X sky130_fd_sc_hd__and2_4
XFILLER_48_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[8\] mprj_dat_i_user[8] max_length1311/X vssd vssd vccd vccd _122_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output513_A wire1143/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1144_A _370_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1409_A wire1410/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] _188_/X vssd vssd vccd vccd _008_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1680_A wire1681/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1778_A wire1779/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__304__A _304_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1945_A wire1946/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput467 wire1063/X vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__buf_8
Xoutput478 _482_/X vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__buf_8
XFILLER_42_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput489 _492_/X vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__buf_8
XFILLER_9_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1209 wire1210/X vssd vssd vccd vccd wire1209/X sky130_fd_sc_hd__buf_6
XFILLER_0_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__A_N _618_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__214__A _214_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4382 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2161_A wire2161/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input244_A la_iena_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1710 wire1710/A vssd vssd vccd vccd _358_/A sky130_fd_sc_hd__buf_6
XFILLER_5_3797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1721 wire1722/X vssd vssd vccd vccd wire1721/X sky130_fd_sc_hd__buf_6
XFILLER_1_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1732 wire1733/X vssd vssd vccd vccd _291_/A sky130_fd_sc_hd__buf_6
XFILLER_46_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1743 wire1743/A vssd vssd vccd vccd wire1743/X sky130_fd_sc_hd__buf_6
XFILLER_19_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1754 wire1754/A vssd vssd vccd vccd wire1754/X sky130_fd_sc_hd__buf_6
XTAP_3010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input411_A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1765 wire1766/X vssd vssd vccd vccd _276_/A sky130_fd_sc_hd__buf_6
XTAP_3021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1776 wire1776/A vssd vssd vccd vccd wire1776/X sky130_fd_sc_hd__buf_6
XFILLER_37_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1787 wire1788/X vssd vssd vccd vccd _264_/A sky130_fd_sc_hd__buf_6
XFILLER_19_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1798 wire1798/A vssd vssd vccd vccd _258_/A sky130_fd_sc_hd__buf_6
XTAP_3054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ _415_/A_N _415_/B _415_/C vssd vssd vccd vccd _415_/X sky130_fd_sc_hd__and3b_4
XTAP_2397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_346_ _346_/A _346_/B vssd vssd vccd vccd _346_/X sky130_fd_sc_hd__and2_4
XFILLER_30_957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_277_ _277_/A _277_/B vssd vssd vccd vccd _277_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output463_A wire1145/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_880 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1261_A _320_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1359_A wire1359/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1526_A wire1526/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1895_A wire1896/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__034__A _034_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1170 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1006 _550_/X vssd vssd vccd vccd wire1006/X sky130_fd_sc_hd__buf_6
Xwire1017 _539_/X vssd vssd vccd vccd wire1017/X sky130_fd_sc_hd__buf_6
Xwire1028 _521_/X vssd vssd vccd vccd wire1028/X sky130_fd_sc_hd__buf_6
XFILLER_38_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1039 _510_/X vssd vssd vccd vccd wire1039/X sky130_fd_sc_hd__buf_6
XFILLER_28_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1903 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__209__A _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_200_ _200_/A _200_/B vssd vssd vccd vccd _200_/X sky130_fd_sc_hd__and2_4
XFILLER_51_2837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2007_A wire2008/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_131_ _131_/A vssd vssd vccd vccd _131_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_36_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input194_A la_iena_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_062_ _062_/A vssd vssd vccd vccd _062_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__386__A_N _514_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input361_A la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input459_A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input55_A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4010 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__598__B _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1540 wire1540/A vssd vssd vccd vccd _574_/A sky130_fd_sc_hd__buf_8
XFILLER_24_1052 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1551 wire1551/A vssd vssd vccd vccd _563_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1573 input31/X vssd vssd vccd vccd _493_/C sky130_fd_sc_hd__buf_6
XFILLER_19_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1584 wire1584/A vssd vssd vccd vccd _619_/A sky130_fd_sc_hd__buf_6
Xwire1595 wire1595/A vssd vssd vccd vccd _608_/A sky130_fd_sc_hd__buf_6
XFILLER_1_2768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__119__A _119_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3146 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output580_A wire1076/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1107_A _406_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_329_ _329_/A _329_/B vssd vssd vccd vccd _329_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output845_A _596_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1476_A wire1476/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] wire1322/X vssd vssd vccd vccd wire965/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_45_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1643_A wire1644/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__301__B _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1908_A wire1909/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__211__B _211_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_810 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2124_A wire2125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input207_A la_iena_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_114_ _114_/A vssd vssd vccd vccd _114_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_045_ _045_/A vssd vssd vccd vccd _045_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_2375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2060 wire2061/X vssd vssd vccd vccd _499_/B sky130_fd_sc_hd__buf_6
Xwire2071 wire2072/X vssd vssd vccd vccd wire2071/X sky130_fd_sc_hd__buf_6
XFILLER_1_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2082 wire2083/X vssd vssd vccd vccd _491_/B sky130_fd_sc_hd__buf_6
XFILLER_38_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2093 wire2093/A vssd vssd vccd vccd wire2093/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1057_A _478_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__401__A_N _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1370 wire1370/A vssd vssd vccd vccd _358_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1381 wire1382/X vssd vssd vccd vccd _351_/B sky130_fd_sc_hd__buf_6
XFILLER_53_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1392 wire1393/X vssd vssd vccd vccd wire1392/X sky130_fd_sc_hd__buf_6
XFILLER_1_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1224_A wire1225/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output795_A wire1005/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[20\] mprj_dat_i_user[20] _294_/X vssd vssd vccd vccd _134_/A sky130_fd_sc_hd__nand2_2
XFILLER_50_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1760_A wire1760/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1858_A wire1858/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__312__A _312_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__206__B _206_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3746 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2074_A wire2075/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input157_A la_iena_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput301 la_oenb_mprj[21] vssd vssd vccd vccd _518_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__424__A_N _552_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput312 la_oenb_mprj[31] vssd vssd vccd vccd _400_/A_N sky130_fd_sc_hd__buf_6
XFILLER_0_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput323 la_oenb_mprj[41] vssd vssd vccd vccd _538_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput334 la_oenb_mprj[51] vssd vssd vccd vccd _420_/A_N sky130_fd_sc_hd__buf_6
XFILLER_2_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput345 la_oenb_mprj[61] vssd vssd vccd vccd _558_/A sky130_fd_sc_hd__clkbuf_4
Xinput356 la_oenb_mprj[71] vssd vssd vccd vccd wire1546/A sky130_fd_sc_hd__buf_6
Xinput367 la_oenb_mprj[81] vssd vssd vccd vccd wire1536/A sky130_fd_sc_hd__buf_6
XANTENNA_input324_A la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput378 la_oenb_mprj[91] vssd vssd vccd vccd _588_/A sky130_fd_sc_hd__buf_6
XFILLER_40_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput389 mprj_adr_o_core[10] vssd vssd vccd vccd wire1521/A sky130_fd_sc_hd__buf_6
XFILLER_53_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input18_A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_594_ _594_/A _594_/B vssd vssd vccd vccd _594_/X sky130_fd_sc_hd__and2_4
XFILLER_16_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1774 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_5 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput808 _562_/X vssd vssd vccd vccd la_oenb_core[65] sky130_fd_sc_hd__buf_8
Xoutput819 _572_/X vssd vssd vccd vccd la_oenb_core[75] sky130_fd_sc_hd__buf_8
X_028_ _028_/A vssd vssd vccd vccd _028_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output543_A wire1084/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__132__A _132_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1174_A wire1175/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3234 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output808_A _562_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1439_A wire1440/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] _218_/X vssd vssd vccd vccd _038_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_48_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4362 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__307__A _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1975_A wire1975/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__447__A_N _575_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_142 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__217__A _217_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input274_A la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2191_A wire2191/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input441_A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput120 la_data_out_mprj[8] vssd vssd vccd vccd _377_/C sky130_fd_sc_hd__clkbuf_4
Xinput131 la_data_out_mprj[9] vssd vssd vccd vccd _378_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_1_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput142 la_iena_mprj[109] vssd vssd vccd vccd _272_/B sky130_fd_sc_hd__clkbuf_4
Xinput153 la_iena_mprj[119] vssd vssd vccd vccd _282_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput164 la_iena_mprj[13] vssd vssd vccd vccd _176_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 la_iena_mprj[23] vssd vssd vccd vccd wire1615/A sky130_fd_sc_hd__buf_6
XTAP_4652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 la_iena_mprj[33] vssd vssd vccd vccd _196_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput197 la_iena_mprj[43] vssd vssd vccd vccd _206_/B sky130_fd_sc_hd__buf_4
XTAP_4674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3314 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_577_ _577_/A _577_/B vssd vssd vccd vccd _577_/X sky130_fd_sc_hd__and2_4
XFILLER_32_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output493_A _496_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__127__A _127_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output660_A _030_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output758_A wire1052/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1291_A wire1292/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput605 _095_/Y vssd vssd vccd vccd la_data_in_mprj[112] sky130_fd_sc_hd__buf_8
XFILLER_9_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1389_A wire1390/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput616 _105_/Y vssd vssd vccd vccd la_data_in_mprj[122] sky130_fd_sc_hd__buf_8
XFILLER_29_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput627 _000_/Y vssd vssd vccd vccd la_data_in_mprj[17] sky130_fd_sc_hd__buf_8
XFILLER_42_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput638 _010_/Y vssd vssd vccd vccd la_data_in_mprj[27] sky130_fd_sc_hd__buf_8
XFILLER_29_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output925_A wire1190/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput649 _020_/Y vssd vssd vccd vccd la_data_in_mprj[37] sky130_fd_sc_hd__buf_8
XFILLER_42_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1723_A wire1724/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__037__A _037_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_B _197_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1903 wire1904/X vssd vssd vccd vccd wire1903/X sky130_fd_sc_hd__buf_6
XANTENNA__500__A _500_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1914 wire1914/A vssd vssd vccd vccd wire1914/X sky130_fd_sc_hd__buf_6
XFILLER_8_1678 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1925 wire1926/X vssd vssd vccd vccd _608_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1936 wire1936/A vssd vssd vccd vccd wire1936/X sky130_fd_sc_hd__buf_6
XFILLER_6_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1947 wire1947/A vssd vssd vccd vccd wire1947/X sky130_fd_sc_hd__buf_6
XTAP_3203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1958 wire1958/A vssd vssd vccd vccd wire1958/X sky130_fd_sc_hd__buf_6
XTAP_3214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1969 wire1970/X vssd vssd vccd vccd _591_/B sky130_fd_sc_hd__buf_6
XTAP_3225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_500_ _500_/A _500_/B vssd vssd vccd vccd _500_/X sky130_fd_sc_hd__and2_4
XFILLER_19_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 _230_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_225 _205_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2037_A wire2038/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_431_ _559_/A _431_/B _431_/C vssd vssd vccd vccd _431_/X sky130_fd_sc_hd__and3b_2
XTAP_2557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_247 _539_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 _480_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_362_ _362_/A _362_/B vssd vssd vccd vccd _362_/X sky130_fd_sc_hd__and2_2
XTAP_1878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_293_ _293_/A _293_/B vssd vssd vccd vccd _293_/X sky130_fd_sc_hd__and2_1
XFILLER_35_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input391_A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input85_A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_856 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output506_A wire1121/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1137_A _377_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1304_A wire1305/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output875_A _310_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] _181_/X vssd vssd vccd vccd _001_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_31_1920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1673_A wire1673/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[16\]_B _179_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[100\]_B _263_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__304__B _304_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1840_A wire1840/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput468 wire1062/X vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__buf_8
XANTENNA_wire1938_A wire1938/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput479 _483_/X vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__buf_8
XFILLER_9_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__320__A _320_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__214__B _214_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_826 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4394 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__230__A _230_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1700 wire1701/X vssd vssd vccd vccd _364_/A sky130_fd_sc_hd__buf_6
Xwire1711 wire1711/A vssd vssd vccd vccd _357_/A sky130_fd_sc_hd__buf_6
Xwire1722 wire1722/A vssd vssd vccd vccd wire1722/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2154_A wire2154/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input237_A la_iena_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1733 wire1734/X vssd vssd vccd vccd wire1733/X sky130_fd_sc_hd__buf_6
Xwire1744 wire1745/X vssd vssd vccd vccd _286_/A sky130_fd_sc_hd__buf_6
XFILLER_46_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1755 wire1756/X vssd vssd vccd vccd _281_/A sky130_fd_sc_hd__buf_6
Xwire1766 wire1766/A vssd vssd vccd vccd wire1766/X sky130_fd_sc_hd__buf_6
XTAP_3011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1777 wire1777/A vssd vssd vccd vccd _270_/A sky130_fd_sc_hd__buf_6
XTAP_3033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1788 wire1788/A vssd vssd vccd vccd wire1788/X sky130_fd_sc_hd__buf_6
XFILLER_41_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1799 wire1799/A vssd vssd vccd vccd _257_/A sky130_fd_sc_hd__buf_6
XTAP_3055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input404_A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ _542_/A _414_/B _414_/C vssd vssd vccd vccd _414_/X sky130_fd_sc_hd__and3b_4
XFILLER_19_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_966 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ _345_/A _345_/B vssd vssd vccd vccd _345_/X sky130_fd_sc_hd__and2_2
XFILLER_50_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2952 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_276_ _276_/A _276_/B vssd vssd vccd vccd _276_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1087_A wire1088/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__140__A _140_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1254_A wire1255/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2530 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1421_A wire1421/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1519_A wire1519/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1888_A wire1888/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__315__A _315_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1182 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__050__A _050_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1007 wire1008/X vssd vssd vccd vccd wire1007/X sky130_fd_sc_hd__buf_6
XFILLER_5_1604 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1018 _538_/X vssd vssd vccd vccd wire1018/X sky130_fd_sc_hd__buf_6
Xwire1029 _520_/X vssd vssd vccd vccd wire1029/X sky130_fd_sc_hd__buf_6
XFILLER_0_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1915 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__209__B _209_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_582 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_130_ _130_/A vssd vssd vccd vccd _130_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_3394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__225__A _225_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_061_ _061_/A vssd vssd vccd vccd _061_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_4423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input187_A la_iena_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input354_A la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input48_A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1530 wire1530/A vssd vssd vccd vccd _584_/A sky130_fd_sc_hd__buf_6
XFILLER_21_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1541 wire1541/A vssd vssd vccd vccd _573_/A sky130_fd_sc_hd__buf_8
XFILLER_47_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1552 wire1552/A vssd vssd vccd vccd _562_/A sky130_fd_sc_hd__buf_6
XFILLER_46_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1563 _415_/A_N vssd vssd vccd vccd _543_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1574 wire1574/A vssd vssd vccd vccd _526_/A sky130_fd_sc_hd__buf_6
XFILLER_38_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1585 wire1585/A vssd vssd vccd vccd _618_/A sky130_fd_sc_hd__buf_6
XFILLER_47_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1596 _479_/A_N vssd vssd vccd vccd _607_/A sky130_fd_sc_hd__buf_4
XFILLER_46_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1002_A wire1003/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_328_ _328_/A _328_/B vssd vssd vccd vccd _328_/X sky130_fd_sc_hd__and2_4
XFILLER_15_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output573_A _453_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__135__A _135_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_259_ _259_/A _259_/B vssd vssd vccd vccd _259_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output740_A _616_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output838_A _589_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1371_A wire1371/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1469_A wire1470/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1014 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__480__A_N _608_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] wire1329/X vssd vssd vccd vccd wire972/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1222 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__045__A _045_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_822 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_538 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input102_A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2117_A wire2118/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_113_ _113_/A vssd vssd vccd vccd _113_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_044_ _044_/A vssd vssd vccd vccd _044_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2050 wire2050/A vssd vssd vccd vccd wire2050/X sky130_fd_sc_hd__buf_6
XFILLER_43_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2061 wire2061/A vssd vssd vccd vccd wire2061/X sky130_fd_sc_hd__buf_6
Xwire2072 wire2072/A vssd vssd vccd vccd wire2072/X sky130_fd_sc_hd__buf_6
Xwire2083 wire2084/X vssd vssd vccd vccd wire2083/X sky130_fd_sc_hd__buf_6
Xwire2094 wire2095/X vssd vssd vccd vccd _487_/B sky130_fd_sc_hd__buf_6
XFILLER_47_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1360 wire1361/X vssd vssd vccd vccd _339_/B sky130_fd_sc_hd__buf_6
Xwire1371 wire1371/A vssd vssd vccd vccd _357_/B sky130_fd_sc_hd__buf_6
Xwire1382 wire1382/A vssd vssd vccd vccd wire1382/X sky130_fd_sc_hd__buf_6
Xwire1393 wire1393/A vssd vssd vccd vccd wire1393/X sky130_fd_sc_hd__buf_6
XFILLER_19_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1217_A wire1218/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output690_A _057_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output788_A _544_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output955_A wire1307/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[13\] mprj_dat_i_user[13] max_length1311/X vssd vssd vccd vccd
+ _127_/A sky130_fd_sc_hd__nand2_2
XFILLER_28_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1753_A wire1754/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__312__B _312_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[1\]_A mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1920_A wire1921/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] _274_/X vssd vssd vccd vccd wire988/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_6_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__376__A_N _504_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput302 la_oenb_mprj[22] vssd vssd vccd vccd _519_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput313 la_oenb_mprj[32] vssd vssd vccd vccd wire1570/A sky130_fd_sc_hd__buf_6
XFILLER_2_4255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput324 la_oenb_mprj[42] vssd vssd vccd vccd _539_/A sky130_fd_sc_hd__buf_4
XFILLER_40_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput335 la_oenb_mprj[52] vssd vssd vccd vccd _549_/A sky130_fd_sc_hd__buf_4
XANTENNA_wire2067_A wire2068/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput346 la_oenb_mprj[62] vssd vssd vccd vccd wire1555/A sky130_fd_sc_hd__buf_6
Xinput357 la_oenb_mprj[72] vssd vssd vccd vccd wire1545/A sky130_fd_sc_hd__buf_6
XFILLER_2_3565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput368 la_oenb_mprj[82] vssd vssd vccd vccd wire1535/A sky130_fd_sc_hd__buf_6
XFILLER_5_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput379 la_oenb_mprj[92] vssd vssd vccd vccd _589_/A sky130_fd_sc_hd__buf_6
XFILLER_29_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input317_A la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_593_ _593_/A _593_/B vssd vssd vccd vccd _593_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_6 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput809 _563_/X vssd vssd vccd vccd la_oenb_core[66] sky130_fd_sc_hd__buf_8
X_027_ _027_/A vssd vssd vccd vccd _027_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_2924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output536_A wire1093/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1167_A wire1168/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__399__A_N _527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1190 wire1191/X vssd vssd vccd vccd wire1190/X sky130_fd_sc_hd__buf_8
XFILLER_39_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] _211_/X vssd vssd vccd vccd _031_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_34_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1501_A wire1502/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__307__B _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1870_A wire1870/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1968_A wire1968/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__323__A _323_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4230 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__233__A _233_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2184_A wire2185/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input267_A la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input434_A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput110 la_data_out_mprj[80] vssd vssd vccd vccd wire1624/A sky130_fd_sc_hd__buf_6
Xinput121 la_data_out_mprj[90] vssd vssd vccd vccd _459_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_input30_A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput132 la_iena_mprj[0] vssd vssd vccd vccd _625_/B sky130_fd_sc_hd__clkbuf_4
Xinput143 la_iena_mprj[10] vssd vssd vccd vccd _173_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput154 la_iena_mprj[11] vssd vssd vccd vccd _174_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput165 la_iena_mprj[14] vssd vssd vccd vccd _177_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput176 la_iena_mprj[24] vssd vssd vccd vccd wire1614/A sky130_fd_sc_hd__buf_6
XTAP_4653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput187 la_iena_mprj[34] vssd vssd vccd vccd _197_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput198 la_iena_mprj[44] vssd vssd vccd vccd _207_/B sky130_fd_sc_hd__buf_4
XFILLER_36_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_576_ _576_/A _576_/B vssd vssd vccd vccd _576_/X sky130_fd_sc_hd__and2_4
XFILLER_16_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output486_A _489_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output653_A _023_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput606 _096_/Y vssd vssd vccd vccd la_data_in_mprj[113] sky130_fd_sc_hd__buf_8
XANTENNA__143__A _143_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput617 _106_/Y vssd vssd vccd vccd la_data_in_mprj[123] sky130_fd_sc_hd__buf_8
XANTENNA_wire1284_A wire1285/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput628 _001_/Y vssd vssd vccd vccd la_data_in_mprj[18] sky130_fd_sc_hd__buf_8
Xoutput639 _011_/Y vssd vssd vccd vccd la_data_in_mprj[28] sky130_fd_sc_hd__buf_8
XFILLER_25_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output820_A _573_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output918_A wire1211/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1451_A wire1451/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1716_A wire1716/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__414__A_N _542_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__053__A _053_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1904 wire1904/A vssd vssd vccd vccd wire1904/X sky130_fd_sc_hd__buf_6
XFILLER_8_1657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__500__B _500_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1915 wire1916/X vssd vssd vccd vccd _611_/B sky130_fd_sc_hd__buf_6
Xwire1926 wire1927/X vssd vssd vccd vccd wire1926/X sky130_fd_sc_hd__buf_6
XTAP_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1937 wire1938/X vssd vssd vccd vccd _604_/B sky130_fd_sc_hd__buf_6
Xwire1948 wire1949/X vssd vssd vccd vccd _599_/B sky130_fd_sc_hd__buf_6
XTAP_3204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1959 wire1960/X vssd vssd vccd vccd _297_/A sky130_fd_sc_hd__buf_6
XTAP_3215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 _205_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_430_ _558_/A _430_/B _430_/C vssd vssd vccd vccd _430_/X sky130_fd_sc_hd__and3b_4
XANTENNA_248 _539_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_259 _480_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__228__A _228_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_361_ _361_/A _361_/B vssd vssd vccd vccd _361_/X sky130_fd_sc_hd__and2_2
XFILLER_13_3212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_292_ _292_/A _292_/B vssd vssd vccd vccd _292_/X sky130_fd_sc_hd__and2_1
XFILLER_42_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input384_A la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input78_A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__410__B _410_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1032_A _517_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__437__A_N _565_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__138__A _138_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_559_ _559_/A _559_/B vssd vssd vccd vccd _559_/X sky130_fd_sc_hd__and2_4
XFILLER_14_2308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output868_A _333_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1499_A wire1500/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1666_A wire1667/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput469 wire1061/X vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__buf_8
XANTENNA__601__A _601_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1833_A wire1834/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__320__B _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__048__A _048_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4362 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__511__A _511_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__230__B _230_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1701 wire1701/A vssd vssd vccd vccd wire1701/X sky130_fd_sc_hd__buf_6
XFILLER_43_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1712 wire1712/A vssd vssd vccd vccd _356_/A sky130_fd_sc_hd__buf_6
Xwire1723 wire1724/X vssd vssd vccd vccd wire1723/X sky130_fd_sc_hd__buf_6
XFILLER_24_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1734 wire1734/A vssd vssd vccd vccd wire1734/X sky130_fd_sc_hd__buf_6
Xwire1745 wire1745/A vssd vssd vccd vccd wire1745/X sky130_fd_sc_hd__buf_6
XTAP_3001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input132_A la_iena_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1756 wire1756/A vssd vssd vccd vccd wire1756/X sky130_fd_sc_hd__buf_6
XFILLER_46_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1767 wire1768/X vssd vssd vccd vccd _275_/A sky130_fd_sc_hd__buf_6
XANTENNA_wire2147_A wire2148/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1778 wire1779/X vssd vssd vccd vccd _269_/A sky130_fd_sc_hd__buf_6
XTAP_3034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1789 wire1790/X vssd vssd vccd vccd _263_/A sky130_fd_sc_hd__buf_6
XFILLER_19_4144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_413_ _541_/A _413_/B _413_/C vssd vssd vccd vccd _413_/X sky130_fd_sc_hd__and3b_4
XTAP_2377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ _344_/A _344_/B vssd vssd vccd vccd _344_/X sky130_fd_sc_hd__and2_2
XFILLER_53_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_3930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_275_ _275_/A _275_/B vssd vssd vccd vccd _275_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2964 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__405__B _405_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output616_A _105_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1247_A wire1248/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1414_A wire1415/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] _193_/X vssd vssd vccd vccd _013_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_33_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__315__B _315_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1950_A wire1951/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__331__A _331_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1008 _549_/X vssd vssd vccd vccd wire1008/X sky130_fd_sc_hd__buf_6
Xwire1019 _536_/X vssd vssd vccd vccd wire1019/X sky130_fd_sc_hd__buf_6
XFILLER_5_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_A mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__506__A _506_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__225__B _225_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_060_ _060_/A vssd vssd vccd vccd _060_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2097_A wire2098/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__241__A _241_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input347_A la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1520 wire1521/X vssd vssd vccd vccd _315_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1531 wire1531/A vssd vssd vccd vccd _583_/A sky130_fd_sc_hd__buf_6
XFILLER_19_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1542 wire1542/A vssd vssd vccd vccd _572_/A sky130_fd_sc_hd__buf_8
XFILLER_21_2643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1553 wire1553/A vssd vssd vccd vccd _561_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1564 _412_/A_N vssd vssd vccd vccd _540_/A sky130_fd_sc_hd__buf_4
XFILLER_24_1076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1575 wire1575/A vssd vssd vccd vccd _524_/A sky130_fd_sc_hd__buf_6
Xwire1586 wire1586/A vssd vssd vccd vccd _617_/A sky130_fd_sc_hd__buf_6
Xwire1597 _478_/A_N vssd vssd vccd vccd _606_/A sky130_fd_sc_hd__buf_6
XFILLER_47_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_327_ _327_/A _327_/B vssd vssd vccd vccd _327_/X sky130_fd_sc_hd__and2_4
XFILLER_15_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_258_ _258_/A _258_/B vssd vssd vccd vccd _258_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output566_A _447_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_189_ _189_/A _189_/B vssd vssd vccd vccd _189_/X sky130_fd_sc_hd__and2_2
XFILLER_45_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output733_A _609_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1364_A wire1364/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2576 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] _241_/X vssd vssd vccd vccd wire978/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_6_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1531_A wire1531/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1629_A wire1629/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1998_A wire1999/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__326__A _326_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1234 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__061__A _061_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1779 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2012_A wire2013/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__236__A _236_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input297_A la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_112_ _112_/A vssd vssd vccd vccd _112_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_043_ _043_/A vssd vssd vccd vccd _043_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input60_A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__402__C _402_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2040 wire2041/X vssd vssd vccd vccd _511_/B sky130_fd_sc_hd__buf_6
Xwire2051 wire2051/A vssd vssd vccd vccd _505_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2062 wire2063/X vssd vssd vccd vccd _498_/B sky130_fd_sc_hd__buf_6
Xwire2073 wire2074/X vssd vssd vccd vccd _494_/B sky130_fd_sc_hd__buf_6
XFILLER_19_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2084 wire2084/A vssd vssd vccd vccd wire2084/X sky130_fd_sc_hd__buf_6
XFILLER_19_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1350 wire1351/X vssd vssd vccd vccd _343_/B sky130_fd_sc_hd__buf_6
Xwire2095 wire2096/X vssd vssd vccd vccd wire2095/X sky130_fd_sc_hd__buf_6
Xwire1361 wire1361/A vssd vssd vccd vccd wire1361/X sky130_fd_sc_hd__buf_6
XFILLER_47_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1372 wire1373/X vssd vssd vccd vccd _338_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1383 wire1384/X vssd vssd vccd vccd _350_/B sky130_fd_sc_hd__buf_6
XFILLER_46_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1394 wire1395/X vssd vssd vccd vccd _298_/B sky130_fd_sc_hd__buf_6
XFILLER_19_377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_870 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output683_A _051_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output850_A wire1268/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output948_A wire1280/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1746_A wire1747/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_B max_length1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1913_A wire1914/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] _267_/X vssd vssd vccd vccd _087_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_17_3700 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__056__A _056_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__503__B _503_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput303 la_oenb_mprj[23] vssd vssd vccd vccd _520_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput314 la_oenb_mprj[33] vssd vssd vccd vccd _530_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput325 la_oenb_mprj[43] vssd vssd vccd vccd _412_/A_N sky130_fd_sc_hd__buf_6
Xinput336 la_oenb_mprj[53] vssd vssd vccd vccd _550_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput347 la_oenb_mprj[63] vssd vssd vccd vccd wire1554/A sky130_fd_sc_hd__buf_6
XFILLER_22_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput358 la_oenb_mprj[73] vssd vssd vccd vccd wire1544/A sky130_fd_sc_hd__buf_6
Xinput369 la_oenb_mprj[83] vssd vssd vccd vccd wire1534/A sky130_fd_sc_hd__buf_6
XFILLER_2_3588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input212_A la_iena_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_592_ _592_/A _592_/B vssd vssd vccd vccd _592_/X sky130_fd_sc_hd__and2_4
XFILLER_43_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__470__A_N _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_7 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_026_ _026_/A vssd vssd vccd vccd _026_/Y sky130_fd_sc_hd__inv_2
XANTENNA__413__B _413_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output529_A wire1100/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1062_A _473_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1180 wire1181/X vssd vssd vccd vccd wire1180/X sky130_fd_sc_hd__buf_6
Xwire1191 wire1192/X vssd vssd vccd vccd wire1191/X sky130_fd_sc_hd__buf_6
XFILLER_1_3098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1327_A _250_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1696_A wire1697/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1362 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__604__A _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1863_A wire1864/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__323__B _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__493__A_N _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__514__A _514_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__233__B _233_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input162_A la_iena_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2177_A wire2178/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput100 la_data_out_mprj[71] vssd vssd vccd vccd wire1633/A sky130_fd_sc_hd__buf_6
XFILLER_2_4042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput111 la_data_out_mprj[81] vssd vssd vccd vccd wire1623/A sky130_fd_sc_hd__buf_6
XFILLER_44_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput122 la_data_out_mprj[91] vssd vssd vccd vccd _460_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput133 la_iena_mprj[100] vssd vssd vccd vccd _263_/B sky130_fd_sc_hd__buf_4
XFILLER_23_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput144 la_iena_mprj[110] vssd vssd vccd vccd _273_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input427_A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput155 la_iena_mprj[120] vssd vssd vccd vccd _283_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 la_iena_mprj[15] vssd vssd vccd vccd _178_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input23_A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput177 la_iena_mprj[25] vssd vssd vccd vccd wire1613/A sky130_fd_sc_hd__buf_6
XTAP_4654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 la_iena_mprj[35] vssd vssd vccd vccd _198_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput199 la_iena_mprj[45] vssd vssd vccd vccd _208_/B sky130_fd_sc_hd__buf_4
XFILLER_29_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_575_ _575_/A _575_/B vssd vssd vccd vccd _575_/X sky130_fd_sc_hd__and2_4
XFILLER_44_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__408__B _408_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output479_A _483_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_29_4157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput607 _097_/Y vssd vssd vccd vccd la_data_in_mprj[114] sky130_fd_sc_hd__buf_8
XFILLER_9_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput618 _107_/Y vssd vssd vccd vccd la_data_in_mprj[124] sky130_fd_sc_hd__buf_8
Xoutput629 _002_/Y vssd vssd vccd vccd la_data_in_mprj[19] sky130_fd_sc_hd__buf_8
XFILLER_29_2733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output646_A _017_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_009_ _009_/A vssd vssd vccd vccd _009_/Y sky130_fd_sc_hd__inv_4
XFILLER_46_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1277_A _312_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output813_A wire1047/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1444_A wire1445/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] _223_/X vssd vssd vccd vccd _043_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_23_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1709_A wire1709/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__318__B _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1980_A wire1980/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4194 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__334__A _334_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_max_length1311_A _294_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1905 wire1906/X vssd vssd vccd vccd _614_/B sky130_fd_sc_hd__buf_6
XTAP_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1916 wire1917/X vssd vssd vccd vccd wire1916/X sky130_fd_sc_hd__buf_6
XFILLER_28_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1927 wire1927/A vssd vssd vccd vccd wire1927/X sky130_fd_sc_hd__buf_6
XFILLER_41_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1938 wire1938/A vssd vssd vccd vccd wire1938/X sky130_fd_sc_hd__buf_6
XTAP_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1949 wire1949/A vssd vssd vccd vccd wire1949/X sky130_fd_sc_hd__buf_6
XFILLER_19_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_205 _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_216 _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_227 _204_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__509__A _509_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_249 _539_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__228__B _228_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ _360_/A _360_/B vssd vssd vccd vccd _360_/X sky130_fd_sc_hd__and2_2
XFILLER_17_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_291_ _291_/A _291_/B vssd vssd vccd vccd _291_/X sky130_fd_sc_hd__and2_1
XFILLER_52_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__244__A _244_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__389__A_N _517_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input377_A la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__410__C _410_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_558_ _558_/A _558_/B vssd vssd vccd vccd _558_/X sky130_fd_sc_hd__and2_2
XANTENNA_wire1025_A _525_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output596_A _087_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_489_ _617_/A _489_/B _489_/C vssd vssd vccd vccd _489_/X sky130_fd_sc_hd__and3b_4
XFILLER_20_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output763_A wire1028/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1394_A wire1395/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output930_A wire1170/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1561_A wire1561/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1659_A wire1660/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__601__B _601_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1826_A wire1826/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__329__A _329_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__064__A _064_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput960 _295_/X vssd vssd vccd vccd user_reset sky130_fd_sc_hd__buf_8
XFILLER_9_3881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__511__B _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1702 wire1703/X vssd vssd vccd vccd _363_/A sky130_fd_sc_hd__buf_6
XFILLER_5_3789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1713 wire1713/A vssd vssd vccd vccd _355_/A sky130_fd_sc_hd__buf_6
XFILLER_8_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1724 wire1725/X vssd vssd vccd vccd wire1724/X sky130_fd_sc_hd__buf_6
XFILLER_1_2908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1735 wire1736/X vssd vssd vccd vccd _290_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1746 wire1747/X vssd vssd vccd vccd _285_/A sky130_fd_sc_hd__buf_6
XTAP_3002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1757 wire1758/X vssd vssd vccd vccd _280_/A sky130_fd_sc_hd__buf_6
Xwire1768 wire1768/A vssd vssd vccd vccd wire1768/X sky130_fd_sc_hd__buf_6
XTAP_3013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1779 wire1779/A vssd vssd vccd vccd wire1779/X sky130_fd_sc_hd__buf_6
XTAP_3035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2042_A wire2043/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input125_A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__239__A _239_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_412_ _412_/A_N _412_/B _412_/C vssd vssd vccd vccd _412_/X sky130_fd_sc_hd__and3b_4
XTAP_2367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_343_ _343_/A _343_/B vssd vssd vccd vccd _343_/X sky130_fd_sc_hd__and2_2
XFILLER_52_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input90_A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_274_ _274_/A _274_/B vssd vssd vccd vccd _274_/X sky130_fd_sc_hd__and2_4
XFILLER_52_2391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__405__C _405_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[6\] mprj_dat_i_user[6] max_length1311/X vssd vssd vccd vccd _120_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_10_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__421__B _421_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__404__A_N _532_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output511_A wire1116/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output609_A _099_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1142_A _372_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1407_A wire1408/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output880_A wire1306/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] _186_/X vssd vssd vccd vccd _006_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_18_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1776_A wire1776/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__612__A _612_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1943_A wire1944/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__331__B _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3802 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1009 wire1010/X vssd vssd vccd vccd wire1009/X sky130_fd_sc_hd__buf_6
XFILLER_20_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__059__A _059_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_B max_length1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__506__B _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__522__A _522_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__427__A_N _555_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__241__B _241_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2200 wire2200/A vssd vssd vccd vccd _306_/A sky130_fd_sc_hd__buf_6
Xoutput790 wire1011/X vssd vssd vccd vccd la_oenb_core[49] sky130_fd_sc_hd__buf_8
XFILLER_1_4118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input242_A la_iena_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3334 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1510 wire1511/X vssd vssd vccd vccd wire1510/X sky130_fd_sc_hd__buf_6
XFILLER_1_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1521 wire1521/A vssd vssd vccd vccd wire1521/X sky130_fd_sc_hd__buf_6
Xwire1532 wire1532/A vssd vssd vccd vccd _582_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1543 wire1543/A vssd vssd vccd vccd _571_/A sky130_fd_sc_hd__buf_6
XFILLER_48_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1554 wire1554/A vssd vssd vccd vccd _560_/A sky130_fd_sc_hd__buf_6
Xwire1565 _409_/A_N vssd vssd vccd vccd _537_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1576 wire1577/X vssd vssd vccd vccd _295_/A_N sky130_fd_sc_hd__buf_6
XFILLER_38_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1587 wire1587/A vssd vssd vccd vccd _616_/A sky130_fd_sc_hd__buf_6
XFILLER_0_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1598 input27/X vssd vssd vccd vccd _489_/C sky130_fd_sc_hd__buf_4
XFILLER_21_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_326_ _326_/A _326_/B vssd vssd vccd vccd _326_/X sky130_fd_sc_hd__and2_4
XFILLER_9_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__416__B _416_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_257_ _257_/A _257_/B vssd vssd vccd vccd _257_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_188_ _188_/A _188_/B vssd vssd vccd vccd _188_/X sky130_fd_sc_hd__and2_2
XANTENNA_output559_A _440_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1092_A _420_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output726_A _603_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1357_A wire1357/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1524_A wire1525/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__607__A _607_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1893_A wire1894/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__326__B _326_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire977_A wire977/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[91\]_B wire1323/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__342__A _342_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__517__A _517_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__236__B _236_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2005_A wire2006/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_111_ _111_/A vssd vssd vccd vccd _111_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_2470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input192_A la_iena_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_042_ _042_/A vssd vssd vccd vccd _042_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__252__A _252_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input457_A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input53_A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2030 wire2030/A vssd vssd vccd vccd _520_/B sky130_fd_sc_hd__buf_6
Xwire2041 wire2041/A vssd vssd vccd vccd wire2041/X sky130_fd_sc_hd__buf_6
Xwire2052 wire2052/A vssd vssd vccd vccd _504_/B sky130_fd_sc_hd__buf_6
XFILLER_38_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2063 wire2063/A vssd vssd vccd vccd wire2063/X sky130_fd_sc_hd__buf_6
Xwire2074 wire2075/X vssd vssd vccd vccd wire2074/X sky130_fd_sc_hd__buf_6
XFILLER_21_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1340 input85/X vssd vssd vccd vccd _427_/C sky130_fd_sc_hd__buf_6
Xwire2085 wire2086/X vssd vssd vccd vccd _490_/B sky130_fd_sc_hd__buf_6
Xwire1351 wire1351/A vssd vssd vccd vccd wire1351/X sky130_fd_sc_hd__buf_6
Xwire2096 wire2096/A vssd vssd vccd vccd wire2096/X sky130_fd_sc_hd__buf_6
Xwire1362 wire1362/A vssd vssd vccd vccd _366_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1373 wire1374/X vssd vssd vccd vccd wire1373/X sky130_fd_sc_hd__buf_6
XFILLER_47_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1384 wire1384/A vssd vssd vccd vccd wire1384/X sky130_fd_sc_hd__buf_6
XFILLER_46_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1395 wire1396/X vssd vssd vccd vccd wire1395/X sky130_fd_sc_hd__buf_6
XFILLER_38_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2802 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_882 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1105_A _408_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_309_ _309_/A _309_/B vssd vssd vccd vccd _309_/X sky130_fd_sc_hd__and2_2
XFILLER_30_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[73\]_B _236_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output843_A _594_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__162__A _162_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1474_A wire1474/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] wire1324/X vssd vssd vccd vccd wire967/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_28_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1641_A wire1642/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1739_A wire1739/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1906_A wire1907/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__337__A _337_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_576 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__072__A _072_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput304 la_oenb_mprj[24] vssd vssd vccd vccd _521_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput315 la_oenb_mprj[34] vssd vssd vccd vccd _531_/A sky130_fd_sc_hd__buf_4
XFILLER_44_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput326 la_oenb_mprj[44] vssd vssd vccd vccd _541_/A sky130_fd_sc_hd__buf_6
Xinput337 la_oenb_mprj[54] vssd vssd vccd vccd _551_/A sky130_fd_sc_hd__buf_8
XFILLER_29_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput348 la_oenb_mprj[64] vssd vssd vccd vccd wire1553/A sky130_fd_sc_hd__buf_6
XFILLER_40_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput359 la_oenb_mprj[74] vssd vssd vccd vccd wire1543/A sky130_fd_sc_hd__buf_6
XFILLER_5_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_591_ _591_/A _591_/B vssd vssd vccd vccd _591_/X sky130_fd_sc_hd__and2_4
XFILLER_35_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2122_A wire2122/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input205_A la_iena_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__247__A _247_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_025_ _025_/A vssd vssd vccd vccd _025_/Y sky130_fd_sc_hd__inv_2
XANTENNA_8 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__413__C _413_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1170 wire1171/X vssd vssd vccd vccd wire1170/X sky130_fd_sc_hd__buf_8
XFILLER_19_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1181 _360_/X vssd vssd vccd vccd wire1181/X sky130_fd_sc_hd__buf_6
XFILLER_47_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1192 wire1193/X vssd vssd vccd vccd wire1192/X sky130_fd_sc_hd__buf_6
XFILLER_1_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__295__A_N _295_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1222_A _348_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output793_A _548_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1076 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1689_A wire1689/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__604__B _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1856_A wire1856/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__620__A _620_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__067__A _067_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[37\]_B _200_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[121\]_B _284_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__514__B _514_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__530__A _530_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input155_A la_iena_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput101 la_data_out_mprj[72] vssd vssd vccd vccd wire1632/A sky130_fd_sc_hd__buf_6
XFILLER_7_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput112 la_data_out_mprj[82] vssd vssd vccd vccd wire1622/A sky130_fd_sc_hd__buf_6
XFILLER_24_2845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput123 la_data_out_mprj[92] vssd vssd vccd vccd _461_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput134 la_iena_mprj[101] vssd vssd vccd vccd _264_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 la_iena_mprj[111] vssd vssd vccd vccd _274_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput156 la_iena_mprj[121] vssd vssd vccd vccd _284_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input322_A la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput167 la_iena_mprj[16] vssd vssd vccd vccd _179_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput178 la_iena_mprj[26] vssd vssd vccd vccd wire1612/A sky130_fd_sc_hd__buf_6
XTAP_4655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 la_iena_mprj[36] vssd vssd vccd vccd _199_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_574_ _574_/A _574_/B vssd vssd vccd vccd _574_/X sky130_fd_sc_hd__and2_4
XANTENNA_user_wb_dat_gates\[30\]_A mprj_dat_i_user[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3940 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__424__B _424_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[112\]_B _275_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput608 _098_/Y vssd vssd vccd vccd la_data_in_mprj[115] sky130_fd_sc_hd__buf_8
Xoutput619 _108_/Y vssd vssd vccd vccd la_data_in_mprj[125] sky130_fd_sc_hd__buf_8
X_008_ _008_/A vssd vssd vccd vccd _008_/Y sky130_fd_sc_hd__inv_4
XFILLER_29_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output541_A wire1087/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output639_A _011_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1172_A wire1173/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output806_A _560_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1437_A wire1438/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] _216_/X vssd vssd vccd vccd _036_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_48_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1604_A _472_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[21\]_A mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__615__A _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1973_A wire1974/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[19\]_B _182_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__334__B _334_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_B wire1316/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__350__A _350_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__460__A_N _588_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input8_A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1906 wire1907/X vssd vssd vccd vccd wire1906/X sky130_fd_sc_hd__buf_6
XTAP_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1917 wire1918/X vssd vssd vccd vccd wire1917/X sky130_fd_sc_hd__buf_6
XTAP_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1928 wire1929/X vssd vssd vccd vccd _607_/B sky130_fd_sc_hd__buf_6
XTAP_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1939 wire1940/X vssd vssd vccd vccd _603_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__509__B _509_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_228 _204_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_239 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[12\]_A mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_290_ _290_/A _290_/B vssd vssd vccd vccd _290_/X sky130_fd_sc_hd__and2_4
XFILLER_17_2682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__525__A _525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__244__B _244_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input272_A la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__260__A _260_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__419__B _419_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_557_ _557_/A _557_/B vssd vssd vccd vccd _557_/X sky130_fd_sc_hd__and2_2
XFILLER_31_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1018_A _538_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_488_ _616_/A _488_/B _488_/C vssd vssd vccd vccd _488_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output491_A _494_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output589_A wire1067/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output756_A wire1034/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1387_A wire1388/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__483__A_N _611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output923_A wire1194/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__170__A _170_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1721_A wire1722/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__329__B _329_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1856 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__345__A _345_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__080__A _080_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput950 wire1299/X vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__buf_8
XFILLER_25_4375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1703 wire1703/A vssd vssd vccd vccd wire1703/X sky130_fd_sc_hd__buf_6
XFILLER_43_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1714 wire1714/A vssd vssd vccd vccd _300_/A sky130_fd_sc_hd__buf_6
Xwire1725 wire1725/A vssd vssd vccd vccd wire1725/X sky130_fd_sc_hd__buf_6
XFILLER_4_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1736 wire1737/X vssd vssd vccd vccd wire1736/X sky130_fd_sc_hd__buf_6
XFILLER_41_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4102 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1747 wire1748/X vssd vssd vccd vccd wire1747/X sky130_fd_sc_hd__buf_6
XTAP_3003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1758 wire1758/A vssd vssd vccd vccd wire1758/X sky130_fd_sc_hd__buf_6
XFILLER_2_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1769 wire1770/X vssd vssd vccd vccd _274_/A sky130_fd_sc_hd__buf_6
XTAP_3014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__239__B _239_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2035_A wire2035/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_411_ _539_/A _411_/B _411_/C vssd vssd vccd vccd _411_/X sky130_fd_sc_hd__and3b_4
XFILLER_27_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_446 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_342_ _342_/A _342_/B vssd vssd vccd vccd _342_/X sky130_fd_sc_hd__and2_2
XTAP_1678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__255__A _255_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_273_ _273_/A _273_/B vssd vssd vccd vccd _273_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input83_A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__421__C _421_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output504_A wire1123/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1135_A _379_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_609_ _609_/A _609_/B vssd vssd vccd vccd _609_/X sky130_fd_sc_hd__and2_4
XFILLER_53_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1302_A _300_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output873_A _308_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__165__A _165_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] _179_/X vssd vssd vccd vccd _163_/A
+ sky130_fd_sc_hd__nand2_4
Xuser_wb_dat_gates\[29\] mprj_dat_i_user[29] max_length1310/X vssd vssd vccd vccd
+ _143_/A sky130_fd_sc_hd__nand2_8
XFILLER_31_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1671_A wire1671/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1769_A wire1770/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__612__B _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1936_A wire1936/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] _290_/X vssd vssd vccd vccd wire979/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__379__A_N _507_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__075__A _075_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_950 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__522__B _522_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput780 wire1050/X vssd vssd vccd vccd la_oenb_core[3] sky130_fd_sc_hd__buf_8
Xwire2201 wire2202/X vssd vssd vccd vccd _305_/A sky130_fd_sc_hd__buf_6
Xoutput791 wire1049/X vssd vssd vccd vccd la_oenb_core[4] sky130_fd_sc_hd__buf_8
XFILLER_40_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1500 wire1500/A vssd vssd vccd vccd wire1500/X sky130_fd_sc_hd__buf_6
XFILLER_8_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3346 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1511 wire1511/A vssd vssd vccd vccd wire1511/X sky130_fd_sc_hd__buf_6
XFILLER_48_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input235_A la_iena_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1522 wire1523/X vssd vssd vccd vccd _305_/B sky130_fd_sc_hd__buf_8
XFILLER_24_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2152_A wire2153/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1533 wire1533/A vssd vssd vccd vccd _581_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1544 wire1544/A vssd vssd vccd vccd _570_/A sky130_fd_sc_hd__buf_6
XFILLER_38_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1555 wire1555/A vssd vssd vccd vccd _559_/A sky130_fd_sc_hd__buf_6
Xwire1566 input32/X vssd vssd vccd vccd _494_/C sky130_fd_sc_hd__buf_6
Xwire1577 wire1578/X vssd vssd vccd vccd wire1577/X sky130_fd_sc_hd__buf_6
XFILLER_24_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1588 wire1588/A vssd vssd vccd vccd _615_/A sky130_fd_sc_hd__buf_6
XFILLER_41_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1599 _477_/A_N vssd vssd vccd vccd _605_/A sky130_fd_sc_hd__buf_4
XFILLER_41_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input402_A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ _325_/A _325_/B vssd vssd vccd vccd _325_/X sky130_fd_sc_hd__and2_4
XFILLER_30_736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__416__C _416_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_256_ _256_/A _256_/B vssd vssd vccd vccd _256_/X sky130_fd_sc_hd__and2_4
XFILLER_7_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_187_ _187_/A _187_/B vssd vssd vccd vccd _187_/X sky130_fd_sc_hd__and2_2
XFILLER_48_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__432__B _432_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1085_A wire1086/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output719_A wire1053/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1252_A _337_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1517_A wire1517/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__607__B _607_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1886_A wire1887/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__623__A _623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__342__B _342_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[4\]_A mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__517__B _517_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_110_ _110_/A vssd vssd vccd vccd _110_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_36_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__533__A _533_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_041_ _041_/A vssd vssd vccd vccd _041_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input185_A la_iena_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__252__B _252_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input352_A la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input46_A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2020 wire2020/A vssd vssd vccd vccd _561_/B sky130_fd_sc_hd__buf_6
XFILLER_1_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2031 wire2031/A vssd vssd vccd vccd _519_/B sky130_fd_sc_hd__buf_6
XFILLER_43_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2042 wire2043/X vssd vssd vccd vccd _510_/B sky130_fd_sc_hd__buf_6
Xwire2053 wire2054/X vssd vssd vccd vccd _503_/B sky130_fd_sc_hd__buf_6
XFILLER_1_3226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2064 wire2065/X vssd vssd vccd vccd _497_/B sky130_fd_sc_hd__buf_6
Xwire1330 _247_/X vssd vssd vccd vccd wire1330/X sky130_fd_sc_hd__buf_8
Xwire2075 wire2075/A vssd vssd vccd vccd wire2075/X sky130_fd_sc_hd__buf_6
Xwire1341 wire1341/A vssd vssd vccd vccd _300_/B sky130_fd_sc_hd__buf_6
Xwire2086 wire2087/X vssd vssd vccd vccd wire2086/X sky130_fd_sc_hd__buf_6
XFILLER_21_3187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1352 wire1353/X vssd vssd vccd vccd _342_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2097 wire2098/X vssd vssd vccd vccd _486_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1363 wire1363/A vssd vssd vccd vccd _365_/B sky130_fd_sc_hd__buf_6
Xwire1374 wire1374/A vssd vssd vccd vccd wire1374/X sky130_fd_sc_hd__buf_6
XFILLER_21_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1385 wire1386/X vssd vssd vccd vccd _349_/B sky130_fd_sc_hd__buf_6
Xwire1396 wire1397/X vssd vssd vccd vccd wire1396/X sky130_fd_sc_hd__buf_6
XFILLER_46_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__427__B _427_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2814 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_308_ _308_/A _308_/B vssd vssd vccd vccd _308_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1000_A wire1001/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output571_A _451_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_239_ _239_/A _239_/B vssd vssd vccd vccd _239_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output836_A wire994/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1467_A wire1468/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] wire1331/X vssd vssd vccd vccd wire974/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_3098 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1634_A wire1634/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__618__A _618_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__337__B _337_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__417__A_N _417_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__353__A _353_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput305 la_oenb_mprj[25] vssd vssd vccd vccd _522_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput316 la_oenb_mprj[35] vssd vssd vccd vccd wire1569/A sky130_fd_sc_hd__buf_6
XFILLER_2_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput327 la_oenb_mprj[45] vssd vssd vccd vccd _542_/A sky130_fd_sc_hd__buf_4
XFILLER_22_3452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput338 la_oenb_mprj[55] vssd vssd vccd vccd _552_/A sky130_fd_sc_hd__buf_4
XFILLER_5_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput349 la_oenb_mprj[65] vssd vssd vccd vccd wire1552/A sky130_fd_sc_hd__buf_6
XFILLER_2_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_590_ _590_/A _590_/B vssd vssd vccd vccd _590_/X sky130_fd_sc_hd__and2_4
XFILLER_2_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__528__A _528_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input100_A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2115_A wire2116/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__263__A _263_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_024_ _024_/A vssd vssd vccd vccd _024_/Y sky130_fd_sc_hd__inv_2
XANTENNA_9 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1160 wire1161/X vssd vssd vccd vccd wire1160/X sky130_fd_sc_hd__buf_6
Xwire1171 wire1172/X vssd vssd vccd vccd wire1171/X sky130_fd_sc_hd__buf_6
Xwire1182 wire1183/X vssd vssd vccd vccd wire1182/X sky130_fd_sc_hd__buf_8
XFILLER_1_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1193 _357_/X vssd vssd vccd vccd wire1193/X sky130_fd_sc_hd__buf_6
XFILLER_47_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1048_A _502_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1215_A wire1216/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output786_A wire1013/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output953_A wire2205/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__173__A _173_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[11\] mprj_dat_i_user[11] _294_/X vssd vssd vccd vccd _125_/A sky130_fd_sc_hd__nand2_2
XFILLER_51_2991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1751_A wire1752/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1849_A wire1849/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__620__B _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__348__A _348_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__083__A _083_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__530__B _530_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput102 la_data_out_mprj[73] vssd vssd vccd vccd wire1631/A sky130_fd_sc_hd__buf_6
Xinput113 la_data_out_mprj[83] vssd vssd vccd vccd wire1621/A sky130_fd_sc_hd__buf_6
XFILLER_7_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput124 la_data_out_mprj[93] vssd vssd vccd vccd _462_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2065_A wire2065/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input148_A la_iena_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput135 la_iena_mprj[102] vssd vssd vccd vccd _265_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput146 la_iena_mprj[112] vssd vssd vccd vccd _275_/B sky130_fd_sc_hd__buf_4
XFILLER_22_3271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput157 la_iena_mprj[122] vssd vssd vccd vccd _285_/B sky130_fd_sc_hd__buf_4
XTAP_4634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 la_iena_mprj[17] vssd vssd vccd vccd _180_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 la_iena_mprj[27] vssd vssd vccd vccd _190_/B sky130_fd_sc_hd__buf_4
XFILLER_29_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input315_A la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__258__A _258_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_573_ _573_/A _573_/B vssd vssd vccd vccd _573_/X sky130_fd_sc_hd__and2_4
XTAP_3988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[30\]_B max_length1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3952 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__424__C _424_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput609 _099_/Y vssd vssd vccd vccd la_data_in_mprj[116] sky130_fd_sc_hd__buf_8
XFILLER_29_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_007_ _007_/A vssd vssd vccd vccd _007_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_46_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__440__B _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output534_A wire1095/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1165_A _364_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1332_A _243_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__168__A _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] _209_/X vssd vssd vccd vccd _029_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_B max_length1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__615__B _615_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] _171_/X vssd vssd vccd vccd _155_/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA__350__B _350_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1907 wire1907/A vssd vssd vccd vccd wire1907/X sky130_fd_sc_hd__buf_6
XFILLER_41_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1918 wire1918/A vssd vssd vccd vccd wire1918/X sky130_fd_sc_hd__buf_6
Xwire1929 wire1930/X vssd vssd vccd vccd wire1929/X sky130_fd_sc_hd__buf_6
XTAP_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__078__A _078_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_207 _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_218 _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 _204_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_978 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[12\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__525__B _525_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__541__A _541_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2182_A wire2183/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input265_A la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__260__B _260_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input432_A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_625_ _625_/A _625_/B vssd vssd vccd vccd _625_/X sky130_fd_sc_hd__and2_1
XTAP_3763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__419__C _419_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_556_ _556_/A _556_/B vssd vssd vccd vccd _556_/X sky130_fd_sc_hd__and2_2
XFILLER_50_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_487_ _615_/A _487_/B _487_/C vssd vssd vccd vccd _487_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__435__B _435_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output484_A _488_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output651_A _022_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output749_A _624_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1282_A wire1283/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output916_A wire1217/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3742 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3786 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1714_A wire1714/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4258 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__345__B _345_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__361__A _361_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput940 wire1238/X vssd vssd vccd vccd mprj_dat_o_user[5] sky130_fd_sc_hd__buf_8
XFILLER_5_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput951 wire1723/X vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_47_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1704 wire1705/X vssd vssd vccd vccd _362_/A sky130_fd_sc_hd__buf_6
XFILLER_28_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1715 wire1715/A vssd vssd vccd vccd _354_/A sky130_fd_sc_hd__buf_6
XFILLER_25_2985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1726 wire1727/X vssd vssd vccd vccd _293_/A sky130_fd_sc_hd__buf_6
XTAP_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1737 wire1737/A vssd vssd vccd vccd wire1737/X sky130_fd_sc_hd__buf_6
Xwire1748 wire1748/A vssd vssd vccd vccd wire1748/X sky130_fd_sc_hd__buf_6
XTAP_3004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1759 wire1760/X vssd vssd vccd vccd _279_/A sky130_fd_sc_hd__buf_6
XFILLER_19_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ _538_/A _410_/B _410_/C vssd vssd vccd vccd _410_/X sky130_fd_sc_hd__and3b_4
XTAP_2347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_341_ _341_/A _341_/B vssd vssd vccd vccd _341_/X sky130_fd_sc_hd__and2_2
XFILLER_36_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__255__B _255_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_272_ _272_/A _272_/B vssd vssd vccd vccd _272_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input382_A la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input76_A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__271__A _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_608_ _608_/A _608_/B vssd vssd vccd vccd _608_/X sky130_fd_sc_hd__and2_4
XTAP_3593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1030_A _519_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1128_A _385_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_539_ _539_/A _539_/B vssd vssd vccd vccd _539_/X sky130_fd_sc_hd__and2_2
XFILLER_32_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__450__A_N _578_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output866_A _331_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1497_A wire1497/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__181__A _181_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1664_A wire1665/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1831_A wire1832/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1929_A wire1930/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__356__A _356_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__091__A _091_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4026 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput770 _527_/X vssd vssd vccd vccd la_oenb_core[30] sky130_fd_sc_hd__buf_8
Xoutput781 _537_/X vssd vssd vccd vccd la_oenb_core[40] sky130_fd_sc_hd__buf_8
XFILLER_47_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2202 wire2202/A vssd vssd vccd vccd wire2202/X sky130_fd_sc_hd__buf_6
Xoutput792 wire1009/X vssd vssd vccd vccd la_oenb_core[50] sky130_fd_sc_hd__buf_8
XFILLER_43_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1501 wire1502/X vssd vssd vccd vccd _321_/B sky130_fd_sc_hd__buf_6
Xwire1512 wire1513/X vssd vssd vccd vccd _318_/B sky130_fd_sc_hd__buf_6
XFILLER_38_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1523 wire1524/X vssd vssd vccd vccd wire1523/X sky130_fd_sc_hd__buf_6
XFILLER_21_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1534 wire1534/A vssd vssd vccd vccd _580_/A sky130_fd_sc_hd__buf_6
Xwire1545 wire1545/A vssd vssd vccd vccd _569_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input130_A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1556 wire1556/A vssd vssd vccd vccd _555_/A sky130_fd_sc_hd__buf_6
XFILLER_38_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2145_A wire2145/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1567 _406_/A_N vssd vssd vccd vccd _534_/A sky130_fd_sc_hd__buf_6
XFILLER_21_2668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1578 input3/X vssd vssd vccd vccd wire1578/X sky130_fd_sc_hd__buf_6
XANTENNA_input228_A la_iena_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1589 wire1589/A vssd vssd vccd vccd _614_/A sky130_fd_sc_hd__buf_6
XTAP_2100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__473__A_N _601_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__266__A _266_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_324_ _324_/A _324_/B vssd vssd vccd vccd _324_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_255_ _255_/A _255_/B vssd vssd vccd vccd _255_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_186_ _186_/A _186_/B vssd vssd vccd vccd _186_/X sky130_fd_sc_hd__and2_2
XFILLER_7_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__432__C _432_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3076 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1245_A _340_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1412_A wire1413/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__176__A _176_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1781_A wire1781/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1879_A wire1880/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__623__B _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[4\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__496__A_N _624_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1162 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__086__A _086_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_040_ _040_/A vssd vssd vccd vccd _040_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2095_A wire2096/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input178_A la_iena_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input345_A la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2010 wire2011/X vssd vssd vccd vccd _569_/B sky130_fd_sc_hd__buf_6
Xwire2021 wire2021/A vssd vssd vccd vccd _560_/B sky130_fd_sc_hd__buf_6
Xwire2032 wire2032/A vssd vssd vccd vccd _518_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input39_A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2043 wire2043/A vssd vssd vccd vccd wire2043/X sky130_fd_sc_hd__buf_6
Xwire2054 wire2054/A vssd vssd vccd vccd wire2054/X sky130_fd_sc_hd__buf_6
XFILLER_43_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1320 _257_/X vssd vssd vccd vccd wire1320/X sky130_fd_sc_hd__buf_6
Xwire2065 wire2065/A vssd vssd vccd vccd wire2065/X sky130_fd_sc_hd__buf_6
Xwire2076 wire2077/X vssd vssd vccd vccd _493_/B sky130_fd_sc_hd__buf_6
Xwire1331 _246_/X vssd vssd vccd vccd wire1331/X sky130_fd_sc_hd__buf_6
XFILLER_1_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1342 wire1343/X vssd vssd vccd vccd _299_/B sky130_fd_sc_hd__buf_6
Xwire2087 wire2087/A vssd vssd vccd vccd wire2087/X sky130_fd_sc_hd__buf_6
XFILLER_1_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1353 wire1353/A vssd vssd vccd vccd wire1353/X sky130_fd_sc_hd__buf_6
Xwire2098 wire2098/A vssd vssd vccd vccd wire2098/X sky130_fd_sc_hd__buf_6
XFILLER_5_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1364 wire1364/A vssd vssd vccd vccd _364_/B sky130_fd_sc_hd__buf_6
XFILLER_46_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1375 wire1375/A vssd vssd vccd vccd _356_/B sky130_fd_sc_hd__buf_6
Xwire1386 wire1386/A vssd vssd vccd vccd wire1386/X sky130_fd_sc_hd__buf_6
Xwire1397 wire1397/A vssd vssd vccd vccd wire1397/X sky130_fd_sc_hd__buf_6
XFILLER_1_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__427__C _427_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_307_ _307_/A _307_/B vssd vssd vccd vccd _307_/X sky130_fd_sc_hd__and2_2
XFILLER_50_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_238_ _238_/A _238_/B vssd vssd vccd vccd _238_/X sky130_fd_sc_hd__and2_4
XANTENNA__443__B _443_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output564_A _445_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__369__A_N _497_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_169_ _169_/A _169_/B vssd vssd vccd vccd _169_/X sky130_fd_sc_hd__and2_2
XFILLER_7_796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1195_A wire1196/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output731_A _607_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output829_A _581_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] _239_/X vssd vssd vccd vccd _059_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_23_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1627_A wire1627/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__618__B _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1996_A wire1997/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__353__B _353_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput306 la_oenb_mprj[26] vssd vssd vccd vccd _523_/A sky130_fd_sc_hd__buf_4
Xinput317 la_oenb_mprj[36] vssd vssd vccd vccd _405_/A_N sky130_fd_sc_hd__buf_6
Xinput328 la_oenb_mprj[46] vssd vssd vccd vccd _415_/A_N sky130_fd_sc_hd__buf_6
Xinput339 la_oenb_mprj[56] vssd vssd vccd vccd _553_/A sky130_fd_sc_hd__buf_4
XFILLER_22_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1382 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3475 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__528__B _528_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2010_A wire2011/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2108_A wire2109/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__544__A _544_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input295_A la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__263__B _263_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_023_ _023_/A vssd vssd vccd vccd _023_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input462_A user_irq_ena[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1150 wire1151/X vssd vssd vccd vccd wire1150/X sky130_fd_sc_hd__buf_8
XFILLER_48_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1161 _365_/X vssd vssd vccd vccd wire1161/X sky130_fd_sc_hd__buf_6
XFILLER_40_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1172 wire1173/X vssd vssd vccd vccd wire1172/X sky130_fd_sc_hd__buf_6
XFILLER_1_2334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1183 wire1184/X vssd vssd vccd vccd wire1183/X sky130_fd_sc_hd__buf_6
Xwire1194 wire1195/X vssd vssd vccd vccd wire1194/X sky130_fd_sc_hd__buf_8
XFILLER_34_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__438__B _438_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1110_A _403_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1208_A wire1209/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output779_A wire1019/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_34_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output946_A wire1289/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1577_A wire1578/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1744_A wire1745/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1911_A wire1912/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] _265_/X vssd vssd vccd vccd _085_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA__348__B _348_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__364__A _364_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput103 la_data_out_mprj[74] vssd vssd vccd vccd wire1630/A sky130_fd_sc_hd__buf_6
Xinput114 la_data_out_mprj[84] vssd vssd vccd vccd wire1620/A sky130_fd_sc_hd__buf_6
XFILLER_49_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput125 la_data_out_mprj[94] vssd vssd vccd vccd _463_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput136 la_iena_mprj[103] vssd vssd vccd vccd _266_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput147 la_iena_mprj[113] vssd vssd vccd vccd _276_/B sky130_fd_sc_hd__buf_4
XTAP_4624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput158 la_iena_mprj[123] vssd vssd vccd vccd _286_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput169 la_iena_mprj[18] vssd vssd vccd vccd _181_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire2058_A wire2059/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__539__A _539_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input210_A la_iena_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_572_ _572_/A _572_/B vssd vssd vccd vccd _572_/X sky130_fd_sc_hd__and2_4
XFILLER_29_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input308_A la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__274__A _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_006_ _006_/A vssd vssd vccd vccd _006_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_29_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__440__C _440_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__407__A_N _535_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output527_A wire1102/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1060_A _475_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1158_A wire1159/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1325_A _252_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output896_A _137_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] _202_/X vssd vssd vccd vccd _022_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_23_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__184__A _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1694_A wire1695/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1861_A wire1861/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1959_A wire1960/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1908 wire1909/X vssd vssd vccd vccd _613_/B sky130_fd_sc_hd__buf_6
XTAP_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1919 wire1920/X vssd vssd vccd vccd _610_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__359__A _359_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__094__A _094_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input160_A la_iena_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input258_A la_iena_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2175_A wire2176/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input425_A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input21_A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__269__A _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_624_ _624_/A _624_/B vssd vssd vccd vccd _624_/X sky130_fd_sc_hd__and2_4
XTAP_4498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_555_ _555_/A _555_/B vssd vssd vccd vccd _555_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_486_ _614_/A _486_/B _486_/C vssd vssd vccd vccd _486_/X sky130_fd_sc_hd__and3b_4
XFILLER_18_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__435__C _435_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output477_A wire1054/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__451__B _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output644_A _015_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1275_A _314_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output811_A _565_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1442_A wire1443/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__179__A _179_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_702 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__361__B _361_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput930 wire1170/X vssd vssd vccd vccd mprj_dat_o_user[25] sky130_fd_sc_hd__buf_8
Xoutput941 wire1235/X vssd vssd vccd vccd mprj_dat_o_user[6] sky130_fd_sc_hd__buf_8
Xoutput952 output952/A vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_5_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1705 wire1705/A vssd vssd vccd vccd wire1705/X sky130_fd_sc_hd__buf_6
Xwire1716 wire1716/A vssd vssd vccd vccd _353_/A sky130_fd_sc_hd__buf_6
XFILLER_28_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1727 wire1728/X vssd vssd vccd vccd wire1727/X sky130_fd_sc_hd__buf_6
XTAP_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__089__A _089_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1738 wire1739/X vssd vssd vccd vccd _289_/A sky130_fd_sc_hd__buf_6
Xwire1749 wire1750/X vssd vssd vccd vccd _284_/A sky130_fd_sc_hd__buf_6
XTAP_3005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ _340_/A _340_/B vssd vssd vccd vccd _340_/X sky130_fd_sc_hd__and2_4
XFILLER_41_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__536__B _536_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_271_ _271_/A _271_/B vssd vssd vccd vccd _271_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__552__A _552_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input375_A la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__271__B _271_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input69_A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_607_ _607_/A _607_/B vssd vssd vccd vccd _607_/X sky130_fd_sc_hd__and2_4
XFILLER_45_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__446__B _446_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_538_ _538_/A _538_/B vssd vssd vccd vccd _538_/X sky130_fd_sc_hd__and2_4
XTAP_2893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output594_A _085_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_469_ _597_/A _469_/B _469_/C vssd vssd vccd vccd _469_/X sky130_fd_sc_hd__and3b_2
XFILLER_32_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output761_A wire1030/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output859_A _306_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1392_A wire1393/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__181__B _181_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1657_A wire1658/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__356__B _356_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_B wire1320/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3738 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1298 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput760 wire1031/X vssd vssd vccd vccd la_oenb_core[21] sky130_fd_sc_hd__buf_8
XFILLER_5_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput771 _528_/X vssd vssd vccd vccd la_oenb_core[31] sky130_fd_sc_hd__buf_8
XFILLER_40_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput782 wire1018/X vssd vssd vccd vccd la_oenb_core[41] sky130_fd_sc_hd__buf_8
XFILLER_8_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2203 wire2204/X vssd vssd vccd vccd _295_/B sky130_fd_sc_hd__buf_6
Xoutput793 _548_/X vssd vssd vccd vccd la_oenb_core[51] sky130_fd_sc_hd__buf_8
XFILLER_47_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1502 wire1503/X vssd vssd vccd vccd wire1502/X sky130_fd_sc_hd__buf_6
XFILLER_24_1014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1513 wire1514/X vssd vssd vccd vccd wire1513/X sky130_fd_sc_hd__buf_6
XFILLER_24_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1524 wire1525/X vssd vssd vccd vccd wire1524/X sky130_fd_sc_hd__buf_6
Xwire1535 wire1535/A vssd vssd vccd vccd _579_/A sky130_fd_sc_hd__buf_6
Xwire1546 wire1546/A vssd vssd vccd vccd _568_/A sky130_fd_sc_hd__buf_6
XFILLER_41_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1557 input34/X vssd vssd vccd vccd _496_/C sky130_fd_sc_hd__buf_4
Xwire1568 _405_/A_N vssd vssd vccd vccd _533_/A sky130_fd_sc_hd__buf_6
XFILLER_38_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1579 wire1579/A vssd vssd vccd vccd _624_/A sky130_fd_sc_hd__buf_6
XANTENNA_input123_A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2040_A wire2041/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2138_A wire2138/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__547__A _547_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__266__B _266_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_323_ _323_/A _323_/B vssd vssd vccd vccd _323_/X sky130_fd_sc_hd__and2_4
XFILLER_42_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[85\]_B wire1329/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_254_ _254_/A _254_/B vssd vssd vccd vccd _254_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__282__A _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_185_ _185_/A _185_/B vssd vssd vccd vccd _185_/X sky130_fd_sc_hd__and2_4
XFILLER_45_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[4\] mprj_dat_i_user[4] max_length1311/X vssd vssd vccd vccd _118_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_6_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1140_A _374_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1238_A wire1239/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1405_A wire1406/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] _184_/X vssd vssd vccd vccd _004_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_50_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_B _239_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__192__A _192_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1774_A wire1774/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1941_A wire1942/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__367__A _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2088_A wire2089/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2000 wire2000/A vssd vssd vccd vccd wire2000/X sky130_fd_sc_hd__buf_6
Xoutput590 wire1136/X vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__buf_8
XFILLER_44_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2011 wire2011/A vssd vssd vccd vccd wire2011/X sky130_fd_sc_hd__buf_6
XFILLER_21_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2022 wire2022/A vssd vssd vccd vccd _559_/B sky130_fd_sc_hd__buf_6
XANTENNA_input240_A la_iena_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2033 wire2033/A vssd vssd vccd vccd _517_/B sky130_fd_sc_hd__buf_6
XANTENNA_input338_A la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2044 wire2044/A vssd vssd vccd vccd _509_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2055 wire2056/X vssd vssd vccd vccd _502_/B sky130_fd_sc_hd__buf_6
XFILLER_40_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__440__A_N _568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1321 _256_/X vssd vssd vccd vccd wire1321/X sky130_fd_sc_hd__buf_6
Xwire2066 wire2067/X vssd vssd vccd vccd _496_/B sky130_fd_sc_hd__buf_6
Xwire2077 wire2078/X vssd vssd vccd vccd wire2077/X sky130_fd_sc_hd__buf_6
XFILLER_8_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1332 _243_/X vssd vssd vccd vccd wire1332/X sky130_fd_sc_hd__buf_6
XFILLER_38_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1343 wire1343/A vssd vssd vccd vccd wire1343/X sky130_fd_sc_hd__buf_6
Xwire2088 wire2089/X vssd vssd vccd vccd _489_/B sky130_fd_sc_hd__buf_6
Xwire2099 wire2100/X vssd vssd vccd vccd _485_/B sky130_fd_sc_hd__buf_6
Xwire1354 wire1355/X vssd vssd vccd vccd _341_/B sky130_fd_sc_hd__buf_6
Xwire1365 wire1365/A vssd vssd vccd vccd _363_/B sky130_fd_sc_hd__buf_6
XFILLER_19_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1376 wire1376/A vssd vssd vccd vccd _355_/B sky130_fd_sc_hd__buf_6
XFILLER_38_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1387 wire1388/X vssd vssd vccd vccd _348_/B sky130_fd_sc_hd__buf_6
Xwire1398 wire1399/X vssd vssd vccd vccd _314_/B sky130_fd_sc_hd__buf_6
XANTENNA__277__A _277_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_370 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_306_ _306_/A _306_/B vssd vssd vccd vccd _306_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_237_ _237_/A _237_/B vssd vssd vccd vccd _237_/X sky130_fd_sc_hd__and2_4
XANTENNA__443__C _443_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_742 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_168_ _168_/A _168_/B vssd vssd vccd vccd _168_/X sky130_fd_sc_hd__and2_2
XFILLER_13_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output557_A wire1139/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_099_ _099_/A vssd vssd vccd vccd _099_/Y sky130_fd_sc_hd__inv_2
XANTENNA_wire1090_A _422_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1188_A wire1189/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output724_A _601_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1355_A wire1355/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] _232_/X vssd vssd vccd vccd _052_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1522_A wire1523/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__187__A _187_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1891_A wire1891/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1989_A wire1989/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__463__A_N _591_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput307 la_oenb_mprj[27] vssd vssd vccd vccd wire1575/A sky130_fd_sc_hd__buf_6
Xinput318 la_oenb_mprj[37] vssd vssd vccd vccd _406_/A_N sky130_fd_sc_hd__buf_6
Xinput329 la_oenb_mprj[47] vssd vssd vccd vccd _416_/A_N sky130_fd_sc_hd__buf_6
XFILLER_6_3695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__097__A _097_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[124\]_B wire1312/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__544__B _544_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2003_A wire2004/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input190_A la_iena_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input288_A la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_022_ _022_/A vssd vssd vccd vccd _022_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__560__A _560_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input455_A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input51_A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1140 _374_/X vssd vssd vccd vccd wire1140/X sky130_fd_sc_hd__buf_6
XFILLER_1_3058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1151 wire1152/X vssd vssd vccd vccd wire1151/X sky130_fd_sc_hd__buf_6
Xwire1162 wire1163/X vssd vssd vccd vccd wire1162/X sky130_fd_sc_hd__buf_8
XFILLER_48_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1173 _362_/X vssd vssd vccd vccd wire1173/X sky130_fd_sc_hd__buf_6
Xwire1184 wire1185/X vssd vssd vccd vccd wire1184/X sky130_fd_sc_hd__buf_6
XFILLER_38_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1195 wire1196/X vssd vssd vccd vccd wire1195/X sky130_fd_sc_hd__buf_6
XANTENNA__438__C _438_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__454__B _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_B _278_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1103_A _410_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__486__A_N _614_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output841_A _592_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output939_A wire1241/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1472_A wire1473/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1904_A wire1904/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[24\]_A mprj_dat_i_user[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[106\]_B _269_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__364__B _364_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput104 la_data_out_mprj[75] vssd vssd vccd vccd wire1629/A sky130_fd_sc_hd__buf_6
XFILLER_40_2105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput115 la_data_out_mprj[85] vssd vssd vccd vccd wire1619/A sky130_fd_sc_hd__buf_6
Xinput126 la_data_out_mprj[95] vssd vssd vccd vccd _464_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput137 la_iena_mprj[104] vssd vssd vccd vccd _267_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput148 la_iena_mprj[114] vssd vssd vccd vccd _277_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput159 la_iena_mprj[124] vssd vssd vccd vccd _287_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__539__B _539_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[15\]_A mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_571_ _571_/A _571_/B vssd vssd vccd vccd _571_/X sky130_fd_sc_hd__and2_4
XTAP_3968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2120_A wire2120/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input203_A la_iena_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__555__A _555_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3932 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__274__B _274_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input99_A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__290__A _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_005_ _005_/A vssd vssd vccd vccd _005_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_4_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__449__B _449_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1053_A _497_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_958 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1220_A wire1221/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output791_A wire1049/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1318_A _259_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1687_A wire1687/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1854_A wire1855/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1909 wire1910/X vssd vssd vccd vccd wire1909/X sky130_fd_sc_hd__buf_6
XTAP_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__359__B _359_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2964 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_209 _232_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2070_A wire2071/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input153_A la_iena_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2168_A wire2168/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__269__B _269_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input320_A la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input418_A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_623_ _623_/A _623_/B vssd vssd vccd vccd _623_/X sky130_fd_sc_hd__and2_4
XFILLER_22_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_554_ _554_/A _554_/B vssd vssd vccd vccd _554_/X sky130_fd_sc_hd__and2_4
XTAP_3798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__285__A _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_485_ _613_/A _485_/B _485_/C vssd vssd vccd vccd _485_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2086 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__451__C _451_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output637_A _009_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1170_A wire1171/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1268_A wire1269/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output804_A wire996/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1435_A wire1436/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] _214_/X vssd vssd vccd vccd _034_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_40_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_714 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__195__A _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1214 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1971_A wire1971/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput920 wire1205/X vssd vssd vccd vccd mprj_dat_o_user[16] sky130_fd_sc_hd__buf_8
XFILLER_2_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput931 wire1166/X vssd vssd vccd vccd mprj_dat_o_user[26] sky130_fd_sc_hd__buf_8
Xoutput942 wire1232/X vssd vssd vccd vccd mprj_dat_o_user[7] sky130_fd_sc_hd__buf_8
XFILLER_8_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput953 wire2205/X vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_9_3885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input6_A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1706 wire1707/X vssd vssd vccd vccd _361_/A sky130_fd_sc_hd__buf_6
XTAP_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1717 wire1717/A vssd vssd vccd vccd _352_/A sky130_fd_sc_hd__buf_6
XTAP_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1728 wire1728/A vssd vssd vccd vccd wire1728/X sky130_fd_sc_hd__buf_6
XFILLER_3_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1739 wire1739/A vssd vssd vccd vccd wire1739/X sky130_fd_sc_hd__buf_6
XFILLER_25_2998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_270_ _270_/A _270_/B vssd vssd vccd vccd _270_/X sky130_fd_sc_hd__and2_1
XFILLER_41_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3902 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__552__B _552_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input270_A la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input368_A la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4052 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_606_ _606_/A _606_/B vssd vssd vccd vccd _606_/X sky130_fd_sc_hd__and2_4
XTAP_3573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_91 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_537_ _537_/A _537_/B vssd vssd vccd vccd _537_/X sky130_fd_sc_hd__and2_4
XTAP_2872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__446__C _446_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_468_ _596_/A _468_/B _468_/C vssd vssd vccd vccd _468_/X sky130_fd_sc_hd__and3b_4
XANTENNA_wire1016_A wire1017/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output587_A wire1069/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_399_ _527_/A _399_/B _399_/C vssd vssd vccd vccd _399_/X sky130_fd_sc_hd__and3b_2
XFILLER_31_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__462__B _462_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output754_A wire1036/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1385_A wire1386/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output921_A wire1202/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] wire1317/X vssd vssd vccd vccd wire961/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_29_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1817_A wire1817/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__372__B _372_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2980 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[7\]_A mprj_dat_i_user[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput750 wire1040/X vssd vssd vccd vccd la_oenb_core[12] sky130_fd_sc_hd__buf_8
Xoutput761 wire1030/X vssd vssd vccd vccd la_oenb_core[22] sky130_fd_sc_hd__buf_8
Xoutput772 _529_/X vssd vssd vccd vccd la_oenb_core[32] sky130_fd_sc_hd__buf_8
XFILLER_5_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput783 wire1016/X vssd vssd vccd vccd la_oenb_core[42] sky130_fd_sc_hd__buf_8
XFILLER_40_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2204 wire2204/A vssd vssd vccd vccd wire2204/X sky130_fd_sc_hd__buf_6
Xoutput794 wire1007/X vssd vssd vccd vccd la_oenb_core[52] sky130_fd_sc_hd__buf_8
XFILLER_5_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2030 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1503 wire1504/X vssd vssd vccd vccd wire1503/X sky130_fd_sc_hd__buf_6
Xwire1514 wire1514/A vssd vssd vccd vccd wire1514/X sky130_fd_sc_hd__buf_6
XFILLER_43_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1525 wire1526/X vssd vssd vccd vccd wire1525/X sky130_fd_sc_hd__buf_6
XFILLER_24_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1536 wire1536/A vssd vssd vccd vccd _578_/A sky130_fd_sc_hd__buf_6
XFILLER_1_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1547 wire1547/A vssd vssd vccd vccd _567_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1558 _420_/A_N vssd vssd vccd vccd _548_/A sky130_fd_sc_hd__buf_6
Xwire1569 wire1569/A vssd vssd vccd vccd _532_/A sky130_fd_sc_hd__buf_6
XFILLER_38_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__547__B _547_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input116_A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2033_A wire2033/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ _322_/A _322_/B vssd vssd vccd vccd _322_/X sky130_fd_sc_hd__and2_4
XTAP_1467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2200_A wire2200/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__563__A _563_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_253_ _253_/A _253_/B vssd vssd vccd vccd _253_/X sky130_fd_sc_hd__and2_4
XFILLER_14_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input81_A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_184_ _184_/A _184_/B vssd vssd vccd vccd _184_/X sky130_fd_sc_hd__and2_1
XFILLER_52_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3238 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output502_A wire1144/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__457__B _457_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1133_A wire1134/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1300_A wire1301/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output871_A _335_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] _177_/X vssd vssd vccd vccd _161_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_31_2210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[27\] mprj_dat_i_user[27] _294_/X vssd vssd vccd vccd _141_/A sky130_fd_sc_hd__nand2_2
XFILLER_33_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__192__B _192_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1767_A wire1768/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4440 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1934_A wire1935/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] _288_/X vssd vssd vccd vccd _108_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_9_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__367__B _367_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__392__A_N _520_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput580 wire1076/X vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__buf_8
XFILLER_40_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2001 wire2002/X vssd vssd vccd vccd _574_/B sky130_fd_sc_hd__buf_6
XFILLER_25_3271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput591 _147_/Y vssd vssd vccd vccd la_data_in_mprj[0] sky130_fd_sc_hd__buf_8
Xwire2012 wire2013/X vssd vssd vccd vccd _568_/B sky130_fd_sc_hd__buf_6
XFILLER_27_2879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2023 wire2023/A vssd vssd vccd vccd _546_/B sky130_fd_sc_hd__buf_4
XFILLER_8_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2034 wire2034/A vssd vssd vccd vccd _516_/B sky130_fd_sc_hd__buf_6
Xwire1300 wire1301/X vssd vssd vccd vccd wire1300/X sky130_fd_sc_hd__buf_6
Xwire2045 wire2046/X vssd vssd vccd vccd _508_/B sky130_fd_sc_hd__buf_6
Xwire2056 wire2056/A vssd vssd vccd vccd wire2056/X sky130_fd_sc_hd__buf_6
XFILLER_21_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1322 _255_/X vssd vssd vccd vccd wire1322/X sky130_fd_sc_hd__buf_6
XFILLER_5_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2067 wire2068/X vssd vssd vccd vccd wire2067/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2150_A wire2151/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input233_A la_iena_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2078 wire2078/A vssd vssd vccd vccd wire2078/X sky130_fd_sc_hd__buf_6
Xwire1333 _242_/X vssd vssd vccd vccd wire1333/X sky130_fd_sc_hd__buf_6
XFILLER_5_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1344 wire1345/X vssd vssd vccd vccd _346_/B sky130_fd_sc_hd__buf_6
Xwire2089 wire2090/X vssd vssd vccd vccd wire2089/X sky130_fd_sc_hd__buf_6
XFILLER_38_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__558__A _558_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1355 wire1355/A vssd vssd vccd vccd wire1355/X sky130_fd_sc_hd__buf_6
Xwire1366 wire1366/A vssd vssd vccd vccd _362_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1377 wire1377/A vssd vssd vccd vccd _354_/B sky130_fd_sc_hd__buf_6
XFILLER_35_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1388 wire1388/A vssd vssd vccd vccd wire1388/X sky130_fd_sc_hd__buf_6
XFILLER_38_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1399 wire1400/X vssd vssd vccd vccd wire1399/X sky130_fd_sc_hd__buf_6
XANTENNA_input400_A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__277__B _277_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__293__A _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_305_ _305_/A _305_/B vssd vssd vccd vccd _305_/X sky130_fd_sc_hd__and2_2
XFILLER_15_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_236_ _236_/A _236_/B vssd vssd vccd vccd _236_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_167_ _167_/A _167_/B vssd vssd vccd vccd _167_/X sky130_fd_sc_hd__and2_1
XFILLER_6_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_098_ _098_/A vssd vssd vccd vccd _098_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_3024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1083_A _427_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output717_A _082_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1250_A _338_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1348_A wire1349/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__187__B _187_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1515_A wire1516/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1884_A wire1885/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire968_A wire968/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput308 la_oenb_mprj[28] vssd vssd vccd vccd _525_/A sky130_fd_sc_hd__buf_4
XFILLER_9_2074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput319 la_oenb_mprj[38] vssd vssd vccd vccd _535_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2859 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_021_ _021_/A vssd vssd vccd vccd _021_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input183_A la_iena_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__560__B _560_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input350_A la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input448_A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input44_A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1130 _383_/X vssd vssd vccd vccd wire1130/X sky130_fd_sc_hd__buf_6
XFILLER_40_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__288__A _288_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1141 _373_/X vssd vssd vccd vccd wire1141/X sky130_fd_sc_hd__buf_6
XFILLER_43_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1152 wire1153/X vssd vssd vccd vccd wire1152/X sky130_fd_sc_hd__buf_6
Xwire1163 wire1164/X vssd vssd vccd vccd wire1163/X sky130_fd_sc_hd__buf_6
XFILLER_38_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1174 wire1175/X vssd vssd vccd vccd wire1174/X sky130_fd_sc_hd__buf_8
Xwire1185 _359_/X vssd vssd vccd vccd wire1185/X sky130_fd_sc_hd__buf_6
XFILLER_34_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1196 wire1197/X vssd vssd vccd vccd wire1196/X sky130_fd_sc_hd__buf_6
XFILLER_35_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_628 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__454__C _454_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_219_ _219_/A _219_/B vssd vssd vccd vccd _219_/X sky130_fd_sc_hd__and2_2
XFILLER_32_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1298_A _301_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__470__B _470_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output834_A wire995/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1465_A wire1466/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] _244_/X vssd vssd vccd vccd wire975/A
+ sky130_fd_sc_hd__nand2_1
XTAP_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__198__A _198_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_606 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[24\]_B _294_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_672 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2747 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__430__A_N _558_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__380__B _380_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput105 la_data_out_mprj[76] vssd vssd vccd vccd wire1628/A sky130_fd_sc_hd__buf_6
Xinput116 la_data_out_mprj[86] vssd vssd vccd vccd wire1618/A sky130_fd_sc_hd__buf_6
XFILLER_24_2849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput127 la_data_out_mprj[96] vssd vssd vccd vccd _465_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput138 la_iena_mprj[105] vssd vssd vccd vccd _268_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput149 la_iena_mprj[115] vssd vssd vccd vccd _278_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_6_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[15\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_570_ _570_/A _570_/B vssd vssd vccd vccd _570_/X sky130_fd_sc_hd__and2_4
XTAP_3958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__555__B _555_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2113_A wire2114/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input398_A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__571__A _571_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_004_ _004_/A vssd vssd vccd vccd _004_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__290__B _290_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1800 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__449__C _449_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_A user_irq_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1046_A _504_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__465__B _465_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1213_A _351_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__453__A_N _581_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output784_A _540_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output951_A wire1723/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1847_A wire1848/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__375__B _375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2063_A wire2063/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input146_A la_iena_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_622_ _622_/A _622_/B vssd vssd vccd vccd _622_/X sky130_fd_sc_hd__and2_4
XFILLER_22_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input313_A la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__476__A_N _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__566__A _566_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_553_ _553_/A _553_/B vssd vssd vccd vccd _553_/X sky130_fd_sc_hd__and2_2
XTAP_3788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4008 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__285__B _285_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_484_ _612_/A _484_/B _484_/C vssd vssd vccd vccd _484_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2098 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3010 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output532_A wire1097/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1163_A wire1164/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1330_A _247_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1428_A wire1429/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] _207_/X vssd vssd vccd vccd _027_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1797_A wire1797/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1964_A wire1964/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput910 _121_/Y vssd vssd vccd vccd mprj_dat_i_core[7] sky130_fd_sc_hd__buf_8
Xoutput921 wire1202/X vssd vssd vccd vccd mprj_dat_o_user[17] sky130_fd_sc_hd__buf_8
Xoutput932 wire1162/X vssd vssd vccd vccd mprj_dat_o_user[27] sky130_fd_sc_hd__buf_8
Xoutput943 wire1229/X vssd vssd vccd vccd mprj_dat_o_user[8] sky130_fd_sc_hd__buf_8
XFILLER_47_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_4379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] _169_/X vssd vssd vccd vccd _153_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_25_2900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput954 output954/A vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_3_4120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1707 wire1707/A vssd vssd vccd vccd wire1707/X sky130_fd_sc_hd__buf_6
XFILLER_3_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1718 wire1718/A vssd vssd vccd vccd _351_/A sky130_fd_sc_hd__buf_6
XFILLER_41_2245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1729 wire1730/X vssd vssd vccd vccd _292_/A sky130_fd_sc_hd__buf_6
XTAP_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input263_A la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2180_A wire2181/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3238 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input430_A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__296__A _296_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_605_ _605_/A _605_/B vssd vssd vccd vccd _605_/X sky130_fd_sc_hd__and2_2
XFILLER_45_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_536_ _536_/A _536_/B vssd vssd vccd vccd _536_/X sky130_fd_sc_hd__and2_4
XFILLER_15_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_467_ _595_/A _467_/B _467_/C vssd vssd vccd vccd _467_/X sky130_fd_sc_hd__and3b_4
XFILLER_14_962 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_398_ _526_/A _398_/B _398_/C vssd vssd vccd vccd _398_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output482_A _486_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1009_A wire1010/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__462__C _462_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output747_A _622_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1280_A wire1281/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1378_A wire1378/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output914_A wire1223/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3818 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1712_A wire1712/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[7\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput740 _616_/X vssd vssd vccd vccd la_oenb_core[119] sky130_fd_sc_hd__buf_8
XFILLER_5_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput751 wire1039/X vssd vssd vccd vccd la_oenb_core[13] sky130_fd_sc_hd__buf_8
XFILLER_47_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput762 wire1029/X vssd vssd vccd vccd la_oenb_core[23] sky130_fd_sc_hd__buf_8
XFILLER_5_3514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput773 wire1024/X vssd vssd vccd vccd la_oenb_core[33] sky130_fd_sc_hd__buf_8
XFILLER_25_3464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput784 _540_/X vssd vssd vccd vccd la_oenb_core[43] sky130_fd_sc_hd__buf_8
XFILLER_40_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2205 wire2206/X vssd vssd vccd vccd wire2205/X sky130_fd_sc_hd__buf_6
Xoutput795 wire1005/X vssd vssd vccd vccd la_oenb_core[53] sky130_fd_sc_hd__buf_8
XFILLER_5_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1504 wire1504/A vssd vssd vccd vccd wire1504/X sky130_fd_sc_hd__buf_6
XFILLER_41_2042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1515 wire1516/X vssd vssd vccd vccd _317_/B sky130_fd_sc_hd__buf_6
Xwire1526 wire1526/A vssd vssd vccd vccd wire1526/X sky130_fd_sc_hd__buf_6
XFILLER_5_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1537 wire1537/A vssd vssd vccd vccd _577_/A sky130_fd_sc_hd__buf_6
XFILLER_5_2868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[7\]_B _170_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1548 wire1548/A vssd vssd vccd vccd _566_/A sky130_fd_sc_hd__buf_6
Xwire1559 _417_/A_N vssd vssd vccd vccd _545_/A sky130_fd_sc_hd__buf_6
XFILLER_3_3293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2026_A wire2026/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input109_A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_321_ _321_/A _321_/B vssd vssd vccd vccd _321_/X sky130_fd_sc_hd__and2_2
XTAP_1457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_252_ _252_/A _252_/B vssd vssd vccd vccd _252_/X sky130_fd_sc_hd__and2_4
XANTENNA__563__B _563_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_183_ _183_/A _183_/B vssd vssd vccd vccd _183_/X sky130_fd_sc_hd__and2_1
XANTENNA_input380_A la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input74_A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__457__C _457_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1126_A _387_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_360 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_519_ _519_/A _519_/B vssd vssd vccd vccd _519_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__473__B _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output864_A _329_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1495_A wire1496/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1662_A wire1662/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1927_A wire1927/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] _281_/X vssd vssd vccd vccd _101_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_3_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__383__B _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput570 _450_/X vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__buf_8
XFILLER_44_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput581 wire1075/X vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__buf_8
XFILLER_47_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2002 wire2002/A vssd vssd vccd vccd wire2002/X sky130_fd_sc_hd__buf_6
XFILLER_40_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput592 _083_/Y vssd vssd vccd vccd la_data_in_mprj[100] sky130_fd_sc_hd__buf_8
XFILLER_5_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2013 wire2013/A vssd vssd vccd vccd wire2013/X sky130_fd_sc_hd__buf_6
Xwire2024 wire2024/A vssd vssd vccd vccd _539_/B sky130_fd_sc_hd__buf_4
XFILLER_43_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2035 wire2035/A vssd vssd vccd vccd _515_/B sky130_fd_sc_hd__buf_6
Xwire1301 wire1302/X vssd vssd vccd vccd wire1301/X sky130_fd_sc_hd__buf_6
XFILLER_8_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2046 wire2046/A vssd vssd vccd vccd wire2046/X sky130_fd_sc_hd__buf_6
XFILLER_21_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1312 _287_/X vssd vssd vccd vccd wire1312/X sky130_fd_sc_hd__buf_8
Xwire2057 wire2057/A vssd vssd vccd vccd _501_/B sky130_fd_sc_hd__buf_6
Xwire2068 wire2068/A vssd vssd vccd vccd wire2068/X sky130_fd_sc_hd__buf_6
Xwire1323 _254_/X vssd vssd vccd vccd wire1323/X sky130_fd_sc_hd__buf_6
XFILLER_43_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1334 input99/X vssd vssd vccd vccd _439_/C sky130_fd_sc_hd__buf_6
Xwire2079 wire2080/X vssd vssd vccd vccd _492_/B sky130_fd_sc_hd__buf_6
XFILLER_19_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1345 wire1345/A vssd vssd vccd vccd wire1345/X sky130_fd_sc_hd__buf_6
XANTENNA__558__B _558_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1356 wire1357/X vssd vssd vccd vccd _340_/B sky130_fd_sc_hd__buf_6
XFILLER_5_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2143_A wire2143/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input226_A la_iena_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1367 wire1367/A vssd vssd vccd vccd _361_/B sky130_fd_sc_hd__buf_6
Xwire1378 wire1378/A vssd vssd vccd vccd _353_/B sky130_fd_sc_hd__buf_6
Xwire1389 wire1390/X vssd vssd vccd vccd _347_/B sky130_fd_sc_hd__buf_6
XFILLER_34_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__574__A _574_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_51_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__293__B _293_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_304_ _304_/A _304_/B vssd vssd vccd vccd _304_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_235_ _235_/A _235_/B vssd vssd vccd vccd _235_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_166_ _166_/A _166_/B vssd vssd vccd vccd _166_/X sky130_fd_sc_hd__and2_1
XFILLER_49_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_097_ _097_/A vssd vssd vccd vccd _097_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1076_A _459_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__468__B _468_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1890 wire1891/X vssd vssd vccd vccd wire1890/X sky130_fd_sc_hd__buf_6
XFILLER_37_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1410_A wire1411/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1508_A wire1508/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_190 _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1638 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1877_A wire1878/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4310 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4102 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput309 la_oenb_mprj[29] vssd vssd vccd vccd wire1574/A sky130_fd_sc_hd__buf_6
XFILLER_29_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__378__B _378_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_16_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_150 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_020_ _020_/A vssd vssd vccd vccd _020_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_14_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2093_A wire2093/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input176_A la_iena_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input343_A la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__569__A _569_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2699 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input37_A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1120 _393_/X vssd vssd vccd vccd wire1120/X sky130_fd_sc_hd__buf_6
XFILLER_19_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1131 _382_/X vssd vssd vccd vccd wire1131/X sky130_fd_sc_hd__buf_6
XFILLER_25_2390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__288__B _288_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1142 _372_/X vssd vssd vccd vccd wire1142/X sky130_fd_sc_hd__buf_6
XFILLER_40_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1153 _367_/X vssd vssd vccd vccd wire1153/X sky130_fd_sc_hd__buf_6
Xwire1164 wire1165/X vssd vssd vccd vccd wire1164/X sky130_fd_sc_hd__buf_6
XFILLER_5_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1175 wire1176/X vssd vssd vccd vccd wire1175/X sky130_fd_sc_hd__buf_6
XFILLER_5_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1186 wire1187/X vssd vssd vccd vccd wire1186/X sky130_fd_sc_hd__buf_8
XFILLER_1_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1197 _356_/X vssd vssd vccd vccd wire1197/X sky130_fd_sc_hd__buf_6
XFILLER_34_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_218_ _218_/A _218_/B vssd vssd vccd vccd _218_/X sky130_fd_sc_hd__and2_2
XFILLER_45_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output562_A _443_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_149_ _149_/A vssd vssd vccd vccd _149_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__470__C _470_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output827_A _579_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__382__A_N _510_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1008 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1360_A wire1361/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1458_A wire1459/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] _237_/X vssd vssd vccd vccd _057_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1625_A wire1625/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1994_A wire1995/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_684 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__380__C _380_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput106 la_data_out_mprj[77] vssd vssd vccd vccd wire1627/A sky130_fd_sc_hd__buf_6
XFILLER_41_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput117 la_data_out_mprj[87] vssd vssd vccd vccd wire1617/A sky130_fd_sc_hd__buf_6
XFILLER_2_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput128 la_data_out_mprj[97] vssd vssd vccd vccd _466_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput139 la_iena_mprj[106] vssd vssd vccd vccd _269_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2106_A wire2107/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1546 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input293_A la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__571__B _571_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_90 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_003_ _003_/A vssd vssd vccd vccd _003_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input460_A user_irq_ena[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__299__A _299_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1039_A _510_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1206_A wire1207/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3422 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output777_A _534_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__481__B _481_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output944_A wire1226/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1742_A wire1743/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__002__A _002_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] _263_/X vssd vssd vccd vccd wire993/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_39_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__391__B _391_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_4027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input139_A la_iena_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2056_A wire2056/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_621_ _621_/A _621_/B vssd vssd vccd vccd _621_/X sky130_fd_sc_hd__and2_4
XTAP_4468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1742 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_552_ _552_/A _552_/B vssd vssd vccd vccd _552_/X sky130_fd_sc_hd__and2_4
XANTENNA__566__B _566_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input306_A la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_483_ _611_/A _483_/B _483_/C vssd vssd vccd vccd _483_/X sky130_fd_sc_hd__and3b_4
XFILLER_44_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__582__A _582_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output525_A wire1104/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1156_A wire1157/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__420__A_N _420_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__476__B _476_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1323_A _254_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output894_A _135_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] _200_/X vssd vssd vccd vccd _020_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_23_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1692_A wire1693/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1957_A wire1958/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput900 _141_/Y vssd vssd vccd vccd mprj_dat_i_core[27] sky130_fd_sc_hd__buf_8
XFILLER_9_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput911 _122_/Y vssd vssd vccd vccd mprj_dat_i_core[8] sky130_fd_sc_hd__buf_8
XFILLER_25_4347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput922 wire1198/X vssd vssd vccd vccd mprj_dat_o_user[18] sky130_fd_sc_hd__buf_8
Xoutput933 wire1158/X vssd vssd vccd vccd mprj_dat_o_user[28] sky130_fd_sc_hd__buf_8
Xoutput944 wire1226/X vssd vssd vccd vccd mprj_dat_o_user[9] sky130_fd_sc_hd__buf_8
XFILLER_28_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput955 wire1307/X vssd vssd vccd vccd user_clock sky130_fd_sc_hd__buf_8
XFILLER_45_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[30\]_B _193_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1708 wire1708/A vssd vssd vccd vccd _360_/A sky130_fd_sc_hd__buf_6
XTAP_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1719 wire1719/A vssd vssd vccd vccd _350_/A sky130_fd_sc_hd__buf_4
XFILLER_45_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__386__B _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[97\]_B _260_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2173_A wire2174/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input256_A la_iena_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__443__A_N _571_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input423_A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__577__A _577_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_604_ _604_/A _604_/B vssd vssd vccd vccd _604_/X sky130_fd_sc_hd__and2_4
XTAP_4298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3962 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_716 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_535_ _535_/A _535_/B vssd vssd vccd vccd _535_/X sky130_fd_sc_hd__and2_1
XFILLER_35_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[88\]_B wire1326/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_466_ _594_/A _466_/B _466_/C vssd vssd vccd vccd _466_/X sky130_fd_sc_hd__and3b_4
XFILLER_53_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_397_ _525_/A _397_/B _397_/C vssd vssd vccd vccd _397_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output475_A wire1056/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output642_A _013_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1273_A _315_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1440_A wire1441/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1538_A wire1538/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_B wire1333/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__466__A_N _594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput730 wire1042/X vssd vssd vccd vccd la_oenb_core[10] sky130_fd_sc_hd__buf_8
XFILLER_9_3651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput741 wire1041/X vssd vssd vccd vccd la_oenb_core[11] sky130_fd_sc_hd__buf_8
Xoutput752 wire1038/X vssd vssd vccd vccd la_oenb_core[14] sky130_fd_sc_hd__buf_8
XFILLER_47_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput763 wire1028/X vssd vssd vccd vccd la_oenb_core[24] sky130_fd_sc_hd__buf_8
Xoutput774 wire1022/X vssd vssd vccd vccd la_oenb_core[34] sky130_fd_sc_hd__buf_8
XFILLER_5_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput785 wire1015/X vssd vssd vccd vccd la_oenb_core[44] sky130_fd_sc_hd__buf_8
Xwire2206 wire2207/X vssd vssd vccd vccd wire2206/X sky130_fd_sc_hd__buf_6
XFILLER_25_3476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput796 _551_/X vssd vssd vccd vccd la_oenb_core[54] sky130_fd_sc_hd__buf_8
XFILLER_48_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1505 wire1506/X vssd vssd vccd vccd _320_/B sky130_fd_sc_hd__buf_6
Xwire1516 wire1517/X vssd vssd vccd vccd wire1516/X sky130_fd_sc_hd__buf_6
XTAP_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2054 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1527 wire1527/A vssd vssd vccd vccd _596_/A sky130_fd_sc_hd__buf_6
XTAP_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1538 wire1538/A vssd vssd vccd vccd _576_/A sky130_fd_sc_hd__buf_6
XTAP_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1549 wire1549/A vssd vssd vccd vccd _565_/A sky130_fd_sc_hd__buf_6
XFILLER_38_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_320_ _320_/A _320_/B vssd vssd vccd vccd _320_/X sky130_fd_sc_hd__and2_4
XFILLER_42_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2019_A wire2019/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_251_ _251_/A _251_/B vssd vssd vccd vccd _251_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_270 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_182_ _182_/A _182_/B vssd vssd vccd vccd _182_/X sky130_fd_sc_hd__and2_2
XFILLER_49_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input373_A la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input67_A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__100__A _100_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_361 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_518_ _518_/A _518_/B vssd vssd vccd vccd _518_/X sky130_fd_sc_hd__and2_4
XTAP_2682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output592_A _083_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1119_A _394_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_449_ _577_/A _449_/B _449_/C vssd vssd vccd vccd _449_/X sky130_fd_sc_hd__and3b_4
XFILLER_15_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__489__A_N _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output857_A _323_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1488_A wire1489/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1655_A wire1656/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1534 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__383__C _383_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2590 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput560 _441_/X vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__buf_8
XFILLER_40_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput571 _451_/X vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__buf_8
XFILLER_43_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput582 wire1074/X vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__buf_8
XFILLER_44_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2003 wire2004/X vssd vssd vccd vccd _573_/B sky130_fd_sc_hd__buf_6
Xoutput593 _084_/Y vssd vssd vccd vccd la_data_in_mprj[101] sky130_fd_sc_hd__buf_8
XFILLER_8_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2014 wire2014/A vssd vssd vccd vccd _567_/B sky130_fd_sc_hd__buf_6
XFILLER_47_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2025 wire2025/A vssd vssd vccd vccd _535_/B sky130_fd_sc_hd__buf_6
XFILLER_47_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2036 wire2036/A vssd vssd vccd vccd _514_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2047 wire2048/X vssd vssd vccd vccd _507_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1302 _300_/X vssd vssd vccd vccd wire1302/X sky130_fd_sc_hd__buf_6
XFILLER_8_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2058 wire2059/X vssd vssd vccd vccd _500_/B sky130_fd_sc_hd__buf_6
Xwire1313 _286_/X vssd vssd vccd vccd wire1313/X sky130_fd_sc_hd__buf_6
Xwire2069 wire2070/X vssd vssd vccd vccd _495_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1324 _253_/X vssd vssd vccd vccd wire1324/X sky130_fd_sc_hd__buf_8
XFILLER_25_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1335 input97/X vssd vssd vccd vccd _438_/C sky130_fd_sc_hd__buf_6
XFILLER_21_2436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1346 wire1347/X vssd vssd vccd vccd _345_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1357 wire1357/A vssd vssd vccd vccd wire1357/X sky130_fd_sc_hd__buf_6
Xwire1368 wire1368/A vssd vssd vccd vccd _360_/B sky130_fd_sc_hd__buf_6
Xwire1379 wire1380/X vssd vssd vccd vccd _352_/B sky130_fd_sc_hd__buf_6
XFILLER_28_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input121_A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input219_A la_iena_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2136_A wire2136/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__574__B _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_B _290_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_303_ _303_/A _303_/B vssd vssd vccd vccd _303_/X sky130_fd_sc_hd__and2_1
XTAP_1288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_234_ _234_/A _234_/B vssd vssd vccd vccd _234_/X sky130_fd_sc_hd__and2_4
XFILLER_7_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__590__A _590_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_165_ _165_/A _165_/B vssd vssd vccd vccd _165_/X sky130_fd_sc_hd__and2_1
XFILLER_6_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[2\] mprj_dat_i_user[2] max_length1310/X vssd vssd vccd vccd _116_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_32_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_096_ _096_/A vssd vssd vccd vccd _096_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_powergood_check_mprj_vdd_logic1 output952/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_940 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__468__C _468_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output605_A _095_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1880 wire1881/X vssd vssd vccd vccd wire1880/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1236_A wire1237/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1891 wire1891/A vssd vssd vccd vccd wire1891/X sky130_fd_sc_hd__buf_6
XFILLER_0_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__484__B _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_B _281_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1403_A wire1404/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_180 _358_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_191 _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1772_A wire1772/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4322 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__005__A _005_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1270 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[27\]_A mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__378__C _378_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__394__B _394_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[109\]_B _272_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2086_A wire2087/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input169_A la_iena_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__569__B _569_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input336_A la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[18\]_A mprj_dat_i_user[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1110 _403_/X vssd vssd vccd vccd wire1110/X sky130_fd_sc_hd__buf_6
XFILLER_25_2380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1121 _392_/X vssd vssd vccd vccd wire1121/X sky130_fd_sc_hd__buf_6
Xwire1132 _381_/X vssd vssd vccd vccd wire1132/X sky130_fd_sc_hd__buf_6
XFILLER_5_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1143 _371_/X vssd vssd vccd vccd wire1143/X sky130_fd_sc_hd__buf_6
Xwire1154 wire1155/X vssd vssd vccd vccd wire1154/X sky130_fd_sc_hd__buf_8
XFILLER_1_2316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1165 _364_/X vssd vssd vccd vccd wire1165/X sky130_fd_sc_hd__buf_6
Xwire1176 wire1177/X vssd vssd vccd vccd wire1176/X sky130_fd_sc_hd__buf_6
XFILLER_38_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1187 wire1188/X vssd vssd vccd vccd wire1187/X sky130_fd_sc_hd__buf_6
XFILLER_5_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1198 wire1199/X vssd vssd vccd vccd wire1198/X sky130_fd_sc_hd__buf_8
XFILLER_53_3907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__585__A _585_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_217_ _217_/A _217_/B vssd vssd vccd vccd _217_/X sky130_fd_sc_hd__and2_1
XFILLER_10_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_148_ _148_/A vssd vssd vccd vccd _148_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output555_A _437_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_079_ _079_/A vssd vssd vccd vccd _079_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_wire1186_A wire1187/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output722_A _599_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__479__B _479_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1353_A wire1353/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] _230_/X vssd vssd vccd vccd _050_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_1_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1520_A wire1521/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1618_A wire1618/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1987_A wire1987/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire973_A wire973/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput107 la_data_out_mprj[78] vssd vssd vccd vccd wire1626/A sky130_fd_sc_hd__buf_6
XFILLER_22_3232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput118 la_data_out_mprj[88] vssd vssd vccd vccd wire1616/A sky130_fd_sc_hd__buf_6
XANTENNA__389__B _389_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput129 la_data_out_mprj[98] vssd vssd vccd vccd _467_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2001_A wire2002/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input286_A la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_80 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_002_ _002_/A vssd vssd vccd vccd _002_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_91 mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input453_A mprj_iena_wb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__299__B _299_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1101_A _412_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__481__C _481_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output937_A wire1146/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1470_A wire1471/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1568_A _405_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1735_A wire1736/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1902_A wire1903/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_620_ _620_/A _620_/B vssd vssd vccd vccd _620_/X sky130_fd_sc_hd__and2_4
XFILLER_22_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2049_A wire2050/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_551_ _551_/A _551_/B vssd vssd vccd vccd _551_/X sky130_fd_sc_hd__and2_4
XTAP_3768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input201_A la_iena_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_482_ _610_/A _482_/B _482_/C vssd vssd vccd vccd _482_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__372__A_N _500_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__582__B _582_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input97_A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__103__A _103_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3758 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output518_A wire1110/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput460 user_irq_ena[0] vssd vssd vccd vccd _291_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1051_A _499_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3632 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__492__B _492_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1685_A wire1685/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput901 _142_/Y vssd vssd vccd vccd mprj_dat_i_core[28] sky130_fd_sc_hd__buf_8
Xoutput912 _123_/Y vssd vssd vccd vccd mprj_dat_i_core[9] sky130_fd_sc_hd__buf_8
XANTENNA_wire1852_A wire1853/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput923 wire1194/X vssd vssd vccd vccd mprj_dat_o_user[19] sky130_fd_sc_hd__buf_8
XFILLER_28_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput934 wire1154/X vssd vssd vccd vccd mprj_dat_o_user[29] sky130_fd_sc_hd__buf_8
XFILLER_47_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput945 wire1294/X vssd vssd vccd vccd mprj_sel_o_user[0] sky130_fd_sc_hd__buf_8
Xoutput956 _297_/X vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__buf_8
XFILLER_45_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1709 wire1709/A vssd vssd vccd vccd _359_/A sky130_fd_sc_hd__buf_6
XFILLER_25_2968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__386__C _386_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__395__A_N _523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2642 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input151_A la_iena_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2166_A wire2166/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input249_A la_iena_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__577__B _577_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input416_A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_603_ _603_/A _603_/B vssd vssd vccd vccd _603_/X sky130_fd_sc_hd__and2_4
XTAP_4288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_534_ _534_/A _534_/B vssd vssd vccd vccd _534_/X sky130_fd_sc_hd__and2_4
XFILLER_15_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__593__A _593_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_465_ _593_/A _465_/B _465_/C vssd vssd vccd vccd _465_/X sky130_fd_sc_hd__and3b_4
XTAP_2897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_396_ _524_/A _396_/B _396_/C vssd vssd vccd vccd _396_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_3551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output468_A wire1062/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1099_A _414_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3923 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output635_A _007_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1266_A wire1267/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output802_A wire1048/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__487__B _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1433_A wire1434/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput290 la_oenb_mprj[127] vssd vssd vccd vccd wire1579/A sky130_fd_sc_hd__buf_6
XFILLER_3_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__008__A _008_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput720 _597_/X vssd vssd vccd vccd la_oenb_core[100] sky130_fd_sc_hd__buf_8
XFILLER_47_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput731 _607_/X vssd vssd vccd vccd la_oenb_core[110] sky130_fd_sc_hd__buf_8
Xoutput742 _617_/X vssd vssd vccd vccd la_oenb_core[120] sky130_fd_sc_hd__buf_8
XFILLER_9_3663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput753 wire1037/X vssd vssd vccd vccd la_oenb_core[15] sky130_fd_sc_hd__buf_8
XFILLER_43_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput764 wire1027/X vssd vssd vccd vccd la_oenb_core[25] sky130_fd_sc_hd__buf_8
XFILLER_47_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput775 _532_/X vssd vssd vccd vccd la_oenb_core[35] sky130_fd_sc_hd__buf_8
XFILLER_9_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput786 wire1013/X vssd vssd vccd vccd la_oenb_core[45] sky130_fd_sc_hd__buf_8
Xwire2207 wire2208/X vssd vssd vccd vccd wire2207/X sky130_fd_sc_hd__buf_6
Xoutput797 wire1004/X vssd vssd vccd vccd la_oenb_core[55] sky130_fd_sc_hd__buf_8
XFILLER_48_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1506 wire1507/X vssd vssd vccd vccd wire1506/X sky130_fd_sc_hd__buf_6
XFILLER_24_1018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1517 wire1517/A vssd vssd vccd vccd wire1517/X sky130_fd_sc_hd__buf_6
XFILLER_47_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1528 wire1528/A vssd vssd vccd vccd _595_/A sky130_fd_sc_hd__buf_6
XTAP_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1539 wire1539/A vssd vssd vccd vccd _575_/A sky130_fd_sc_hd__buf_8
XTAP_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__397__B _397_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_250_ _250_/A _250_/B vssd vssd vccd vccd _250_/X sky130_fd_sc_hd__and2_4
XFILLER_36_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_181_ _181_/A _181_/B vssd vssd vccd vccd _181_/X sky130_fd_sc_hd__and2_1
XFILLER_52_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input199_A la_iena_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__410__A_N _538_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input366_A la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_irq_gates\[1\] user_irq_core[1] _292_/X vssd vssd vccd vccd _112_/A sky130_fd_sc_hd__nand2_2
XFILLER_8_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__588__A _588_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_340 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_351 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_517_ _517_/A _517_/B vssd vssd vccd vccd _517_/X sky130_fd_sc_hd__and2_4
XTAP_2672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_362 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_448_ _576_/A _448_/B _448_/C vssd vssd vccd vccd _448_/X sky130_fd_sc_hd__and3b_4
XTAP_1982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output585_A wire1071/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3370 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_379_ _507_/A _379_/B _379_/C vssd vssd vccd vccd _379_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output752_A wire1038/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1383_A wire1384/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] _260_/X vssd vssd vccd vccd _080_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_3825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1648_A wire1649/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__498__A _498_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__433__A_N _561_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput550 _432_/X vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__buf_8
Xoutput561 _442_/X vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__buf_8
XFILLER_27_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput572 _452_/X vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__buf_8
XFILLER_47_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput583 wire1073/X vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__buf_8
Xwire2004 wire2004/A vssd vssd vccd vccd wire2004/X sky130_fd_sc_hd__buf_6
Xoutput594 _085_/Y vssd vssd vccd vccd la_data_in_mprj[102] sky130_fd_sc_hd__buf_8
XFILLER_5_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2015 wire2015/A vssd vssd vccd vccd _566_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2026 wire2026/A vssd vssd vccd vccd _531_/B sky130_fd_sc_hd__buf_6
Xwire2037 wire2038/X vssd vssd vccd vccd _513_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1303 wire1304/X vssd vssd vccd vccd wire1303/X sky130_fd_sc_hd__buf_6
Xwire2048 wire2048/A vssd vssd vccd vccd wire2048/X sky130_fd_sc_hd__buf_6
XFILLER_43_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__201__A _201_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2059 wire2059/A vssd vssd vccd vccd wire2059/X sky130_fd_sc_hd__buf_6
XFILLER_21_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1314 _277_/X vssd vssd vccd vccd wire1314/X sky130_fd_sc_hd__buf_6
Xwire1325 _252_/X vssd vssd vccd vccd wire1325/X sky130_fd_sc_hd__buf_8
XFILLER_25_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1336 input96/X vssd vssd vccd vccd _437_/C sky130_fd_sc_hd__buf_6
Xwire1347 wire1347/A vssd vssd vccd vccd wire1347/X sky130_fd_sc_hd__buf_6
XFILLER_3_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1358 wire1358/A vssd vssd vccd vccd _368_/B sky130_fd_sc_hd__buf_6
Xwire1369 wire1369/A vssd vssd vccd vccd _359_/B sky130_fd_sc_hd__buf_6
XFILLER_38_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2031_A wire2031/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input114_A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2129_A wire2129/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ _302_/A _302_/B vssd vssd vccd vccd _302_/X sky130_fd_sc_hd__and2_2
XTAP_1278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_233_ _233_/A _233_/B vssd vssd vccd vccd _233_/X sky130_fd_sc_hd__and2_2
XFILLER_50_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__590__B _590_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_164_ _164_/A _164_/B vssd vssd vccd vccd _164_/X sky130_fd_sc_hd__and2_1
XFILLER_10_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_095_ _095_/A vssd vssd vccd vccd _095_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_40_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1870 wire1870/A vssd vssd vccd vccd wire1870/X sky130_fd_sc_hd__buf_6
XANTENNA_output500_A wire1126/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1881 wire1882/X vssd vssd vccd vccd wire1881/X sky130_fd_sc_hd__buf_6
XFILLER_37_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1892 wire1893/X vssd vssd vccd vccd _618_/B sky130_fd_sc_hd__buf_6
XFILLER_20_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1131_A _382_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1229_A wire1230/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__456__A_N _584_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__484__C _484_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_181 _358_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_192 _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] _175_/X vssd vssd vccd vccd _159_/A
+ sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_gates\[25\] mprj_dat_i_user[25] _294_/X vssd vssd vccd vccd _139_/A sky130_fd_sc_hd__nand2_4
XFILLER_50_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1765_A wire1766/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1932_A wire1933/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2954 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__021__A _021_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[27\]_B _294_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] wire1313/X vssd vssd vccd vccd
+ wire981/A sky130_fd_sc_hd__nand2_2
XFILLER_2_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2079_A wire2080/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1100 _413_/X vssd vssd vccd vccd wire1100/X sky130_fd_sc_hd__buf_6
XANTENNA_user_wb_dat_gates\[18\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1111 _402_/X vssd vssd vccd vccd wire1111/X sky130_fd_sc_hd__buf_6
Xwire1122 _391_/X vssd vssd vccd vccd wire1122/X sky130_fd_sc_hd__buf_6
XFILLER_43_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input231_A la_iena_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1133 wire1134/X vssd vssd vccd vccd wire1133/X sky130_fd_sc_hd__buf_6
XANTENNA_input329_A la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__479__A_N _479_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1144 _370_/X vssd vssd vccd vccd wire1144/X sky130_fd_sc_hd__buf_6
Xwire1155 wire1156/X vssd vssd vccd vccd wire1155/X sky130_fd_sc_hd__buf_6
Xwire1166 wire1167/X vssd vssd vccd vccd wire1166/X sky130_fd_sc_hd__buf_8
XFILLER_47_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1177 _361_/X vssd vssd vccd vccd wire1177/X sky130_fd_sc_hd__buf_6
Xwire1188 wire1189/X vssd vssd vccd vccd wire1188/X sky130_fd_sc_hd__buf_6
XFILLER_5_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1199 wire1200/X vssd vssd vccd vccd wire1199/X sky130_fd_sc_hd__buf_6
XFILLER_38_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__585__B _585_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_216_ _216_/A _216_/B vssd vssd vccd vccd _216_/X sky130_fd_sc_hd__and2_2
XFILLER_11_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__106__A _106_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_147_ _147_/A vssd vssd vccd vccd _147_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1083 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_078_ _078_/A vssd vssd vccd vccd _078_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output548_A wire1079/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1081_A _428_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1179_A wire1180/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__479__C _479_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output715_A _080_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1346_A wire1347/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__495__B _495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1513_A wire1514/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1882_A wire1882/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire966_A wire966/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__016__A _016_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput108 la_data_out_mprj[79] vssd vssd vccd vccd wire1625/A sky130_fd_sc_hd__buf_6
XANTENNA__389__C _389_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput119 la_data_out_mprj[89] vssd vssd vccd vccd _458_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_642 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3936 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_70 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_001_ _001_/A vssd vssd vccd vccd _001_/Y sky130_fd_sc_hd__inv_2
XANTENNA_81 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_92 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input181_A la_iena_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2196_A wire2196/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input279_A la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input446_A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input42_A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__596__A _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output498_A wire1128/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1296_A wire1297/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output832_A _584_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1463_A wire1464/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1630_A wire1630/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1728_A wire1728/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput90 la_data_out_mprj[62] vssd vssd vccd vccd _431_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_550_ _550_/A _550_/B vssd vssd vccd vccd _550_/X sky130_fd_sc_hd__and2_2
XFILLER_17_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_940 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_481_ _609_/A _481_/B _481_/C vssd vssd vccd vccd _481_/X sky130_fd_sc_hd__and3b_1
XFILLER_16_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2111_A wire2111/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2209_A wire2209/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input396_A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput450 mprj_dat_o_core[7] vssd vssd vccd vccd wire1349/A sky130_fd_sc_hd__buf_6
XFILLER_23_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput461 user_irq_ena[1] vssd vssd vccd vccd _292_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1044_A _506_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3644 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1211_A wire1212/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output782_A wire1018/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1309_A _296_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__492__C _492_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3254 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1678_A wire1679/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput902 _143_/Y vssd vssd vccd vccd mprj_dat_i_core[29] sky130_fd_sc_hd__buf_8
XFILLER_29_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput913 wire1251/X vssd vssd vccd vccd mprj_dat_o_user[0] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput924 wire1249/X vssd vssd vccd vccd mprj_dat_o_user[1] sky130_fd_sc_hd__buf_8
XFILLER_9_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput935 wire1246/X vssd vssd vccd vccd mprj_dat_o_user[2] sky130_fd_sc_hd__buf_8
XFILLER_25_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput946 wire1289/X vssd vssd vccd vccd mprj_sel_o_user[1] sky130_fd_sc_hd__buf_8
Xoutput957 _111_/Y vssd vssd vccd vccd user_irq[0] sky130_fd_sc_hd__buf_8
XFILLER_3_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1845_A wire1845/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_4062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_442 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__204__A _204_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3090 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input144_A la_iena_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2061_A wire2061/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2159_A wire2160/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_602_ _602_/A _602_/B vssd vssd vccd vccd _602_/X sky130_fd_sc_hd__and2_4
XTAP_4278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input311_A la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input409_A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_533_ _533_/A _533_/B vssd vssd vccd vccd _533_/X sky130_fd_sc_hd__and2_4
XFILLER_2_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1574 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__593__B _593_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_464_ _592_/A _464_/B _464_/C vssd vssd vccd vccd _464_/X sky130_fd_sc_hd__and3b_4
XTAP_2898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_395_ _523_/A _395_/B _395_/C vssd vssd vccd vccd _395_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output530_A wire1099/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1161_A _365_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1259_A _322_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__487__C _487_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput280 la_oenb_mprj[118] vssd vssd vccd vccd wire1588/A sky130_fd_sc_hd__buf_6
Xinput291 la_oenb_mprj[12] vssd vssd vccd vccd _509_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] _205_/X vssd vssd vccd vccd _025_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_3430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1795_A wire1796/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1962_A wire1962/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput710 _075_/Y vssd vssd vccd vccd la_data_in_mprj[92] sky130_fd_sc_hd__buf_8
Xoutput721 _598_/X vssd vssd vccd vccd la_oenb_core[101] sky130_fd_sc_hd__buf_8
XANTENNA__024__A _024_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput732 _608_/X vssd vssd vccd vccd la_oenb_core[111] sky130_fd_sc_hd__buf_8
XFILLER_47_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput743 _618_/X vssd vssd vccd vccd la_oenb_core[121] sky130_fd_sc_hd__buf_8
Xoutput754 wire1036/X vssd vssd vccd vccd la_oenb_core[16] sky130_fd_sc_hd__buf_8
XFILLER_9_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput765 wire1026/X vssd vssd vccd vccd la_oenb_core[26] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] _167_/X vssd vssd vccd vccd _151_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput776 _533_/X vssd vssd vccd vccd la_oenb_core[36] sky130_fd_sc_hd__buf_8
XFILLER_28_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput787 _543_/X vssd vssd vccd vccd la_oenb_core[46] sky130_fd_sc_hd__buf_8
Xwire2208 wire2209/X vssd vssd vccd vccd wire2208/X sky130_fd_sc_hd__buf_6
Xoutput798 wire1002/X vssd vssd vccd vccd la_oenb_core[56] sky130_fd_sc_hd__buf_8
XFILLER_42_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1507 wire1508/X vssd vssd vccd vccd wire1507/X sky130_fd_sc_hd__buf_6
XFILLER_3_3241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1518 wire1519/X vssd vssd vccd vccd _316_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1529 wire1529/A vssd vssd vccd vccd _585_/A sky130_fd_sc_hd__buf_6
XTAP_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__397__C _397_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_751 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_180_ _180_/A _180_/B vssd vssd vccd vccd _180_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_294 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input261_A la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_622 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input359_A la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__588__B _588_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_330 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_341 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_352 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_516_ _516_/A _516_/B vssd vssd vccd vccd _516_/X sky130_fd_sc_hd__and2_4
XANTENNA_363 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__109__A _109_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_447_ _575_/A _447_/B _447_/C vssd vssd vccd vccd _447_/X sky130_fd_sc_hd__and3b_4
XTAP_1994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1007_A wire1008/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_378_ _506_/A _378_/B _378_/C vssd vssd vccd vccd _378_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output480_A _484_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output578_A wire1077/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output745_A _620_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__385__A_N _513_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1376_A wire1376/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output912_A _123_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__498__B _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1543_A wire1543/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1710_A wire1710/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1808_A wire1808/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire996_A _558_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__019__A _019_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput540 wire1089/X vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__buf_8
XFILLER_25_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput551 _433_/X vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__buf_8
XFILLER_9_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput562 _443_/X vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__buf_8
Xoutput573 _453_/X vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__buf_8
XFILLER_43_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput584 wire1072/X vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__buf_8
Xwire2005 wire2006/X vssd vssd vccd vccd _572_/B sky130_fd_sc_hd__buf_6
Xoutput595 _086_/Y vssd vssd vccd vccd la_data_in_mprj[103] sky130_fd_sc_hd__buf_8
XFILLER_21_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2016 wire2016/A vssd vssd vccd vccd _565_/B sky130_fd_sc_hd__buf_6
Xwire2027 wire2027/A vssd vssd vccd vccd _525_/B sky130_fd_sc_hd__buf_6
Xwire2038 wire2038/A vssd vssd vccd vccd wire2038/X sky130_fd_sc_hd__buf_6
XFILLER_25_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1304 wire1305/X vssd vssd vccd vccd wire1304/X sky130_fd_sc_hd__buf_6
Xwire2049 wire2050/X vssd vssd vccd vccd _506_/B sky130_fd_sc_hd__buf_6
Xwire1315 _270_/X vssd vssd vccd vccd wire1315/X sky130_fd_sc_hd__buf_6
XFILLER_8_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1326 _251_/X vssd vssd vccd vccd wire1326/X sky130_fd_sc_hd__buf_8
Xwire1337 input95/X vssd vssd vccd vccd _436_/C sky130_fd_sc_hd__buf_6
XFILLER_19_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1348 wire1349/X vssd vssd vccd vccd _344_/B sky130_fd_sc_hd__buf_6
XFILLER_28_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1359 wire1359/A vssd vssd vccd vccd _367_/B sky130_fd_sc_hd__buf_6
XFILLER_3_3093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_301_ _301_/A _301_/B vssd vssd vccd vccd _301_/X sky130_fd_sc_hd__and2_4
XTAP_1268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_232_ _232_/A _232_/B vssd vssd vccd vccd _232_/X sky130_fd_sc_hd__and2_2
XFILLER_24_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_163_ _163_/A vssd vssd vccd vccd _163_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input72_A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_094_ _094_/A vssd vssd vccd vccd _094_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__599__A _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1860 wire1860/A vssd vssd vccd vccd wire1860/X sky130_fd_sc_hd__buf_6
Xwire1871 wire1871/A vssd vssd vccd vccd _625_/A sky130_fd_sc_hd__buf_6
Xwire1882 wire1882/A vssd vssd vccd vccd wire1882/X sky130_fd_sc_hd__buf_6
XFILLER_24_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1893 wire1894/X vssd vssd vccd vccd wire1893/X sky130_fd_sc_hd__buf_6
XFILLER_18_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1124_A _389_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _221_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_171 _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_182 _358_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_193 _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output862_A wire1254/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[18\] mprj_dat_i_user[18] max_length1311/X vssd vssd vccd vccd
+ _132_/A sky130_fd_sc_hd__nand2_4
XFILLER_31_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1660_A wire1660/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1758_A wire1758/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__302__A _302_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1925_A wire1926/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] _279_/X vssd vssd vccd vccd _099_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_28_128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__400__A_N _400_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__212__A _212_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1101 _412_/X vssd vssd vccd vccd wire1101/X sky130_fd_sc_hd__buf_6
XFILLER_0_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1112 _401_/X vssd vssd vccd vccd wire1112/X sky130_fd_sc_hd__buf_6
Xwire1123 _390_/X vssd vssd vccd vccd wire1123/X sky130_fd_sc_hd__buf_6
XFILLER_5_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1134 _380_/X vssd vssd vccd vccd wire1134/X sky130_fd_sc_hd__buf_6
XFILLER_43_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1145 _369_/X vssd vssd vccd vccd wire1145/X sky130_fd_sc_hd__buf_6
Xwire1156 wire1157/X vssd vssd vccd vccd wire1156/X sky130_fd_sc_hd__buf_6
Xwire1167 wire1168/X vssd vssd vccd vccd wire1167/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2141_A wire2141/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input224_A la_iena_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1178 wire1179/X vssd vssd vccd vccd wire1178/X sky130_fd_sc_hd__buf_8
XFILLER_1_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1189 _358_/X vssd vssd vccd vccd wire1189/X sky130_fd_sc_hd__buf_6
XFILLER_28_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_215_ _215_/A _215_/B vssd vssd vccd vccd _215_/X sky130_fd_sc_hd__and2_2
XFILLER_11_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_146_ _146_/A vssd vssd vccd vccd _146_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_077_ _077_/A vssd vssd vccd vccd _077_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__122__A _122_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1074_A _461_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__423__A_N _551_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3779 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output610_A _100_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1241_A wire1242/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__495__C _495_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1690 wire1691/X vssd vssd vccd vccd _368_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1828 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1506_A wire1507/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput109 la_data_out_mprj[7] vssd vssd vccd vccd _376_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_654 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2206 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__207__A _207_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_60 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_000_ _000_/A vssd vssd vccd vccd _000_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_71 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_82 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_93 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2091_A wire2092/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input174_A la_iena_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2189_A wire2190/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_97 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__446__A_N _574_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input341_A la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input439_A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input35_A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__596__B _596_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output560_A _441_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output658_A _028_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_129_ _129_/A vssd vssd vccd vccd _129_/Y sky130_fd_sc_hd__inv_2
XANTENNA_wire1191_A wire1192/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1289_A wire1290/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output825_A _577_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1456_A wire1456/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] _235_/X vssd vssd vccd vccd _055_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1623_A wire1623/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1992_A wire1993/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__469__A_N _597_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput80 la_data_out_mprj[53] vssd vssd vccd vccd _422_/C sky130_fd_sc_hd__clkbuf_4
Xinput91 la_data_out_mprj[63] vssd vssd vccd vccd _432_/C sky130_fd_sc_hd__buf_4
XFILLER_43_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[33\]_B _196_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_480_ _608_/A _480_/B _480_/C vssd vssd vccd vccd _480_/X sky130_fd_sc_hd__and3b_2
XFILLER_26_952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1302 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3756 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input291_A la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input389_A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2506 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput440 mprj_dat_o_core[27] vssd vssd vccd vccd wire1364/A sky130_fd_sc_hd__buf_6
Xinput451 mprj_dat_o_core[8] vssd vssd vccd vccd wire1347/A sky130_fd_sc_hd__buf_6
Xinput462 user_irq_ena[2] vssd vssd vccd vccd _293_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1037_A _512_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1204_A _354_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output775_A _532_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output942_A wire1232/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput903 _116_/Y vssd vssd vccd vccd mprj_dat_i_core[2] sky130_fd_sc_hd__buf_8
Xoutput914 wire1223/X vssd vssd vccd vccd mprj_dat_o_user[10] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[15\]_B _178_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput925 wire1190/X vssd vssd vccd vccd mprj_dat_o_user[20] sky130_fd_sc_hd__buf_8
XFILLER_47_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput936 wire1150/X vssd vssd vccd vccd mprj_dat_o_user[30] sky130_fd_sc_hd__buf_8
XFILLER_9_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput947 wire1284/X vssd vssd vccd vccd mprj_sel_o_user[2] sky130_fd_sc_hd__buf_8
Xoutput958 _112_/Y vssd vssd vccd vccd user_irq[1] sky130_fd_sc_hd__buf_8
XFILLER_42_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1740_A wire1741/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1838_A wire1838/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__310__A _310_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_454 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2790 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__204__B _204_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input137_A la_iena_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_601_ _601_/A _601_/B vssd vssd vccd vccd _601_/X sky130_fd_sc_hd__and2_4
XTAP_4268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_532_ _532_/A _532_/B vssd vssd vccd vccd _532_/X sky130_fd_sc_hd__and2_4
XTAP_2822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input304_A la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_463_ _591_/A _463_/B _463_/C vssd vssd vccd vccd _463_/X sky130_fd_sc_hd__and3b_4
XTAP_2877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_394_ _522_/A _394_/B _394_/C vssd vssd vccd vccd _394_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output523_A wire1105/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__130__A _130_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1154_A wire1155/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput270 la_oenb_mprj[109] vssd vssd vccd vccd _478_/A_N sky130_fd_sc_hd__buf_6
XFILLER_20_3579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput281 la_oenb_mprj[119] vssd vssd vccd vccd wire1587/A sky130_fd_sc_hd__buf_6
XFILLER_7_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput292 la_oenb_mprj[13] vssd vssd vccd vccd _510_/A sky130_fd_sc_hd__buf_4
XFILLER_36_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1321_A _256_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1419_A wire1420/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] _198_/X vssd vssd vccd vccd _018_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_51_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1690_A wire1691/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1788_A wire1788/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__305__A _305_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1955_A wire1956/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput700 _066_/Y vssd vssd vccd vccd la_data_in_mprj[83] sky130_fd_sc_hd__buf_8
XFILLER_9_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput711 _076_/Y vssd vssd vccd vccd la_data_in_mprj[93] sky130_fd_sc_hd__buf_8
Xoutput722 _599_/X vssd vssd vccd vccd la_oenb_core[102] sky130_fd_sc_hd__buf_8
Xoutput733 _609_/X vssd vssd vccd vccd la_oenb_core[112] sky130_fd_sc_hd__buf_8
Xoutput744 _619_/X vssd vssd vccd vccd la_oenb_core[122] sky130_fd_sc_hd__buf_8
Xoutput755 wire1035/X vssd vssd vccd vccd la_oenb_core[17] sky130_fd_sc_hd__buf_8
XFILLER_47_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput766 _524_/X vssd vssd vccd vccd la_oenb_core[27] sky130_fd_sc_hd__buf_8
XFILLER_9_3687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput777 _534_/X vssd vssd vccd vccd la_oenb_core[37] sky130_fd_sc_hd__buf_8
XFILLER_5_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput788 _544_/X vssd vssd vccd vccd la_oenb_core[47] sky130_fd_sc_hd__buf_8
Xoutput799 _554_/X vssd vssd vccd vccd la_oenb_core[57] sky130_fd_sc_hd__buf_8
Xwire2209 wire2209/A vssd vssd vccd vccd wire2209/X sky130_fd_sc_hd__buf_6
XFILLER_28_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1508 wire1508/A vssd vssd vccd vccd wire1508/X sky130_fd_sc_hd__buf_6
XFILLER_28_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1519 wire1519/A vssd vssd vccd vccd wire1519/X sky130_fd_sc_hd__buf_6
XTAP_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_763 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__215__A _215_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1750 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2171_A wire2172/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input254_A la_iena_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_678 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input421_A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_320 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_331 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_342 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_515_ _515_/A _515_/B vssd vssd vccd vccd _515_/X sky130_fd_sc_hd__and2_2
XTAP_2652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_353 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_364 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_446_ _574_/A _446_/B _446_/C vssd vssd vccd vccd _446_/X sky130_fd_sc_hd__and3b_4
XTAP_1962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_377_ _505_/A _377_/B _377_/C vssd vssd vccd vccd _377_/X sky130_fd_sc_hd__and3b_4
XFILLER_48_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output473_A wire1057/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output640_A _012_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output738_A _614_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3755 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1271_A wire1272/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1369_A wire1369/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3310 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1536_A wire1536/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__035__A _035_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput530 wire1099/X vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__buf_8
Xoutput541 wire1087/X vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__buf_8
Xoutput552 _434_/X vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__buf_8
XFILLER_25_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput563 _444_/X vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__buf_8
XFILLER_47_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput574 _454_/X vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__buf_8
Xoutput585 wire1071/X vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__buf_8
Xwire2006 wire2006/A vssd vssd vccd vccd wire2006/X sky130_fd_sc_hd__buf_6
Xoutput596 _087_/Y vssd vssd vccd vccd la_data_in_mprj[104] sky130_fd_sc_hd__buf_8
Xwire2017 wire2017/A vssd vssd vccd vccd _564_/B sky130_fd_sc_hd__buf_6
XFILLER_5_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2028 wire2028/A vssd vssd vccd vccd _523_/B sky130_fd_sc_hd__buf_6
XFILLER_25_3287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2039 wire2039/A vssd vssd vccd vccd _512_/B sky130_fd_sc_hd__buf_6
Xwire1305 _299_/X vssd vssd vccd vccd wire1305/X sky130_fd_sc_hd__buf_6
Xwire1316 _266_/X vssd vssd vccd vccd wire1316/X sky130_fd_sc_hd__buf_6
Xwire1327 _250_/X vssd vssd vccd vccd wire1327/X sky130_fd_sc_hd__buf_8
XFILLER_3_3061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1338 input94/X vssd vssd vccd vccd _435_/C sky130_fd_sc_hd__buf_6
Xwire1349 wire1349/A vssd vssd vccd vccd wire1349/X sky130_fd_sc_hd__buf_6
XFILLER_41_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3924 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_858 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_300_ _300_/A _300_/B vssd vssd vccd vccd _300_/X sky130_fd_sc_hd__and2_4
XFILLER_42_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2017_A wire2017/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_4393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_231_ _231_/A _231_/B vssd vssd vccd vccd _231_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_162_ _162_/A vssd vssd vccd vccd _162_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_3534 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input371_A la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_093_ _093_/A vssd vssd vccd vccd _093_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_910 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input65_A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__599__B _599_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1850 wire1851/X vssd vssd vccd vccd _176_/A sky130_fd_sc_hd__buf_6
XFILLER_21_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1861 wire1861/A vssd vssd vccd vccd _169_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1872 wire1873/X vssd vssd vccd vccd _624_/B sky130_fd_sc_hd__buf_6
Xwire1883 wire1884/X vssd vssd vccd vccd _621_/B sky130_fd_sc_hd__buf_6
Xwire1894 wire1894/A vssd vssd vccd vccd wire1894/X sky130_fd_sc_hd__buf_6
XTAP_3150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 _210_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_161 _222_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_183 wire1459/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output590_A wire1136/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_194 _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1117_A _396_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output688_A _055_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_429_ _557_/A _429_/B _429_/C vssd vssd vccd vccd _429_/X sky130_fd_sc_hd__and3b_4
XTAP_1792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output855_A wire1260/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1486_A wire1487/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4242 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1653_A wire1653/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__302__B _302_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[0\]_A mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput1 caravel_clk vssd vssd vccd vccd _296_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_37_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] _272_/X vssd vssd vccd vccd _092_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_0_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__212__B _212_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1102 _411_/X vssd vssd vccd vccd wire1102/X sky130_fd_sc_hd__buf_6
XFILLER_5_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1113 _400_/X vssd vssd vccd vccd wire1113/X sky130_fd_sc_hd__buf_6
XFILLER_22_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1124 _389_/X vssd vssd vccd vccd wire1124/X sky130_fd_sc_hd__buf_6
Xwire1135 _379_/X vssd vssd vccd vccd wire1135/X sky130_fd_sc_hd__buf_6
XFILLER_19_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1146 wire1147/X vssd vssd vccd vccd wire1146/X sky130_fd_sc_hd__buf_8
XFILLER_5_2477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1157 _366_/X vssd vssd vccd vccd wire1157/X sky130_fd_sc_hd__buf_6
XFILLER_47_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1168 wire1169/X vssd vssd vccd vccd wire1168/X sky130_fd_sc_hd__buf_6
Xwire1179 wire1180/X vssd vssd vccd vccd wire1179/X sky130_fd_sc_hd__buf_6
XFILLER_19_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2134_A wire2134/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input217_A la_iena_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3754 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_214_ _214_/A _214_/B vssd vssd vccd vccd _214_/X sky130_fd_sc_hd__and2_2
XFILLER_7_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_145_ _145_/A vssd vssd vccd vccd _145_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[0\] mprj_dat_i_user[0] max_length1310/X vssd vssd vccd vccd _114_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_32_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_076_ _076_/A vssd vssd vccd vccd _076_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_4404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1067_A _468_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output603_A _093_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1680 wire1681/X vssd vssd vccd vccd _373_/B sky130_fd_sc_hd__buf_6
XFILLER_39_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1691 wire1691/A vssd vssd vccd vccd wire1691/X sky130_fd_sc_hd__buf_6
XFILLER_34_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1401_A wire1402/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[30\] mprj_dat_i_user[30] max_length1310/X vssd vssd vccd vccd
+ _144_/A sky130_fd_sc_hd__nand2_8
XFILLER_33_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1770_A wire1770/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1868_A wire1868/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__313__A _313_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__398__A_N _526_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__207__B _207_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_50 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_61 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_72 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_83 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_94 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2084_A wire2084/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input167_A la_iena_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input334_A la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input28_A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_128_ _128_/A vssd vssd vccd vccd _128_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output553_A _435_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__133__A _133_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_059_ _059_/A vssd vssd vccd vccd _059_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1184_A wire1185/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output720_A _597_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output818_A _571_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1351_A wire1351/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1449_A wire1450/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] _228_/X vssd vssd vccd vccd _048_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_40_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1616_A wire1616/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__308__A _308_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1985_A wire1985/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire971_A wire971/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput70 la_data_out_mprj[44] vssd vssd vccd vccd _413_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_8_4239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput81 la_data_out_mprj[54] vssd vssd vccd vccd _423_/C sky130_fd_sc_hd__clkbuf_4
Xinput92 la_data_out_mprj[64] vssd vssd vccd vccd _433_/C sky130_fd_sc_hd__buf_4
XFILLER_45_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__218__A _218_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1314 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__413__A_N _541_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input284_A la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input451_A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3936 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput430 mprj_dat_o_core[18] vssd vssd vccd vccd wire1376/A sky130_fd_sc_hd__buf_6
XFILLER_23_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput441 mprj_dat_o_core[28] vssd vssd vccd vccd wire1363/A sky130_fd_sc_hd__buf_6
XFILLER_48_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput452 mprj_dat_o_core[9] vssd vssd vccd vccd wire1345/A sky130_fd_sc_hd__buf_6
XFILLER_2_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output768_A _526_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1399_A wire1400/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output935_A wire1246/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput904 _144_/Y vssd vssd vccd vccd mprj_dat_i_core[30] sky130_fd_sc_hd__buf_8
Xoutput915 wire1220/X vssd vssd vccd vccd mprj_dat_o_user[11] sky130_fd_sc_hd__buf_8
XFILLER_28_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput926 wire1186/X vssd vssd vccd vccd mprj_dat_o_user[21] sky130_fd_sc_hd__buf_8
Xoutput937 wire1146/X vssd vssd vccd vccd mprj_dat_o_user[31] sky130_fd_sc_hd__buf_8
XFILLER_47_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput948 wire1280/X vssd vssd vccd vccd mprj_sel_o_user[3] sky130_fd_sc_hd__buf_8
XFILLER_25_3639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput959 _113_/Y vssd vssd vccd vccd user_irq[2] sky130_fd_sc_hd__buf_8
XTAP_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1733_A wire1734/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__310__B _310_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1900_A wire1901/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2302 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__436__A_N _564_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__038__A _038_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__501__A _501_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_600_ _600_/A _600_/B vssd vssd vccd vccd _600_/X sky130_fd_sc_hd__and2_4
XTAP_4258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2047_A wire2048/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_531_ _531_/A _531_/B vssd vssd vccd vccd _531_/X sky130_fd_sc_hd__and2_1
XTAP_2812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_462_ _590_/A _462_/B _462_/C vssd vssd vccd vccd _462_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_393_ _521_/A _393_/B _393_/C vssd vssd vccd vccd _393_/X sky130_fd_sc_hd__and3b_4
XFILLER_25_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input95_A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1707 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output516_A wire1112/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput260 la_oenb_mprj[0] vssd vssd vccd vccd _497_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput271 la_oenb_mprj[10] vssd vssd vccd vccd _507_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput282 la_oenb_mprj[11] vssd vssd vccd vccd _508_/A sky130_fd_sc_hd__buf_4
Xinput293 la_oenb_mprj[14] vssd vssd vccd vccd _511_/A sky130_fd_sc_hd__buf_4
XANTENNA_wire1147_A wire1148/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__459__A_N _587_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1314_A _277_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] _191_/X vssd vssd vccd vccd _011_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1683_A wire1683/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__305__B _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput701 _067_/Y vssd vssd vccd vccd la_data_in_mprj[84] sky130_fd_sc_hd__buf_8
Xoutput712 _077_/Y vssd vssd vccd vccd la_data_in_mprj[94] sky130_fd_sc_hd__buf_8
XANTENNA_wire1850_A wire1851/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput723 _600_/X vssd vssd vccd vccd la_oenb_core[103] sky130_fd_sc_hd__buf_8
XANTENNA_wire1948_A wire1949/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput734 _610_/X vssd vssd vccd vccd la_oenb_core[113] sky130_fd_sc_hd__buf_8
XFILLER_29_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput745 _620_/X vssd vssd vccd vccd la_oenb_core[123] sky130_fd_sc_hd__buf_8
Xoutput756 wire1034/X vssd vssd vccd vccd la_oenb_core[18] sky130_fd_sc_hd__buf_8
XFILLER_42_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput767 wire1025/X vssd vssd vccd vccd la_oenb_core[28] sky130_fd_sc_hd__buf_8
Xoutput778 wire1020/X vssd vssd vccd vccd la_oenb_core[38] sky130_fd_sc_hd__buf_8
Xoutput789 _545_/X vssd vssd vccd vccd la_oenb_core[48] sky130_fd_sc_hd__buf_8
XFILLER_42_4484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__321__A _321_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_powergood_check_mprj2_vdd_logic1 output954/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1509 wire1510/X vssd vssd vccd vccd _319_/B sky130_fd_sc_hd__buf_6
XTAP_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3863 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__215__B _215_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__231__A _231_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input247_A la_iena_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3834 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input414_A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_310 _437_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_321 wire1985/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_332 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_514_ _514_/A _514_/B vssd vssd vccd vccd _514_/X sky130_fd_sc_hd__and2_4
XTAP_2653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_343 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_354 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_365 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_445_ _573_/A _445_/B _445_/C vssd vssd vccd vccd _445_/X sky130_fd_sc_hd__and3b_4
XTAP_1963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ _504_/A _376_/B _376_/C vssd vssd vccd vccd _376_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output466_A wire1064/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1097_A _416_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output633_A _005_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__141__A _141_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1264_A wire1265/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output800_A wire1000/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1529_A wire1529/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1898_A wire1899/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__316__A _316_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput520 wire1108/X vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__buf_8
Xoutput531 wire1098/X vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__buf_8
XFILLER_44_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput542 wire1085/X vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__buf_8
XFILLER_9_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput553 _435_/X vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__buf_8
XFILLER_43_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput564 _445_/X vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__buf_8
Xoutput575 _455_/X vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__buf_8
XFILLER_47_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__051__A _051_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput586 wire1070/X vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__buf_8
Xwire2007 wire2008/X vssd vssd vccd vccd _571_/B sky130_fd_sc_hd__buf_6
Xoutput597 _088_/Y vssd vssd vccd vccd la_data_in_mprj[105] sky130_fd_sc_hd__buf_8
Xwire2018 wire2018/A vssd vssd vccd vccd _563_/B sky130_fd_sc_hd__buf_6
Xwire2029 wire2029/A vssd vssd vccd vccd _521_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1306 _298_/X vssd vssd vccd vccd wire1306/X sky130_fd_sc_hd__buf_6
XFILLER_5_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input2_A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1317 _262_/X vssd vssd vccd vccd wire1317/X sky130_fd_sc_hd__buf_6
XFILLER_47_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1328 _249_/X vssd vssd vccd vccd wire1328/X sky130_fd_sc_hd__buf_8
XFILLER_41_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1339 input93/X vssd vssd vccd vccd _434_/C sky130_fd_sc_hd__buf_6
XFILLER_3_3073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_230_ _230_/A _230_/B vssd vssd vccd vccd _230_/X sky130_fd_sc_hd__and2_2
XFILLER_23_583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__226__A _226_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_161_ _161_/A vssd vssd vccd vccd _161_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input197_A la_iena_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_092_ _092_/A vssd vssd vccd vccd _092_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input364_A la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input58_A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_966 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_454 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1840 wire1840/A vssd vssd vccd vccd _184_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1851 wire1851/A vssd vssd vccd vccd wire1851/X sky130_fd_sc_hd__buf_6
XFILLER_20_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1862 wire1862/A vssd vssd vccd vccd _168_/A sky130_fd_sc_hd__buf_6
XFILLER_1_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1873 wire1874/X vssd vssd vccd vccd wire1873/X sky130_fd_sc_hd__buf_6
Xwire1884 wire1885/X vssd vssd vccd vccd wire1884/X sky130_fd_sc_hd__buf_6
XTAP_3140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1895 wire1896/X vssd vssd vccd vccd _617_/B sky130_fd_sc_hd__buf_6
XTAP_3151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _210_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _222_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_173 _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_184 wire1461/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _524_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_428_ _556_/A _428_/B _428_/C vssd vssd vccd vccd _428_/X sky130_fd_sc_hd__and3b_4
XFILLER_18_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output583_A wire1073/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__136__A _136_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_359_ _359_/A _359_/B vssd vssd vccd vccd _359_/X sky130_fd_sc_hd__and2_1
XFILLER_35_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output750_A wire1040/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1381_A wire1382/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1479_A wire1480/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] wire1319/X vssd vssd vccd vccd wire962/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_44_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1646_A wire1647/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[0\]_B max_length1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput2 caravel_clk2 vssd vssd vccd vccd _297_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__046__A _046_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1103 _410_/X vssd vssd vccd vccd wire1103/X sky130_fd_sc_hd__buf_6
XFILLER_5_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1114 _399_/X vssd vssd vccd vccd wire1114/X sky130_fd_sc_hd__buf_6
XFILLER_48_929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1125 _388_/X vssd vssd vccd vccd wire1125/X sky130_fd_sc_hd__buf_6
XFILLER_9_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1136 _378_/X vssd vssd vccd vccd wire1136/X sky130_fd_sc_hd__buf_6
Xwire1147 wire1148/X vssd vssd vccd vccd wire1147/X sky130_fd_sc_hd__buf_6
Xwire1158 wire1159/X vssd vssd vccd vccd wire1158/X sky130_fd_sc_hd__buf_8
XFILLER_0_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1169 _363_/X vssd vssd vccd vccd wire1169/X sky130_fd_sc_hd__buf_6
XFILLER_38_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input112_A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_213_ _213_/A _213_/B vssd vssd vccd vccd _213_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_144_ _144_/A vssd vssd vccd vccd _144_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_075_ _075_/A vssd vssd vccd vccd _075_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_4541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__403__B _403_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1670 wire1671/X vssd vssd vccd vccd _377_/B sky130_fd_sc_hd__buf_6
XFILLER_20_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1681 wire1681/A vssd vssd vccd vccd wire1681/X sky130_fd_sc_hd__buf_6
XFILLER_18_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1692 wire1693/X vssd vssd vccd vccd _367_/A sky130_fd_sc_hd__buf_6
XFILLER_0_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1227_A wire1228/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output798_A wire1002/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] _173_/X vssd vssd vccd vccd _157_/A
+ sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_gates\[23\] mprj_dat_i_user[23] max_length1310/X vssd vssd vccd vccd
+ _137_/A sky130_fd_sc_hd__nand2_4
XFILLER_50_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1596_A _479_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1763_A wire1764/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__313__B _313_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1930_A wire1930/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] _284_/X vssd vssd vccd vccd _104_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_40 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_51 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_62 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_73 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_84 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_95 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__504__A _504_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2077_A wire2078/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input327_A la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_954 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__492__A_N _620_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_49_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_127_ _127_/A vssd vssd vccd vccd _127_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_058_ _058_/A vssd vssd vccd vccd _058_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output546_A wire1140/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output713_A _078_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1344_A wire1345/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2190 wire2190/A vssd vssd vccd vccd wire2190/X sky130_fd_sc_hd__buf_6
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] _221_/X vssd vssd vccd vccd _041_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_19_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1511_A wire1511/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__308__B _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1880_A wire1881/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1978_A wire1978/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire964_A wire964/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__324__A _324_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput60 la_data_out_mprj[35] vssd vssd vccd vccd _404_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput71 la_data_out_mprj[45] vssd vssd vccd vccd _414_/C sky130_fd_sc_hd__clkbuf_4
Xinput82 la_data_out_mprj[55] vssd vssd vccd vccd _424_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput93 la_data_out_mprj[65] vssd vssd vccd vccd input93/X sky130_fd_sc_hd__buf_6
XFILLER_41_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_792 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_4404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__234__A _234_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2194_A wire2194/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input277_A la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input444_A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input40_A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput420 mprj_cyc_o_core vssd vssd vccd vccd wire1397/A sky130_fd_sc_hd__buf_6
Xinput431 mprj_dat_o_core[19] vssd vssd vccd vccd wire1375/A sky130_fd_sc_hd__buf_6
XFILLER_40_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput442 mprj_dat_o_core[29] vssd vssd vccd vccd wire1362/A sky130_fd_sc_hd__buf_6
XANTENNA__400__C _400_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput453 mprj_iena_wb vssd vssd vccd vccd _294_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output496_A wire1130/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__144__A _144_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__388__A_N _516_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1294_A wire1295/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput905 _145_/Y vssd vssd vccd vccd mprj_dat_i_core[31] sky130_fd_sc_hd__buf_8
XFILLER_49_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput916 wire1217/X vssd vssd vccd vccd mprj_dat_o_user[12] sky130_fd_sc_hd__buf_8
XFILLER_29_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output830_A _582_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput927 wire1182/X vssd vssd vccd vccd mprj_dat_o_user[22] sky130_fd_sc_hd__buf_8
XFILLER_28_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput938 wire1244/X vssd vssd vccd vccd mprj_dat_o_user[3] sky130_fd_sc_hd__buf_8
XANTENNA_output928_A wire1178/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput949 wire1303/X vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__buf_8
XFILLER_45_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1461_A wire1461/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1559_A _417_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1726_A wire1727/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__054__A _054_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__501__B _501_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_530_ _530_/A _530_/B vssd vssd vccd vccd _530_/X sky130_fd_sc_hd__and2_4
XTAP_3558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__229__A _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_461_ _589_/A _461_/B _461_/C vssd vssd vccd vccd _461_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_392_ _520_/A _392_/B _392_/C vssd vssd vccd vccd _392_/X sky130_fd_sc_hd__and3b_4
XFILLER_17_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2207_A wire2208/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input394_A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input88_A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__411__B _411_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput250 la_iena_mprj[91] vssd vssd vccd vccd _254_/B sky130_fd_sc_hd__clkbuf_4
Xinput261 la_oenb_mprj[100] vssd vssd vccd vccd wire1607/A sky130_fd_sc_hd__buf_6
Xinput272 la_oenb_mprj[110] vssd vssd vccd vccd _479_/A_N sky130_fd_sc_hd__buf_6
Xinput283 la_oenb_mprj[120] vssd vssd vccd vccd wire1586/A sky130_fd_sc_hd__buf_6
XFILLER_23_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output509_A wire1118/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput294 la_oenb_mprj[15] vssd vssd vccd vccd _512_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1042_A wire1043/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__139__A _139_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output780_A wire1050/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1307_A wire1308/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output878_A wire1276/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2342 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1676_A wire1677/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput702 _068_/Y vssd vssd vccd vccd la_data_in_mprj[85] sky130_fd_sc_hd__buf_8
XFILLER_9_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput713 _078_/Y vssd vssd vccd vccd la_data_in_mprj[95] sky130_fd_sc_hd__buf_8
Xoutput724 _601_/X vssd vssd vccd vccd la_oenb_core[104] sky130_fd_sc_hd__buf_8
XFILLER_9_3645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput735 _611_/X vssd vssd vccd vccd la_oenb_core[114] sky130_fd_sc_hd__buf_8
XANTENNA__602__A _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput746 _621_/X vssd vssd vccd vccd la_oenb_core[124] sky130_fd_sc_hd__buf_8
XFILLER_29_2861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput757 wire1033/X vssd vssd vccd vccd la_oenb_core[19] sky130_fd_sc_hd__buf_8
XFILLER_47_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1843_A wire1843/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput768 _526_/X vssd vssd vccd vccd la_oenb_core[29] sky130_fd_sc_hd__buf_8
Xoutput779 wire1019/X vssd vssd vccd vccd la_oenb_core[39] sky130_fd_sc_hd__buf_8
XANTENNA__321__B _321_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__403__A_N _531_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__049__A _049_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__512__A _512_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__231__B _231_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3846 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input142_A la_iena_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2157_A wire2158/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input407_A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_300 wire1907/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_311 _341_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_322 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_513_ _513_/A _513_/B vssd vssd vccd vccd _513_/X sky130_fd_sc_hd__and2_4
XTAP_2632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_344 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_355 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_366 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_444_ _572_/A _444_/B _444_/C vssd vssd vccd vccd _444_/X sky130_fd_sc_hd__and3b_4
XTAP_2687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_375_ _503_/A _375_/B _375_/C vssd vssd vccd vccd _375_/X sky130_fd_sc_hd__and3b_4
XTAP_1997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__406__B _406_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__426__A_N _554_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1257_A _324_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1424_A wire1425/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] _203_/X vssd vssd vccd vccd _023_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_24_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1793_A wire1794/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__316__B _316_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1960_A wire1961/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[90\]_B wire1324/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput510 wire1117/X vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__buf_8
XANTENNA__332__A _332_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput521 wire1107/X vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__buf_8
XFILLER_9_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput532 wire1097/X vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__buf_8
XFILLER_44_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput543 wire1084/X vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__buf_8
Xoutput554 _436_/X vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] _165_/X vssd vssd vccd vccd _149_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput565 _446_/X vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__buf_8
XFILLER_5_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput576 _456_/X vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__buf_8
Xoutput587 wire1069/X vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__buf_8
Xwire2008 wire2008/A vssd vssd vccd vccd wire2008/X sky130_fd_sc_hd__buf_6
Xoutput598 _089_/Y vssd vssd vccd vccd la_data_in_mprj[106] sky130_fd_sc_hd__buf_8
Xwire2019 wire2019/A vssd vssd vccd vccd _562_/B sky130_fd_sc_hd__buf_6
XFILLER_25_3278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1307 wire1308/X vssd vssd vccd vccd wire1307/X sky130_fd_sc_hd__buf_6
XFILLER_3_3041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1318 _259_/X vssd vssd vccd vccd wire1318/X sky130_fd_sc_hd__buf_8
Xwire1329 _248_/X vssd vssd vccd vccd wire1329/X sky130_fd_sc_hd__buf_8
XFILLER_28_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__507__A _507_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_160_ _160_/A vssd vssd vccd vccd _160_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__226__B _226_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_091_ _091_/A vssd vssd vccd vccd _091_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_B _244_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__449__A_N _577_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__242__A _242_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input357_A la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1830 wire1830/A vssd vssd vccd vccd _190_/A sky130_fd_sc_hd__buf_6
XFILLER_19_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1841 wire1841/A vssd vssd vccd vccd _183_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1852 wire1853/X vssd vssd vccd vccd _175_/A sky130_fd_sc_hd__buf_6
Xwire1863 wire1864/X vssd vssd vccd vccd _167_/A sky130_fd_sc_hd__buf_6
Xwire1874 wire1875/X vssd vssd vccd vccd wire1874/X sky130_fd_sc_hd__buf_6
XFILLER_37_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1885 wire1885/A vssd vssd vccd vccd wire1885/X sky130_fd_sc_hd__buf_6
XTAP_3141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1896 wire1897/X vssd vssd vccd vccd wire1896/X sky130_fd_sc_hd__buf_6
XTAP_3152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _527_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_141 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_152 _212_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 _228_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _559_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_196 _618_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_427_ _555_/A _427_/B _427_/C vssd vssd vccd vccd _427_/X sky130_fd_sc_hd__and3b_4
XTAP_1783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_358_ _358_/A _358_/B vssd vssd vccd vccd _358_/X sky130_fd_sc_hd__and2_1
XFILLER_50_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1005_A wire1006/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output576_A _456_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_289_ _289_/A _289_/B vssd vssd vccd vccd _289_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[72\]_B _235_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output743_A _618_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1374_A wire1374/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] wire1326/X vssd vssd vccd vccd wire969/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_3587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1541_A wire1541/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1639_A wire1640/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput3 caravel_rstn vssd vssd vccd vccd input3/X sky130_fd_sc_hd__buf_6
XFILLER_4_2671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire994_A _587_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__327__A _327_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__062__A _062_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1104 _409_/X vssd vssd vccd vccd wire1104/X sky130_fd_sc_hd__buf_6
XFILLER_44_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1115 _398_/X vssd vssd vccd vccd wire1115/X sky130_fd_sc_hd__buf_6
Xwire1126 _387_/X vssd vssd vccd vccd wire1126/X sky130_fd_sc_hd__buf_6
XFILLER_5_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1137 _377_/X vssd vssd vccd vccd wire1137/X sky130_fd_sc_hd__buf_6
XFILLER_47_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1148 wire1149/X vssd vssd vccd vccd wire1148/X sky130_fd_sc_hd__buf_6
XFILLER_21_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1159 wire1160/X vssd vssd vccd vccd wire1159/X sky130_fd_sc_hd__buf_6
XFILLER_0_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2022_A wire2022/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__237__A _237_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_690 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_212_ _212_/A _212_/B vssd vssd vccd vccd _212_/X sky130_fd_sc_hd__and2_1
XFILLER_10_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_143_ _143_/A vssd vssd vccd vccd _143_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_52_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input70_A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_074_ _074_/A vssd vssd vccd vccd _074_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__403__C _403_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_230 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1660 wire1660/A vssd vssd vccd vccd wire1660/X sky130_fd_sc_hd__buf_6
Xwire1671 wire1671/A vssd vssd vccd vccd wire1671/X sky130_fd_sc_hd__buf_6
XFILLER_1_2844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1682 wire1683/X vssd vssd vccd vccd _372_/B sky130_fd_sc_hd__buf_6
Xwire1693 wire1693/A vssd vssd vccd vccd wire1693/X sky130_fd_sc_hd__buf_6
XFILLER_18_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1122_A _391_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output860_A wire1256/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[16\] mprj_dat_i_user[16] max_length1311/X vssd vssd vccd vccd
+ _130_/A sky130_fd_sc_hd__nand2_4
XFILLER_31_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1491_A wire1492/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire990 wire990/A vssd vssd vccd vccd _091_/A sky130_fd_sc_hd__buf_6
XFILLER_41_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1756_A wire1756/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__610__A _610_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_2503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1923_A wire1924/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] wire1314/X vssd vssd vccd vccd
+ wire985/A sky130_fd_sc_hd__nand2_4
XFILLER_39_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_602 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__057__A _057_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_30 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_41 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_52 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_63 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_74 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_85 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_B _199_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_96 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__504__B _504_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_B _283_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__520__A _520_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input222_A la_iena_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_126_ _126_/A vssd vssd vccd vccd _126_/Y sky130_fd_sc_hd__inv_2
XANTENNA__414__B _414_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_B _274_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_057_ _057_/A vssd vssd vccd vccd _057_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3671 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output539_A wire1090/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1072_A _463_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_4190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2180 wire2181/X vssd vssd vccd vccd _444_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2191 wire2191/A vssd vssd vccd vccd _438_/B sky130_fd_sc_hd__buf_6
XANTENNA_wire1337_A input95/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1490 wire1491/X vssd vssd vccd vccd _324_/B sky130_fd_sc_hd__buf_6
XFILLER_19_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1504_A wire1504/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[20\]_A mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__605__A _605_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1873_A wire1874/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__324__B _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[102\]_B _265_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput50 la_data_out_mprj[26] vssd vssd vccd vccd _395_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput61 la_data_out_mprj[36] vssd vssd vccd vccd _405_/C sky130_fd_sc_hd__clkbuf_4
Xinput72 la_data_out_mprj[46] vssd vssd vccd vccd _415_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput83 la_data_out_mprj[56] vssd vssd vccd vccd _425_/C sky130_fd_sc_hd__buf_4
XFILLER_28_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput94 la_data_out_mprj[66] vssd vssd vccd vccd input94/X sky130_fd_sc_hd__buf_6
XFILLER_28_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[11\]_A mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__515__A _515_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__234__B _234_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input172_A la_iena_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__250__A _250_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2266 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input437_A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput410 mprj_adr_o_core[2] vssd vssd vccd vccd wire1441/A sky130_fd_sc_hd__buf_6
Xinput421 mprj_dat_o_core[0] vssd vssd vccd vccd wire1393/A sky130_fd_sc_hd__buf_6
XFILLER_24_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input33_A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput432 mprj_dat_o_core[1] vssd vssd vccd vccd wire1374/A sky130_fd_sc_hd__buf_6
XFILLER_0_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput443 mprj_dat_o_core[2] vssd vssd vccd vccd wire1361/A sky130_fd_sc_hd__buf_6
XFILLER_40_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput454 mprj_sel_o_core[0] vssd vssd vccd vccd _301_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__409__B _409_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output489_A _492_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output656_A _026_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_109_ _109_/A vssd vssd vccd vccd _109_/Y sky130_fd_sc_hd__clkinv_2
Xoutput906 _117_/Y vssd vssd vccd vccd mprj_dat_i_core[3] sky130_fd_sc_hd__buf_8
Xoutput917 wire1214/X vssd vssd vccd vccd mprj_dat_o_user[13] sky130_fd_sc_hd__buf_8
XFILLER_45_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput928 wire1178/X vssd vssd vccd vccd mprj_dat_o_user[23] sky130_fd_sc_hd__buf_8
XFILLER_7_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1287_A wire1288/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput939 wire1241/X vssd vssd vccd vccd mprj_dat_o_user[4] sky130_fd_sc_hd__buf_8
XFILLER_45_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output823_A _576_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1454_A wire1455/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] _233_/X vssd vssd vccd vccd _053_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1621_A wire1621/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__319__B _319_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1990_A wire1991/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__335__A _335_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__A_N _610_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__070__A _070_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_460_ _588_/A _460_/B _460_/C vssd vssd vccd vccd _460_/X sky130_fd_sc_hd__and3b_4
XTAP_2847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__229__B _229_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_391_ _519_/A _391_/B _391_/C vssd vssd vccd vccd _391_/X sky130_fd_sc_hd__and3b_4
XFILLER_53_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2102_A wire2103/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__245__A _245_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input387_A la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4386 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput240 la_iena_mprj[82] vssd vssd vccd vccd _245_/B sky130_fd_sc_hd__buf_4
XFILLER_20_3549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput251 la_iena_mprj[92] vssd vssd vccd vccd _255_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput262 la_oenb_mprj[101] vssd vssd vccd vccd wire1606/A sky130_fd_sc_hd__buf_6
Xinput273 la_oenb_mprj[111] vssd vssd vccd vccd wire1595/A sky130_fd_sc_hd__buf_6
XFILLER_48_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput284 la_oenb_mprj[121] vssd vssd vccd vccd wire1585/A sky130_fd_sc_hd__buf_6
Xinput295 la_oenb_mprj[16] vssd vssd vccd vccd _513_/A sky130_fd_sc_hd__buf_4
XFILLER_18_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1035_A _514_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_589_ _589_/A _589_/B vssd vssd vccd vccd _589_/X sky130_fd_sc_hd__and2_4
XFILLER_18_3489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1202_A wire1203/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output773_A wire1024/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__155__A _155_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2354 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output940_A wire1238/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput703 _069_/Y vssd vssd vccd vccd la_data_in_mprj[86] sky130_fd_sc_hd__buf_8
XANTENNA_wire1571_A _400_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput714 _079_/Y vssd vssd vccd vccd la_data_in_mprj[96] sky130_fd_sc_hd__buf_8
XANTENNA_wire1669_A wire1669/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput725 _602_/X vssd vssd vccd vccd la_oenb_core[105] sky130_fd_sc_hd__buf_8
XFILLER_47_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput736 _612_/X vssd vssd vccd vccd la_oenb_core[115] sky130_fd_sc_hd__buf_8
XANTENNA__602__B _602_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput747 _622_/X vssd vssd vccd vccd la_oenb_core[125] sky130_fd_sc_hd__buf_8
Xoutput758 wire1052/X vssd vssd vccd vccd la_oenb_core[1] sky130_fd_sc_hd__buf_8
XFILLER_42_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput769 wire1051/X vssd vssd vccd vccd la_oenb_core[2] sky130_fd_sc_hd__buf_8
XFILLER_47_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1836_A wire1836/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__065__A _065_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__512__B _512_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2052_A wire2052/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input135_A la_iena_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__378__A_N _506_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_301 wire1951/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_512_ _512_/A _512_/B vssd vssd vccd vccd _512_/X sky130_fd_sc_hd__and2_4
XFILLER_19_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 _351_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_323 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input302_A la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_334 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_345 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_356 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_443_ _571_/A _443_/B _443_/C vssd vssd vccd vccd _443_/X sky130_fd_sc_hd__and3b_4
XTAP_2677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_374_ _502_/A _374_/B _374_/C vssd vssd vccd vccd _374_/X sky130_fd_sc_hd__and3b_4
XTAP_1987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output521_A wire1107/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1152_A wire1153/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1417_A wire1418/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] _196_/X vssd vssd vccd vccd _016_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_51_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__613__A _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1953_A wire1954/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput500 wire1126/X vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__buf_8
Xoutput511 wire1116/X vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__buf_8
Xoutput522 wire1106/X vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__buf_8
XANTENNA__332__B _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput533 wire1096/X vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__buf_8
XFILLER_47_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput544 wire1082/X vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__buf_8
Xoutput555 _437_/X vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__buf_8
XFILLER_47_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput566 _447_/X vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__buf_8
XANTENNA_user_wb_dat_gates\[3\]_A mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput577 _457_/X vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__buf_8
XFILLER_5_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput588 wire1068/X vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__buf_8
Xwire2009 wire2009/A vssd vssd vccd vccd _570_/B sky130_fd_sc_hd__buf_6
Xoutput599 _090_/Y vssd vssd vccd vccd la_data_in_mprj[107] sky130_fd_sc_hd__buf_8
XFILLER_42_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1308 wire1309/X vssd vssd vccd vccd wire1308/X sky130_fd_sc_hd__buf_6
XFILLER_25_2578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1319 _258_/X vssd vssd vccd vccd wire1319/X sky130_fd_sc_hd__buf_6
XFILLER_25_2589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__507__B _507_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_090_ _090_/A vssd vssd vccd vccd _090_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__523__A _523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input252_A la_iena_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1820 wire1820/A vssd vssd vccd vccd _206_/A sky130_fd_sc_hd__buf_6
Xwire1831 wire1832/X vssd vssd vccd vccd _189_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1842 wire1842/A vssd vssd vccd vccd _329_/A sky130_fd_sc_hd__buf_6
XFILLER_21_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1853 wire1853/A vssd vssd vccd vccd wire1853/X sky130_fd_sc_hd__buf_6
Xwire1864 wire1864/A vssd vssd vccd vccd wire1864/X sky130_fd_sc_hd__buf_6
XFILLER_19_836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1875 wire1875/A vssd vssd vccd vccd wire1875/X sky130_fd_sc_hd__buf_6
XFILLER_18_324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1886 wire1887/X vssd vssd vccd vccd _620_/B sky130_fd_sc_hd__buf_6
XFILLER_37_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1897 wire1897/A vssd vssd vccd vccd wire1897/X sky130_fd_sc_hd__buf_6
XTAP_3153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _527_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_142 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _212_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_164 _228_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_175 _341_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_186 _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_426_ _554_/A _426_/B _426_/C vssd vssd vccd vccd _426_/X sky130_fd_sc_hd__and3b_4
XTAP_1773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__417__B _417_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_197 _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ _357_/A _357_/B vssd vssd vccd vccd _357_/X sky130_fd_sc_hd__and2_1
XFILLER_32_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_288_ _288_/A _288_/B vssd vssd vccd vccd _288_/X sky130_fd_sc_hd__and2_4
XANTENNA_output471_A wire1059/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output569_A _449_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_740 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output736_A _612_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1367_A wire1367/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1534_A wire1534/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput4 la_data_out_mprj[0] vssd vssd vccd vccd _369_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_20_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1701_A wire1701/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__608__A _608_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__327__B _327_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire987_A wire987/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__343__A _343_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1105 _408_/X vssd vssd vccd vccd wire1105/X sky130_fd_sc_hd__buf_6
XFILLER_40_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1116 _397_/X vssd vssd vccd vccd wire1116/X sky130_fd_sc_hd__buf_6
Xwire1127 _386_/X vssd vssd vccd vccd wire1127/X sky130_fd_sc_hd__buf_6
XFILLER_9_1893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1138 _376_/X vssd vssd vccd vccd wire1138/X sky130_fd_sc_hd__buf_6
Xwire1149 _368_/X vssd vssd vccd vccd wire1149/X sky130_fd_sc_hd__buf_6
XFILLER_27_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__518__A _518_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__237__B _237_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2015_A wire2015/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__416__A_N _416_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_211_ _211_/A _211_/B vssd vssd vccd vccd _211_/X sky130_fd_sc_hd__and2_1
XFILLER_49_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_142_ _142_/A vssd vssd vccd vccd _142_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__253__A _253_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_073_ _073_/A vssd vssd vccd vccd _073_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input63_A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1650 wire1651/X vssd vssd vccd vccd _386_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1661 wire1662/X vssd vssd vccd vccd _381_/B sky130_fd_sc_hd__buf_6
XFILLER_47_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1672 wire1673/X vssd vssd vccd vccd _376_/B sky130_fd_sc_hd__buf_6
Xwire1683 wire1683/A vssd vssd vccd vccd wire1683/X sky130_fd_sc_hd__buf_6
XFILLER_19_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1694 wire1695/X vssd vssd vccd vccd _366_/A sky130_fd_sc_hd__buf_6
XFILLER_19_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1115_A _398_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output686_A _053_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_409_ _409_/A_N _409_/B _409_/C vssd vssd vccd vccd _409_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output853_A wire1262/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__163__A _163_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1484_A wire1484/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire980 wire980/A vssd vssd vccd vccd _109_/A sky130_fd_sc_hd__buf_6
XFILLER_31_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire991 wire991/A vssd vssd vccd vccd _090_/A sky130_fd_sc_hd__buf_6
XFILLER_6_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1749_A wire1750/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__610__B _610_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1916_A wire1917/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] wire1315/X vssd vssd vccd vccd
+ wire991/A sky130_fd_sc_hd__nand2_1
XFILLER_53_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__439__A_N _567_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__338__A _338_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_20 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_31 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_42 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_53 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_64 mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_75 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__073__A _073_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_86 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_97 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__520__B _520_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3750 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input215_A la_iena_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2132_A wire2132/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__248__A _248_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_125_ _125_/A vssd vssd vccd vccd _125_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__414__C _414_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_056_ _056_/A vssd vssd vccd vccd _056_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__430__B _430_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_4055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3490 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1065_A _470_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2170 wire2170/A vssd vssd vccd vccd wire2170/X sky130_fd_sc_hd__buf_6
XFILLER_21_3271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2181 wire2181/A vssd vssd vccd vccd wire2181/X sky130_fd_sc_hd__buf_6
Xwire2192 wire2192/A vssd vssd vccd vccd _437_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1480 wire1481/X vssd vssd vccd vccd wire1480/X sky130_fd_sc_hd__buf_6
Xwire1491 wire1492/X vssd vssd vccd vccd wire1491/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1232_A wire1233/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[20\]_B _294_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1699_A wire1699/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__605__B _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput40 la_data_out_mprj[17] vssd vssd vccd vccd _386_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1866_A wire1866/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput51 la_data_out_mprj[27] vssd vssd vccd vccd _396_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput62 la_data_out_mprj[37] vssd vssd vccd vccd _406_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput73 la_data_out_mprj[47] vssd vssd vccd vccd _416_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput84 la_data_out_mprj[57] vssd vssd vccd vccd _426_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_7_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput95 la_data_out_mprj[67] vssd vssd vccd vccd input95/X sky130_fd_sc_hd__buf_6
XFILLER_45_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__621__A _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__340__B _340_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__068__A _068_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[11\]_B _294_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__515__B _515_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__531__A _531_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input165_A la_iena_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2082_A wire2083/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2278 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput400 mprj_adr_o_core[20] vssd vssd vccd vccd wire1484/A sky130_fd_sc_hd__buf_6
XFILLER_2_4353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput411 mprj_adr_o_core[30] vssd vssd vccd vccd wire1436/A sky130_fd_sc_hd__buf_6
XFILLER_40_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput422 mprj_dat_o_core[10] vssd vssd vccd vccd wire1390/A sky130_fd_sc_hd__buf_6
XFILLER_7_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input332_A la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput433 mprj_dat_o_core[20] vssd vssd vccd vccd wire1371/A sky130_fd_sc_hd__buf_6
XFILLER_48_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput444 mprj_dat_o_core[30] vssd vssd vccd vccd wire1359/A sky130_fd_sc_hd__buf_6
XFILLER_0_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput455 mprj_sel_o_core[1] vssd vssd vccd vccd _302_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input26_A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__409__C _409_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3362 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__425__B _425_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_108_ _108_/A vssd vssd vccd vccd _108_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput907 _118_/Y vssd vssd vccd vccd mprj_dat_i_core[4] sky130_fd_sc_hd__buf_8
XFILLER_49_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output551_A _433_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput918 wire1211/X vssd vssd vccd vccd mprj_dat_o_user[14] sky130_fd_sc_hd__buf_8
Xoutput929 wire1174/X vssd vssd vccd vccd mprj_dat_o_user[24] sky130_fd_sc_hd__buf_8
XANTENNA_output649_A _020_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_039_ _039_/A vssd vssd vccd vccd _039_/Y sky130_fd_sc_hd__inv_2
XANTENNA_wire1182_A wire1183/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output816_A _569_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1447_A wire1448/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] _226_/X vssd vssd vccd vccd _046_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_36_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__616__A _616_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1983_A wire1983/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__335__B _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__351__A _351_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_390_ _518_/A _390_/B _390_/C vssd vssd vccd vccd _390_/X sky130_fd_sc_hd__and3b_4
XFILLER_52_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__526__A _526_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__245__B _245_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input282_A la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__261__A _261_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4354 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput230 la_iena_mprj[73] vssd vssd vccd vccd _236_/B sky130_fd_sc_hd__clkbuf_4
Xinput241 la_iena_mprj[83] vssd vssd vccd vccd _246_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput252 la_iena_mprj[93] vssd vssd vccd vccd _256_/B sky130_fd_sc_hd__clkbuf_4
Xinput263 la_oenb_mprj[102] vssd vssd vccd vccd wire1605/A sky130_fd_sc_hd__buf_6
Xinput274 la_oenb_mprj[112] vssd vssd vccd vccd wire1594/A sky130_fd_sc_hd__buf_6
XFILLER_49_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput285 la_oenb_mprj[122] vssd vssd vccd vccd wire1584/A sky130_fd_sc_hd__buf_6
XFILLER_18_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput296 la_oenb_mprj[17] vssd vssd vccd vccd _514_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_588_ _588_/A _588_/B vssd vssd vccd vccd _588_/X sky130_fd_sc_hd__and2_4
XFILLER_34_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_970 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output766_A _524_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1397_A wire1397/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1080 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output933_A wire1158/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput704 _070_/Y vssd vssd vccd vccd la_data_in_mprj[87] sky130_fd_sc_hd__buf_8
XFILLER_29_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput715 _080_/Y vssd vssd vccd vccd la_data_in_mprj[97] sky130_fd_sc_hd__buf_8
XANTENNA__171__A _171_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput726 _603_/X vssd vssd vccd vccd la_oenb_core[106] sky130_fd_sc_hd__buf_8
XFILLER_42_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput737 _613_/X vssd vssd vccd vccd la_oenb_core[116] sky130_fd_sc_hd__buf_8
XFILLER_47_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1564_A _412_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput748 _623_/X vssd vssd vccd vccd la_oenb_core[126] sky130_fd_sc_hd__buf_8
XFILLER_7_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput759 wire1032/X vssd vssd vccd vccd la_oenb_core[20] sky130_fd_sc_hd__buf_8
XFILLER_42_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1731_A wire1731/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1829_A wire1829/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__346__A _346_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__081__A _081_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_506 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input128_A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2045_A wire2046/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_302 wire1954/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_511_ _511_/A _511_/B vssd vssd vccd vccd _511_/X sky130_fd_sc_hd__and2_4
XTAP_3368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_313 wire1885/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_335 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_357 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ _570_/A _442_/B _442_/C vssd vssd vccd vccd _442_/X sky130_fd_sc_hd__and3b_4
XFILLER_19_3788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__256__A _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_373_ _501_/A _373_/B _373_/C vssd vssd vccd vccd _373_/X sky130_fd_sc_hd__and3b_4
XFILLER_39_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input93_A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[9\] mprj_dat_i_user[9] _294_/X vssd vssd vccd vccd _123_/A sky130_fd_sc_hd__nand2_2
XFILLER_29_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__422__C _422_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output514_A wire1114/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1145_A _369_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1312_A _287_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__472__A_N _472_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__166__A _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] _189_/X vssd vssd vccd vccd _009_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_14_2417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1681_A wire1681/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1779_A wire1779/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__613__B _613_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput501 wire1125/X vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__buf_8
Xoutput512 wire1115/X vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__buf_8
XFILLER_5_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput523 wire1105/X vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__buf_8
XFILLER_25_3203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput534 wire1095/X vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__buf_8
XFILLER_44_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1946_A wire1947/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput545 wire1081/X vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__buf_8
XFILLER_25_3236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput556 _438_/X vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__buf_8
XANTENNA_user_wb_dat_gates\[3\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput567 _448_/X vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__buf_8
XFILLER_5_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput578 wire1077/X vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__buf_8
Xoutput589 wire1067/X vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__buf_8
XFILLER_47_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1309 _296_/X vssd vssd vccd vccd wire1309/X sky130_fd_sc_hd__buf_6
XFILLER_38_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_358 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_4391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__076__A _076_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__523__B _523_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2162_A wire2163/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input245_A la_iena_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1810 wire1810/A vssd vssd vccd vccd _233_/A sky130_fd_sc_hd__buf_6
XFILLER_41_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1821 wire1821/A vssd vssd vccd vccd _205_/A sky130_fd_sc_hd__buf_6
Xwire1832 wire1832/A vssd vssd vccd vccd wire1832/X sky130_fd_sc_hd__buf_6
XFILLER_46_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1843 wire1843/A vssd vssd vccd vccd _182_/A sky130_fd_sc_hd__buf_6
XFILLER_21_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1854 wire1855/X vssd vssd vccd vccd _174_/A sky130_fd_sc_hd__buf_6
XTAP_3110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1865 wire1866/X vssd vssd vccd vccd _166_/A sky130_fd_sc_hd__buf_6
XTAP_3121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input412_A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1876 wire1877/X vssd vssd vccd vccd _623_/B sky130_fd_sc_hd__buf_6
XFILLER_46_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1887 wire1888/X vssd vssd vccd vccd wire1887/X sky130_fd_sc_hd__buf_6
XANTENNA__495__A_N _623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1898 wire1899/X vssd vssd vccd vccd _616_/B sky130_fd_sc_hd__buf_6
XFILLER_19_4253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 _547_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_154 _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _228_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _342_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_187 _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_425_ _553_/A _425_/B _425_/C vssd vssd vccd vccd _425_/X sky130_fd_sc_hd__and3b_2
XTAP_2497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__417__C _417_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_356_ _356_/A _356_/B vssd vssd vccd vccd _356_/X sky130_fd_sc_hd__and2_1
XFILLER_31_2027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_287_ _287_/A _287_/B vssd vssd vccd vccd _287_/X sky130_fd_sc_hd__and2_2
XFILLER_31_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__433__B _433_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output464_A wire1066/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1095_A _418_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output729_A _606_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1262_A wire1263/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput5 la_data_out_mprj[100] vssd vssd vccd vccd _469_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__608__B _608_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1896_A wire1897/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__624__A _624_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__343__B _343_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1106 _407_/X vssd vssd vccd vccd wire1106/X sky130_fd_sc_hd__buf_6
Xwire1117 _396_/X vssd vssd vccd vccd wire1117/X sky130_fd_sc_hd__buf_6
Xwire1128 _385_/X vssd vssd vccd vccd wire1128/X sky130_fd_sc_hd__buf_6
XFILLER_38_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1139 _375_/X vssd vssd vccd vccd wire1139/X sky130_fd_sc_hd__buf_6
XFILLER_19_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4426 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__518__B _518_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_210_ _210_/A _210_/B vssd vssd vccd vccd _210_/X sky130_fd_sc_hd__and2_1
XFILLER_51_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__534__A _534_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
X_141_ _141_/A vssd vssd vccd vccd _141_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_49_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input195_A la_iena_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__253__B _253_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_072_ _072_/A vssd vssd vccd vccd _072_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_2645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input362_A la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input56_A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1640 wire1640/A vssd vssd vccd vccd wire1640/X sky130_fd_sc_hd__buf_6
XFILLER_1_2824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1651 wire1651/A vssd vssd vccd vccd wire1651/X sky130_fd_sc_hd__buf_6
XFILLER_5_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1662 wire1662/A vssd vssd vccd vccd wire1662/X sky130_fd_sc_hd__buf_6
XFILLER_19_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1673 wire1673/A vssd vssd vccd vccd wire1673/X sky130_fd_sc_hd__buf_6
XFILLER_47_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1684 wire1685/X vssd vssd vccd vccd _371_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1695 wire1695/A vssd vssd vccd vccd wire1695/X sky130_fd_sc_hd__buf_6
XFILLER_46_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__428__B _428_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ _536_/A _408_/B _408_/C vssd vssd vccd vccd _408_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output581_A wire1075/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1108_A _405_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_32_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_339_ _339_/A _339_/B vssd vssd vccd vccd _339_/X sky130_fd_sc_hd__and2_1
XFILLER_35_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire970 wire970/A vssd vssd vccd vccd _070_/A sky130_fd_sc_hd__buf_6
XANTENNA_output846_A wire1044/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire981 wire981/A vssd vssd vccd vccd _106_/A sky130_fd_sc_hd__buf_6
Xwire992 wire992/A vssd vssd vccd vccd _086_/A sky130_fd_sc_hd__buf_6
XFILLER_45_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1477_A wire1478/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] wire1321/X vssd vssd vccd vccd wire964/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_41_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1644_A wire1644/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1811_A wire1811/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1909_A wire1910/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__619__A _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__338__B _338_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_10 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_21 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_32 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__354__A _354_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_43 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_54 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_65 mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_76 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_87 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_98 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__529__A _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__248__B _248_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input110_A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2125_A wire2125/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input208_A la_iena_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__264__A _264_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_124_ _124_/A vssd vssd vccd vccd _124_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3198 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_055_ _055_/A vssd vssd vccd vccd _055_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1730 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__430__C _430_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2160 wire2161/X vssd vssd vccd vccd wire2160/X sky130_fd_sc_hd__buf_6
Xwire2171 wire2172/X vssd vssd vccd vccd _448_/B sky130_fd_sc_hd__buf_6
XFILLER_1_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2182 wire2183/X vssd vssd vccd vccd _443_/B sky130_fd_sc_hd__buf_6
Xwire2193 wire2193/A vssd vssd vccd vccd _436_/B sky130_fd_sc_hd__buf_6
XANTENNA_wire1058_A _477_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1470 wire1471/X vssd vssd vccd vccd wire1470/X sky130_fd_sc_hd__buf_6
XFILLER_53_209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1481 wire1481/A vssd vssd vccd vccd wire1481/X sky130_fd_sc_hd__buf_6
Xwire1492 wire1493/X vssd vssd vccd vccd wire1492/X sky130_fd_sc_hd__buf_6
XFILLER_34_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1225_A _347_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output796_A _551_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__174__A _174_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[21\] mprj_dat_i_user[21] max_length1310/X vssd vssd vccd vccd
+ _135_/A sky130_fd_sc_hd__nand2_4
XFILLER_30_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput30 la_data_out_mprj[123] vssd vssd vccd vccd _492_/C sky130_fd_sc_hd__buf_4
XFILLER_50_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput41 la_data_out_mprj[18] vssd vssd vccd vccd _387_/C sky130_fd_sc_hd__clkbuf_4
Xinput52 la_data_out_mprj[28] vssd vssd vccd vccd _397_/C sky130_fd_sc_hd__clkbuf_4
Xinput63 la_data_out_mprj[38] vssd vssd vccd vccd _407_/C sky130_fd_sc_hd__clkbuf_4
Xinput74 la_data_out_mprj[48] vssd vssd vccd vccd _417_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1761_A wire1762/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput85 la_data_out_mprj[58] vssd vssd vccd vccd input85/X sky130_fd_sc_hd__buf_6
XFILLER_41_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput96 la_data_out_mprj[68] vssd vssd vccd vccd input96/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1859_A wire1860/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__621__B _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__406__A_N _406_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__349__A _349_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__531__B _531_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2075_A wire2075/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input158_A la_iena_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput401 mprj_adr_o_core[21] vssd vssd vccd vccd wire1481/A sky130_fd_sc_hd__buf_6
Xinput412 mprj_adr_o_core[31] vssd vssd vccd vccd wire1431/A sky130_fd_sc_hd__buf_6
XFILLER_22_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput423 mprj_dat_o_core[11] vssd vssd vccd vccd wire1388/A sky130_fd_sc_hd__buf_6
XFILLER_40_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput434 mprj_dat_o_core[21] vssd vssd vccd vccd wire1370/A sky130_fd_sc_hd__buf_6
XFILLER_40_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput445 mprj_dat_o_core[31] vssd vssd vccd vccd wire1358/A sky130_fd_sc_hd__buf_6
XFILLER_2_4387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput456 mprj_sel_o_core[2] vssd vssd vccd vccd _303_/B sky130_fd_sc_hd__buf_4
XANTENNA_input325_A la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__259__A _259_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input19_A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__425__C _425_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_107_ _107_/A vssd vssd vccd vccd _107_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput908 _119_/Y vssd vssd vccd vccd mprj_dat_i_core[5] sky130_fd_sc_hd__buf_8
Xoutput919 wire1208/X vssd vssd vccd vccd mprj_dat_o_user[15] sky130_fd_sc_hd__buf_8
XFILLER_45_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__429__A_N _557_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_038_ _038_/A vssd vssd vccd vccd _038_/Y sky130_fd_sc_hd__inv_2
XANTENNA__441__B _441_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output544_A wire1082/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1175_A wire1176/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output809_A _563_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1342_A wire1343/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__169__A _169_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] _219_/X vssd vssd vccd vccd _039_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_19_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__616__B _616_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1976_A wire1976/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__351__B _351_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__079__A _079_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__526__B _526_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__542__A _542_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2192_A wire2192/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input275_A la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__261__B _261_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input442_A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput220 la_iena_mprj[64] vssd vssd vccd vccd _227_/B sky130_fd_sc_hd__buf_4
XFILLER_1_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput231 la_iena_mprj[74] vssd vssd vccd vccd _237_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput242 la_iena_mprj[84] vssd vssd vccd vccd _247_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput253 la_iena_mprj[94] vssd vssd vccd vccd _257_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput264 la_oenb_mprj[103] vssd vssd vccd vccd _472_/A_N sky130_fd_sc_hd__buf_6
Xinput275 la_oenb_mprj[113] vssd vssd vccd vccd wire1593/A sky130_fd_sc_hd__buf_6
XFILLER_2_3483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput286 la_oenb_mprj[123] vssd vssd vccd vccd wire1583/A sky130_fd_sc_hd__buf_6
Xinput297 la_oenb_mprj[18] vssd vssd vccd vccd _515_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1046 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_587_ _587_/A _587_/B vssd vssd vccd vccd _587_/X sky130_fd_sc_hd__and2_2
XFILLER_32_724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__436__B _436_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output494_A wire1132/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_779 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_982 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output661_A _031_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output759_A wire1032/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1292_A wire1293/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput705 _071_/Y vssd vssd vccd vccd la_data_in_mprj[88] sky130_fd_sc_hd__buf_8
Xoutput716 _081_/Y vssd vssd vccd vccd la_data_in_mprj[98] sky130_fd_sc_hd__buf_8
XFILLER_29_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput727 _604_/X vssd vssd vccd vccd la_oenb_core[107] sky130_fd_sc_hd__buf_8
XFILLER_29_2831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput738 _614_/X vssd vssd vccd vccd la_oenb_core[117] sky130_fd_sc_hd__buf_8
XFILLER_42_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput749 _624_/X vssd vssd vccd vccd la_oenb_core[127] sky130_fd_sc_hd__buf_8
XANTENNA_output926_A wire1186/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_2897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2430 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1724_A wire1725/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_890 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__346__B _346_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[93\]_B wire1321/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__362__A _362_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_510_ _510_/A _510_/B vssd vssd vccd vccd _510_/X sky130_fd_sc_hd__and2_4
XFILLER_22_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 wire1956/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_314 wire2109/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_325 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_336 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__537__A _537_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_347 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_441_ _569_/A _441_/B _441_/C vssd vssd vccd vccd _441_/X sky130_fd_sc_hd__and3b_4
XTAP_2657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_358 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__256__B _256_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_372_ _500_/A _372_/B _372_/C vssd vssd vccd vccd _372_/X sky130_fd_sc_hd__and3b_4
XTAP_1967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2205_A wire2206/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input392_A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_B wire1330/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input86_A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__272__A _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output507_A wire1120/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1040_A _509_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1138_A _376_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1305_A _299_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output876_A wire1278/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] _182_/X vssd vssd vccd vccd _002_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_32_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[75\]_B _238_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__182__A _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1674_A wire1675/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput502 wire1144/X vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__buf_8
XFILLER_44_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput513 wire1143/X vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__buf_8
XFILLER_48_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput524 wire1142/X vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__buf_8
Xoutput535 wire1141/X vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__buf_8
Xoutput546 wire1140/X vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__buf_8
XFILLER_44_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput557 wire1139/X vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__buf_8
XANTENNA_wire1841_A wire1841/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput568 wire1138/X vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__buf_8
XFILLER_25_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1939_A wire1940/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput579 wire1137/X vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__buf_8
XFILLER_5_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__357__A _357_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1964 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1352 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__092__A _092_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1800 wire1800/A vssd vssd vccd vccd _256_/A sky130_fd_sc_hd__buf_6
XANTENNA_input140_A la_iena_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1811 wire1811/A vssd vssd vccd vccd _298_/A sky130_fd_sc_hd__buf_6
XANTENNA_wire2155_A wire2155/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1822 wire1822/A vssd vssd vccd vccd _204_/A sky130_fd_sc_hd__buf_6
XANTENNA_input238_A la_iena_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1833 wire1834/X vssd vssd vccd vccd _188_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1844 wire1844/A vssd vssd vccd vccd _181_/A sky130_fd_sc_hd__buf_6
XFILLER_46_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1855 wire1855/A vssd vssd vccd vccd wire1855/X sky130_fd_sc_hd__buf_6
XFILLER_18_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1866 wire1866/A vssd vssd vccd vccd wire1866/X sky130_fd_sc_hd__buf_6
XTAP_3122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1877 wire1878/X vssd vssd vccd vccd wire1877/X sky130_fd_sc_hd__buf_6
XTAP_3133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1888 wire1888/A vssd vssd vccd vccd wire1888/X sky130_fd_sc_hd__buf_6
XFILLER_41_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1899 wire1900/X vssd vssd vccd vccd wire1899/X sky130_fd_sc_hd__buf_6
XTAP_3155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input405_A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__267__A _267_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _547_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1706 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_155 _219_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_424_ _552_/A _424_/B _424_/C vssd vssd vccd vccd _424_/X sky130_fd_sc_hd__and3b_1
XTAP_1742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _380_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_355_ _355_/A _355_/B vssd vssd vccd vccd _355_/X sky130_fd_sc_hd__and2_1
XFILLER_50_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_286_ _286_/A _286_/B vssd vssd vccd vccd _286_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__433__C _433_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1255_A _327_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2674 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput6 la_data_out_mprj[101] vssd vssd vccd vccd _470_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1422_A wire1423/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__177__A _177_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1791_A wire1792/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1889_A wire1890/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__624__B _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] _625_/X vssd vssd vccd vccd _147_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_40_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1107 _406_/X vssd vssd vccd vccd wire1107/X sky130_fd_sc_hd__buf_6
XFILLER_29_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1118 _395_/X vssd vssd vccd vccd wire1118/X sky130_fd_sc_hd__buf_6
Xwire1129 _384_/X vssd vssd vccd vccd wire1129/X sky130_fd_sc_hd__buf_6
XFILLER_25_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__087__A _087_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4438 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[39\]_B _202_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_140_ _140_/A vssd vssd vccd vccd _140_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[123\]_B wire1313/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_071_ _071_/A vssd vssd vccd vccd _071_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input188_A la_iena_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__550__A _550_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input355_A la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__462__A_N _590_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input49_A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1630 wire1630/A vssd vssd vccd vccd _443_/C sky130_fd_sc_hd__buf_6
Xwire1641 wire1642/X vssd vssd vccd vccd _391_/B sky130_fd_sc_hd__buf_6
XFILLER_47_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1652 wire1653/X vssd vssd vccd vccd _385_/B sky130_fd_sc_hd__buf_6
XFILLER_46_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1663 wire1664/X vssd vssd vccd vccd _380_/B sky130_fd_sc_hd__buf_6
Xwire1674 wire1675/X vssd vssd vccd vccd _375_/B sky130_fd_sc_hd__buf_6
XFILLER_19_4040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1685 wire1685/A vssd vssd vccd vccd wire1685/X sky130_fd_sc_hd__buf_6
XFILLER_47_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1696 wire1697/X vssd vssd vccd vccd _365_/A sky130_fd_sc_hd__buf_6
XFILLER_38_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__428__C _428_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ _535_/A _407_/B _407_/C vssd vssd vccd vccd _407_/X sky130_fd_sc_hd__and3b_4
XTAP_1572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__444__B _444_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_B wire1314/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_338_ _338_/A _338_/B vssd vssd vccd vccd _338_/X sky130_fd_sc_hd__and2_4
XANTENNA_output574_A _454_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_269_ _269_/A _269_/B vssd vssd vccd vccd _269_/X sky130_fd_sc_hd__and2_4
Xwire971 wire971/A vssd vssd vccd vccd _069_/A sky130_fd_sc_hd__buf_6
XFILLER_31_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire982 wire982/A vssd vssd vccd vccd _105_/A sky130_fd_sc_hd__buf_6
Xwire993 wire993/A vssd vssd vccd vccd _083_/A sky130_fd_sc_hd__buf_6
XANTENNA_output741_A wire1041/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output839_A _590_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1372_A wire1373/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] wire1328/X vssd vssd vccd vccd wire971/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_39_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1637_A wire1638/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__619__B _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[23\]_A mprj_dat_i_user[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_11 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_22 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_B _268_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__354__B _354_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_33 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_44 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_55 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_66 mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_77 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_88 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_99 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__485__A_N _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2382 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_A mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2020_A wire2020/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input103_A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2118_A wire2118/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__545__A _545_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__264__B _264_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_123_ _123_/A vssd vssd vccd vccd _123_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_2421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_054_ _054_/A vssd vssd vccd vccd _054_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__280__A _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2150 wire2151/X vssd vssd vccd vccd wire2150/X sky130_fd_sc_hd__buf_6
XFILLER_1_4068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2161 wire2161/A vssd vssd vccd vccd wire2161/X sky130_fd_sc_hd__buf_6
XFILLER_40_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2172 wire2172/A vssd vssd vccd vccd wire2172/X sky130_fd_sc_hd__buf_6
XFILLER_8_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2183 wire2183/A vssd vssd vccd vccd wire2183/X sky130_fd_sc_hd__buf_6
XFILLER_5_2780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2194 wire2194/A vssd vssd vccd vccd _435_/B sky130_fd_sc_hd__buf_6
XFILLER_47_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1460 wire1461/X vssd vssd vccd vccd wire1460/X sky130_fd_sc_hd__buf_6
XFILLER_1_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1471 wire1471/A vssd vssd vccd vccd wire1471/X sky130_fd_sc_hd__buf_6
XANTENNA__439__B _439_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1482 wire1483/X vssd vssd vccd vccd _325_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1493 wire1493/A vssd vssd vccd vccd wire1493/X sky130_fd_sc_hd__buf_6
XFILLER_47_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1120_A _393_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1218_A wire1219/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output691_A _058_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output789_A _545_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[14\] mprj_dat_i_user[14] _294_/X vssd vssd vccd vccd _128_/A sky130_fd_sc_hd__nand2_2
Xinput20 la_data_out_mprj[114] vssd vssd vccd vccd _483_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput31 la_data_out_mprj[124] vssd vssd vccd vccd input31/X sky130_fd_sc_hd__buf_6
XFILLER_50_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput42 la_data_out_mprj[19] vssd vssd vccd vccd _388_/C sky130_fd_sc_hd__clkbuf_4
Xinput53 la_data_out_mprj[29] vssd vssd vccd vccd _398_/C sky130_fd_sc_hd__clkbuf_4
Xinput64 la_data_out_mprj[39] vssd vssd vccd vccd _408_/C sky130_fd_sc_hd__clkbuf_4
Xinput75 la_data_out_mprj[49] vssd vssd vccd vccd _418_/C sky130_fd_sc_hd__clkbuf_4
Xinput86 la_data_out_mprj[59] vssd vssd vccd vccd _428_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__190__A _190_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput97 la_data_out_mprj[69] vssd vssd vccd vccd input97/X sky130_fd_sc_hd__buf_6
XFILLER_6_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1921_A wire1921/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] _275_/X vssd vssd vccd vccd wire987/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA__349__B _349_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__365__A _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput402 mprj_adr_o_core[22] vssd vssd vccd vccd wire1476/A sky130_fd_sc_hd__buf_6
XFILLER_7_1629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput413 mprj_adr_o_core[3] vssd vssd vccd vccd wire1426/A sky130_fd_sc_hd__buf_6
XFILLER_9_2190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput424 mprj_dat_o_core[12] vssd vssd vccd vccd wire1386/A sky130_fd_sc_hd__buf_6
XFILLER_6_3790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2068_A wire2068/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput435 mprj_dat_o_core[22] vssd vssd vccd vccd wire1369/A sky130_fd_sc_hd__buf_6
XFILLER_0_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput446 mprj_dat_o_core[3] vssd vssd vccd vccd wire1357/A sky130_fd_sc_hd__buf_6
XFILLER_2_3643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput457 mprj_sel_o_core[3] vssd vssd vccd vccd _304_/B sky130_fd_sc_hd__buf_4
XFILLER_22_3582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input220_A la_iena_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input318_A la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__275__A _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2554 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_106_ _106_/A vssd vssd vccd vccd _106_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput909 _120_/Y vssd vssd vccd vccd mprj_dat_i_core[6] sky130_fd_sc_hd__buf_8
X_037_ _037_/A vssd vssd vccd vccd _037_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__441__C _441_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4036 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output537_A wire1092/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1070_A _465_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1168_A wire1169/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1290 wire1291/X vssd vssd vccd vccd wire1290/X sky130_fd_sc_hd__buf_8
XFILLER_39_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] _212_/X vssd vssd vccd vccd _032_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_34_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1502_A wire1503/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__185__A _185_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1871_A wire1871/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1969_A wire1970/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__095__A _095_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__542__B _542_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input170_A la_iena_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input268_A la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input435_A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput210 la_iena_mprj[55] vssd vssd vccd vccd _218_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_4_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input31_A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput221 la_iena_mprj[65] vssd vssd vccd vccd _228_/B sky130_fd_sc_hd__buf_4
XFILLER_23_1207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput232 la_iena_mprj[75] vssd vssd vccd vccd _238_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput243 la_iena_mprj[85] vssd vssd vccd vccd _248_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput254 la_iena_mprj[95] vssd vssd vccd vccd _258_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput265 la_oenb_mprj[104] vssd vssd vccd vccd wire1603/A sky130_fd_sc_hd__buf_6
XFILLER_48_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput276 la_oenb_mprj[114] vssd vssd vccd vccd wire1592/A sky130_fd_sc_hd__buf_6
Xinput287 la_oenb_mprj[124] vssd vssd vccd vccd wire1582/A sky130_fd_sc_hd__buf_6
XFILLER_18_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput298 la_oenb_mprj[19] vssd vssd vccd vccd _516_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_586_ _586_/A _586_/B vssd vssd vccd vccd _586_/X sky130_fd_sc_hd__and2_2
XFILLER_16_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__436__C _436_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output487_A _490_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__452__B _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output654_A _024_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput706 _072_/Y vssd vssd vccd vccd la_data_in_mprj[89] sky130_fd_sc_hd__buf_8
Xoutput717 _082_/Y vssd vssd vccd vccd la_data_in_mprj[99] sky130_fd_sc_hd__buf_8
XFILLER_29_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput728 _605_/X vssd vssd vccd vccd la_oenb_core[108] sky130_fd_sc_hd__buf_8
XANTENNA_wire1285_A wire1286/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput739 _615_/X vssd vssd vccd vccd la_oenb_core[118] sky130_fd_sc_hd__buf_8
XFILLER_42_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output821_A _574_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output919_A wire1208/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3290 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1452_A wire1453/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3824 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1458 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__362__B _362_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[6\]_A mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_304 _582_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_315 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 wire2078/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_337 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_440_ _568_/A _440_/B _440_/C vssd vssd vccd vccd _440_/X sky130_fd_sc_hd__and3b_4
XTAP_1913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_348 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_359 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__419__A_N _547_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_371_ _499_/A _371_/B _371_/C vssd vssd vccd vccd _371_/X sky130_fd_sc_hd__and3b_4
XFILLER_18_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2100_A wire2101/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__553__A _553_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input385_A la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__272__B _272_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input79_A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__447__B _447_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1033_A _516_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_569_ _569_/A _569_/B vssd vssd vccd vccd _569_/X sky130_fd_sc_hd__and2_4
XFILLER_31_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1200_A wire1201/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output771_A _528_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output869_A _334_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput503 wire1124/X vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__buf_8
XFILLER_9_3424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput514 wire1114/X vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__buf_8
XFILLER_44_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1667_A wire1667/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput525 wire1104/X vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__buf_8
XFILLER_48_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput536 wire1093/X vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__buf_8
XFILLER_29_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput547 wire1080/X vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__buf_8
XFILLER_42_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2662 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput558 _439_/X vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__buf_8
Xoutput569 _449_/X vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__buf_8
XFILLER_47_1549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1834_A wire1834/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__357__B _357_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3783 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1801 wire1801/A vssd vssd vccd vccd _255_/A sky130_fd_sc_hd__buf_4
XFILLER_1_3708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1812 wire1812/A vssd vssd vccd vccd _334_/A sky130_fd_sc_hd__buf_6
Xwire1823 wire1823/A vssd vssd vccd vccd _331_/A sky130_fd_sc_hd__buf_6
Xwire1834 wire1834/A vssd vssd vccd vccd wire1834/X sky130_fd_sc_hd__buf_6
Xwire1845 wire1845/A vssd vssd vccd vccd _180_/A sky130_fd_sc_hd__buf_6
XFILLER_19_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input133_A la_iena_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2050_A wire2050/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1856 wire1856/A vssd vssd vccd vccd _173_/A sky130_fd_sc_hd__buf_6
XTAP_3101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1867 wire1868/X vssd vssd vccd vccd _165_/A sky130_fd_sc_hd__buf_6
XFILLER_45_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1878 wire1878/A vssd vssd vccd vccd wire1878/X sky130_fd_sc_hd__buf_6
XANTENNA__548__A _548_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1889 wire1890/X vssd vssd vccd vccd _619_/B sky130_fd_sc_hd__buf_6
XTAP_3145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1070 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_112 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input300_A la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__267__B _267_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_123 mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _547_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _219_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1718 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_423_ _551_/A _423_/B _423_/C vssd vssd vccd vccd _423_/X sky130_fd_sc_hd__and3b_4
XANTENNA_167 _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_178 _400_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__391__A_N _519_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_354_ _354_/A _354_/B vssd vssd vccd vccd _354_/X sky130_fd_sc_hd__and2_4
XTAP_1798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__283__A _283_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_285_ _285_/A _285_/B vssd vssd vccd vccd _285_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1246 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1150_A wire1151/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput7 la_data_out_mprj[102] vssd vssd vccd vccd _471_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2686 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__177__B _177_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1415_A wire1416/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] _194_/X vssd vssd vccd vccd _014_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_138 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__193__A _193_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1784_A wire1784/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1951_A wire1952/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2542 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1108 _405_/X vssd vssd vccd vccd wire1108/X sky130_fd_sc_hd__buf_6
XFILLER_5_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1119 _394_/X vssd vssd vccd vccd wire1119/X sky130_fd_sc_hd__buf_6
XFILLER_0_4453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__368__A _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_070_ _070_/A vssd vssd vccd vccd _070_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2098_A wire2098/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__550__B _550_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input250_A la_iena_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input348_A la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1620 wire1620/A vssd vssd vccd vccd _453_/C sky130_fd_sc_hd__buf_6
XFILLER_5_2962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1631 wire1631/A vssd vssd vccd vccd _442_/C sky130_fd_sc_hd__buf_6
XFILLER_19_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1642 wire1642/A vssd vssd vccd vccd wire1642/X sky130_fd_sc_hd__buf_6
Xwire1653 wire1653/A vssd vssd vccd vccd wire1653/X sky130_fd_sc_hd__buf_6
XFILLER_47_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__278__A _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1664 wire1665/X vssd vssd vccd vccd wire1664/X sky130_fd_sc_hd__buf_6
XFILLER_24_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1675 wire1675/A vssd vssd vccd vccd wire1675/X sky130_fd_sc_hd__buf_6
XFILLER_46_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1686 wire1687/X vssd vssd vccd vccd _370_/B sky130_fd_sc_hd__buf_6
Xwire1697 wire1697/A vssd vssd vccd vccd wire1697/X sky130_fd_sc_hd__buf_6
XFILLER_47_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_406_ _406_/A_N _406_/B _406_/C vssd vssd vccd vccd _406_/X sky130_fd_sc_hd__and3b_4
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_337_ _337_/A _337_/B vssd vssd vccd vccd _337_/X sky130_fd_sc_hd__and2_4
XANTENNA__444__C _444_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_268_ _268_/A _268_/B vssd vssd vccd vccd _268_/X sky130_fd_sc_hd__and2_4
XANTENNA_output567_A _448_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire961 wire961/A vssd vssd vccd vccd _082_/A sky130_fd_sc_hd__buf_6
XFILLER_28_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire972 wire972/A vssd vssd vccd vccd _068_/A sky130_fd_sc_hd__buf_6
XFILLER_45_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire983 wire983/A vssd vssd vccd vccd _100_/A sky130_fd_sc_hd__buf_6
XFILLER_31_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire994 _587_/X vssd vssd vccd vccd wire994/X sky130_fd_sc_hd__buf_6
X_199_ _199_/A _199_/B vssd vssd vccd vccd _199_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1198_A wire1199/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__460__B _460_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output734_A _610_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1365_A wire1365/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output901_A _142_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] wire1333/X vssd vssd vccd vccd wire977/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_39_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1532_A wire1532/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__188__A _188_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[23\]_B max_length1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1999_A wire2000/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire985_A wire985/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_12 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_23 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_34 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_45 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_56 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_67 mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_78 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_89 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__370__B _370_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__098__A _098_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[14\]_B _294_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__545__B _545_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input298_A la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_122_ _122_/A vssd vssd vccd vccd _122_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_11_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__561__A _561_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_053_ _053_/A vssd vssd vccd vccd _053_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_4343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__280__B _280_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input61_A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2140 wire2140/A vssd vssd vccd vccd _464_/B sky130_fd_sc_hd__buf_6
Xwire2151 wire2151/A vssd vssd vccd vccd wire2151/X sky130_fd_sc_hd__buf_6
XFILLER_43_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2162 wire2163/X vssd vssd vccd vccd _452_/B sky130_fd_sc_hd__buf_6
Xwire2173 wire2174/X vssd vssd vccd vccd _447_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2184 wire2185/X vssd vssd vccd vccd _442_/B sky130_fd_sc_hd__buf_6
Xwire1450 wire1451/X vssd vssd vccd vccd wire1450/X sky130_fd_sc_hd__buf_6
XFILLER_5_2792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2195 wire2195/A vssd vssd vccd vccd _308_/A sky130_fd_sc_hd__buf_6
Xwire1461 wire1461/A vssd vssd vccd vccd wire1461/X sky130_fd_sc_hd__buf_6
XFILLER_47_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1472 wire1473/X vssd vssd vccd vccd _328_/B sky130_fd_sc_hd__buf_6
XANTENNA__439__C _439_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1483 wire1484/X vssd vssd vccd vccd wire1483/X sky130_fd_sc_hd__buf_6
XFILLER_1_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1494 wire1495/X vssd vssd vccd vccd _323_/B sky130_fd_sc_hd__buf_6
XFILLER_19_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__455__B _455_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output684_A _052_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput10 la_data_out_mprj[105] vssd vssd vccd vccd _474_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_output851_A wire1266/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput21 la_data_out_mprj[115] vssd vssd vccd vccd _484_/C sky130_fd_sc_hd__buf_4
XFILLER_28_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput32 la_data_out_mprj[125] vssd vssd vccd vccd input32/X sky130_fd_sc_hd__buf_6
XFILLER_11_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output949_A wire1303/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput43 la_data_out_mprj[1] vssd vssd vccd vccd _370_/C sky130_fd_sc_hd__clkbuf_4
Xinput54 la_data_out_mprj[2] vssd vssd vccd vccd _371_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput65 la_data_out_mprj[3] vssd vssd vccd vccd _372_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1482_A wire1483/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput76 la_data_out_mprj[4] vssd vssd vccd vccd _373_/C sky130_fd_sc_hd__clkbuf_4
Xinput87 la_data_out_mprj[5] vssd vssd vccd vccd _374_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__190__B _190_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput98 la_data_out_mprj[6] vssd vssd vccd vccd _375_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1747_A wire1748/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] _268_/X vssd vssd vccd vccd _088_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_0_2144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj2_logic_high_inst wire2209/A vccd2_uq0 vssd2_uq0 mprj2_logic_high
XFILLER_11_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__365__B _365_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__452__A_N _580_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput403 mprj_adr_o_core[23] vssd vssd vccd vccd wire1474/A sky130_fd_sc_hd__buf_6
XFILLER_44_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput414 mprj_adr_o_core[4] vssd vssd vccd vccd wire1421/A sky130_fd_sc_hd__buf_6
XFILLER_22_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput425 mprj_dat_o_core[13] vssd vssd vccd vccd wire1384/A sky130_fd_sc_hd__buf_6
XFILLER_22_3550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput436 mprj_dat_o_core[23] vssd vssd vccd vccd wire1368/A sky130_fd_sc_hd__buf_6
XFILLER_40_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput447 mprj_dat_o_core[4] vssd vssd vccd vccd wire1355/A sky130_fd_sc_hd__buf_6
Xinput458 mprj_stb_o_core vssd vssd vccd vccd wire1343/A sky130_fd_sc_hd__buf_6
XFILLER_25_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2130_A wire2131/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input213_A la_iena_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_959 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__556__A _556_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__275__B _275_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__291__A _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_105_ _105_/A vssd vssd vccd vccd _105_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_036_ _036_/A vssd vssd vccd vccd _036_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4048 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1063_A _472_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1280 wire1281/X vssd vssd vccd vccd wire1280/X sky130_fd_sc_hd__buf_8
Xwire1291 wire1292/X vssd vssd vccd vccd wire1291/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1230_A wire1231/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__475__A_N _603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1328_A _249_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__185__B _185_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1697_A wire1697/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1864_A wire1864/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1906 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high_inst wire2204/A _395_/B _396_/B _397_/B _398_/B _399_/B _400_/B _401_/B
+ _402_/B _403_/B _404_/B wire2202/A _405_/B _406_/B _407_/B _408_/B _409_/B _410_/B
+ _411_/B _412_/B _413_/B _414_/B wire2200/A _415_/B _416_/B _417_/B _418_/B _419_/B
+ _420_/B _421_/B _422_/B _423_/B _424_/B wire2199/A _425_/B _426_/B _427_/B _428_/B
+ _429_/B _430_/B _431_/B wire2198/A wire2197/A wire2196/A wire2195/A wire2194/A wire2193/A
+ wire2192/A wire2191/A wire2190/A wire2188/A wire2187/A wire2185/A wire2183/A wire2181/A
+ wire2179/A wire2178/A wire2176/A wire2174/A wire2172/A wire2170/A wire2168/A wire2166/A
+ wire2164/A wire2161/A wire2158/A wire2155/A wire2154/A wire2151/A wire2148/A wire2145/A
+ wire2144/A wire2143/A wire2142/A _462_/B wire2141/A wire2140/A _311_/A wire2139/A
+ wire2138/A wire2136/A wire2135/A wire2134/A wire2132/A wire2131/A wire2129/A wire2127/A
+ wire2125/A _312_/A wire2123/A wire2122/A wire2120/A wire2118/A wire2116/A wire2114/A
+ wire2111/A wire2109/A wire2107/A wire2104/A _313_/A wire2101/A wire2098/A wire2096/A
+ wire2093/A wire2090/A wire2087/A wire2084/A wire2081/A wire2078/A wire2075/A _314_/A
+ _296_/A wire2072/A wire2068/A wire2065/A wire2063/A wire2061/A wire2059/A wire2057/A
+ wire2056/A wire2054/A wire2052/A _315_/A wire2051/A wire2050/A wire2048/A wire2046/A
+ wire2044/A wire2043/A wire2041/A wire2039/A wire2038/A wire2036/A _316_/A wire2035/A
+ wire2034/A wire2033/A wire2032/A wire2031/A wire2030/A wire2029/A _522_/B wire2028/A
+ _524_/B _317_/A wire2027/A _526_/B _527_/B _528_/B _529_/B _530_/B wire2026/A _532_/B
+ _533_/B _534_/B _318_/A wire2025/A _536_/B _537_/B _538_/B wire2024/A _540_/B _541_/B
+ _542_/B _543_/B _544_/B _319_/A _545_/B wire2023/A _547_/B _548_/B _549_/B _550_/B
+ _551_/B _552_/B _553_/B _554_/B _320_/A _555_/B _556_/B _557_/B _558_/B wire2022/A
+ wire2021/A wire2020/A wire2019/A wire2018/A wire2017/A _321_/A wire2016/A wire2015/A
+ wire2014/A wire2013/A wire2011/A wire2009/A wire2008/A wire2006/A wire2004/A wire2002/A
+ _322_/A wire2000/A wire1997/A wire1995/A wire1993/A wire1991/A wire1989/A wire1987/A
+ wire1985/A wire1983/A wire1980/A _323_/A wire1978/A wire1976/A wire1975/A wire1974/A
+ wire1972/A wire1971/A wire1970/A wire1968/A wire1966/A wire1964/A _324_/A wire1962/A
+ wire1958/A wire1956/A wire1954/A wire1952/A wire1949/A wire1947/A wire1944/A wire1942/A
+ wire1940/A wire1938/A _325_/A wire1936/A wire1933/A wire1930/A wire1927/A wire1924/A
+ wire1921/A wire1918/A wire1914/A wire1910/A wire1907/A _326_/A wire1904/A wire1901/A
+ wire1897/A wire1894/A wire1891/A wire1888/A wire1885/A wire1882/A wire1878/A wire1875/A
+ _327_/A wire1871/A wire1870/A wire1868/A wire1866/A wire1864/A wire1862/A wire1861/A
+ wire1860/A wire1858/A wire1857/A _328_/A wire1856/A wire1855/A wire1853/A wire1851/A
+ wire1849/A wire1848/A wire1846/A wire1845/A wire1844/A wire1843/A wire1842/A wire1841/A
+ wire1840/A wire1839/A wire1838/A wire1836/A wire1834/A wire1832/A wire1830/A wire1829/A
+ wire1828/A wire1827/A wire1826/A wire1825/A wire1824/A _196_/A _197_/A _198_/A _199_/A
+ _200_/A _201_/A _202_/A wire1823/A _203_/A wire1822/A wire1821/A wire1820/A wire1819/A
+ wire1818/A _209_/A _210_/A _211_/A _212_/A wire1817/A _213_/A _214_/A _215_/A _216_/A
+ _217_/A _218_/A _219_/A _220_/A _221_/A _222_/A wire1816/A _223_/A _224_/A _225_/A
+ _226_/A _227_/A _228_/A _229_/A wire1815/A wire1814/A wire1813/A wire1812/A wire1811/A
+ wire1810/A _234_/A _235_/A _236_/A _237_/A _238_/A _239_/A _240_/A _241_/A _242_/A
+ wire1809/A _243_/A wire1808/A wire1807/A _246_/A _247_/A _248_/A wire1806/A wire1805/A
+ wire1804/A _252_/A wire1803/A _253_/A wire1802/A wire1801/A wire1800/A wire1799/A
+ wire1798/A wire1797/A wire1796/A wire1794/A wire1792/A _337_/A wire1790/A wire1788/A
+ wire1786/A wire1784/A wire1783/A wire1781/A wire1779/A wire1777/A wire1776/A wire1774/A
+ _338_/A wire1772/A wire1770/A wire1768/A wire1766/A wire1764/A wire1762/A wire1760/A
+ wire1758/A wire1756/A wire1754/A _339_/A wire1752/A wire1750/A wire1748/A wire1745/A
+ wire1743/A wire1741/A wire1739/A wire1737/A wire1734/A wire1731/A _340_/A wire1728/A
+ wire1725/A wire1722/A _341_/A _342_/A _343_/A _344_/A _299_/A _345_/A _346_/A _347_/A
+ _348_/A _349_/A wire1719/A wire1718/A wire1717/A wire1716/A wire1715/A wire1714/A
+ wire1713/A wire1712/A wire1711/A wire1710/A wire1709/A wire1708/A wire1707/A wire1705/A
+ wire1703/A wire1701/A wire1699/A wire1697/A wire1695/A wire1693/A wire1691/A wire1689/A
+ wire1687/A wire1685/A wire1683/A wire1681/A wire1679/A wire1677/A wire1675/A wire1673/A
+ wire1671/A wire1669/A wire1667/A wire1665/A wire1662/A wire1660/A wire1658/A wire1656/A
+ wire1654/A wire1653/A wire1651/A wire1649/A wire1647/A wire1645/A wire1644/A wire1642/A
+ wire1640/A wire1638/A wire1636/A wire1634/A vccd1_uq1 vssd1_uq1 mprj_logic_high
XTAP_3508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2080_A wire2081/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input163_A la_iena_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2178_A wire2178/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput200 la_iena_mprj[46] vssd vssd vccd vccd _209_/B sky130_fd_sc_hd__buf_4
Xinput211 la_iena_mprj[56] vssd vssd vccd vccd _219_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput222 la_iena_mprj[66] vssd vssd vccd vccd _229_/B sky130_fd_sc_hd__buf_4
XFILLER_0_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput233 la_iena_mprj[76] vssd vssd vccd vccd _239_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_input330_A la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput244 la_iena_mprj[86] vssd vssd vccd vccd _249_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_input428_A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput255 la_iena_mprj[96] vssd vssd vccd vccd _259_/B sky130_fd_sc_hd__clkbuf_4
Xinput266 la_oenb_mprj[105] vssd vssd vccd vccd wire1602/A sky130_fd_sc_hd__buf_6
XFILLER_40_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input24_A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput277 la_oenb_mprj[115] vssd vssd vccd vccd wire1591/A sky130_fd_sc_hd__buf_6
XFILLER_40_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput288 la_oenb_mprj[125] vssd vssd vccd vccd wire1581/A sky130_fd_sc_hd__buf_6
Xinput299 la_oenb_mprj[1] vssd vssd vccd vccd _498_/A sky130_fd_sc_hd__buf_4
XFILLER_18_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__286__A _286_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_585_ _585_/A _585_/B vssd vssd vccd vccd _585_/X sky130_fd_sc_hd__and2_4
XFILLER_17_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__452__C _452_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput707 _155_/Y vssd vssd vccd vccd la_data_in_mprj[8] sky130_fd_sc_hd__buf_8
Xoutput718 _156_/Y vssd vssd vccd vccd la_data_in_mprj[9] sky130_fd_sc_hd__buf_8
XFILLER_10_2082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput729 _606_/X vssd vssd vccd vccd la_oenb_core[109] sky130_fd_sc_hd__buf_8
XANTENNA_output647_A _018_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_019_ _019_/A vssd vssd vccd vccd _019_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1180_A wire1181/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1278_A wire1279/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output814_A _567_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1445_A wire1446/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] _224_/X vssd vssd vccd vccd _044_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_23_2498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__196__A _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1981_A wire1982/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[6\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_305 _579_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_316 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_327 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_349 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ _498_/A _370_/B _370_/C vssd vssd vccd vccd _370_/X sky130_fd_sc_hd__and3b_4
XTAP_1947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__553__B _553_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input280_A la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input378_A la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_542 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__447__C _447_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_568_ _568_/A _568_/B vssd vssd vccd vccd _568_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1026_A _523_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output597_A _088_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2578 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_499_ _499_/A _499_/B vssd vssd vccd vccd _499_/X sky130_fd_sc_hd__and2_4
XFILLER_31_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__463__B _463_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output764_A wire1027/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1395_A wire1396/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput504 wire1123/X vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__buf_8
XANTENNA_output931_A wire1166/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput515 wire1113/X vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__buf_8
XFILLER_44_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput526 wire1103/X vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__buf_8
Xoutput537 wire1092/X vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__buf_8
Xoutput548 wire1079/X vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__buf_8
XFILLER_47_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput559 _440_/X vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__buf_8
XFILLER_25_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2674 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1827_A wire1827/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__373__B _373_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1802 wire1802/A vssd vssd vccd vccd _254_/A sky130_fd_sc_hd__buf_6
XFILLER_5_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1813 wire1813/A vssd vssd vccd vccd _232_/A sky130_fd_sc_hd__buf_6
Xwire1824 wire1824/A vssd vssd vccd vccd _195_/A sky130_fd_sc_hd__buf_4
XFILLER_41_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1835 wire1836/X vssd vssd vccd vccd _187_/A sky130_fd_sc_hd__buf_6
Xwire1846 wire1846/A vssd vssd vccd vccd _179_/A sky130_fd_sc_hd__buf_6
XTAP_3102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1857 wire1857/A vssd vssd vccd vccd _172_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1868 wire1868/A vssd vssd vccd vccd wire1868/X sky130_fd_sc_hd__buf_6
XFILLER_41_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1879 wire1880/X vssd vssd vccd vccd _622_/B sky130_fd_sc_hd__buf_6
XFILLER_46_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__548__B _548_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2043_A wire2043/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input126_A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_113 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _431_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_135 _547_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_146 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _220_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_422_ _550_/A _422_/B _422_/C vssd vssd vccd vccd _422_/X sky130_fd_sc_hd__and3b_4
XTAP_1722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_179 _550_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__564__A _564_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XTAP_1777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_353_ _353_/A _353_/B vssd vssd vccd vccd _353_/X sky130_fd_sc_hd__and2_4
XTAP_1788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input91_A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_284_ _284_/A _284_/B vssd vssd vccd vccd _284_/X sky130_fd_sc_hd__and2_4
XFILLER_52_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[7\] mprj_dat_i_user[7] max_length1311/X vssd vssd vccd vccd _121_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_48_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1258 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output512_A wire1115/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput8 la_data_out_mprj[103] vssd vssd vccd vccd _472_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__458__B _458_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1143_A _371_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1408_A wire1408/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_36_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] _187_/X vssd vssd vccd vccd _007_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__193__B _193_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1777_A wire1777/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1944_A wire1944/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__409__A_N _409_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2554 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1109 _404_/X vssd vssd vccd vccd wire1109/X sky130_fd_sc_hd__buf_6
XFILLER_5_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__368__B _368_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1474 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_51_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3802 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput890 _132_/Y vssd vssd vccd vccd mprj_dat_i_core[18] sky130_fd_sc_hd__buf_8
XFILLER_43_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2160_A wire2161/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input243_A la_iena_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1610 wire1610/A vssd vssd vccd vccd _230_/B sky130_fd_sc_hd__buf_4
XANTENNA__559__A _559_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1621 wire1621/A vssd vssd vccd vccd _452_/C sky130_fd_sc_hd__buf_6
XFILLER_4_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1632 wire1632/A vssd vssd vccd vccd _441_/C sky130_fd_sc_hd__buf_6
Xwire1643 wire1644/X vssd vssd vccd vccd _390_/B sky130_fd_sc_hd__buf_6
XFILLER_46_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1654 wire1654/A vssd vssd vccd vccd _303_/A sky130_fd_sc_hd__buf_6
XANTENNA_input410_A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__278__B _278_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1665 wire1665/A vssd vssd vccd vccd wire1665/X sky130_fd_sc_hd__buf_6
Xwire1676 wire1677/X vssd vssd vccd vccd _302_/A sky130_fd_sc_hd__buf_6
XFILLER_46_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1687 wire1687/A vssd vssd vccd vccd wire1687/X sky130_fd_sc_hd__buf_6
XFILLER_34_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1698 wire1699/X vssd vssd vccd vccd _301_/A sky130_fd_sc_hd__buf_6
XTAP_2220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__294__A _294_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_405_ _405_/A_N _405_/B _405_/C vssd vssd vccd vccd _405_/X sky130_fd_sc_hd__and3b_4
XTAP_1552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_336_ _336_/A _336_/B vssd vssd vccd vccd _336_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_267_ _267_/A _267_/B vssd vssd vccd vccd _267_/X sky130_fd_sc_hd__and2_4
Xwire962 wire962/A vssd vssd vccd vccd _078_/A sky130_fd_sc_hd__buf_6
XFILLER_10_3883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire973 wire973/A vssd vssd vccd vccd _067_/A sky130_fd_sc_hd__buf_6
X_198_ _198_/A _198_/B vssd vssd vccd vccd _198_/X sky130_fd_sc_hd__and2_2
Xwire984 wire984/A vssd vssd vccd vccd _098_/A sky130_fd_sc_hd__buf_6
XFILLER_45_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire995 _586_/X vssd vssd vccd vccd wire995/X sky130_fd_sc_hd__buf_6
XFILLER_26_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__460__C _460_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1093_A wire1094/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output727_A _604_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1358_A wire1358/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__188__B _188_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1525_A wire1526/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1894_A wire1894/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_13 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_24 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_35 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_46 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1947 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_57 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_68 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_79 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__370__C _370_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__381__A_N _509_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2006_A wire2006/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_121_ _121_/A vssd vssd vccd vccd _121_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input193_A la_iena_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_052_ _052_/A vssd vssd vccd vccd _052_/Y sky130_fd_sc_hd__inv_2
XANTENNA__561__B _561_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input360_A la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input458_A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input54_A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2130 wire2131/X vssd vssd vccd vccd _471_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2141 wire2141/A vssd vssd vccd vccd _463_/B sky130_fd_sc_hd__buf_6
XANTENNA__289__A _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2152 wire2153/X vssd vssd vccd vccd _455_/B sky130_fd_sc_hd__buf_6
XFILLER_38_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2163 wire2164/X vssd vssd vccd vccd wire2163/X sky130_fd_sc_hd__buf_6
Xwire2174 wire2174/A vssd vssd vccd vccd wire2174/X sky130_fd_sc_hd__buf_6
XFILLER_47_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1440 wire1441/X vssd vssd vccd vccd wire1440/X sky130_fd_sc_hd__buf_6
Xwire2185 wire2185/A vssd vssd vccd vccd wire2185/X sky130_fd_sc_hd__buf_6
XFILLER_1_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1451 wire1451/A vssd vssd vccd vccd wire1451/X sky130_fd_sc_hd__buf_6
XFILLER_21_2552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2196 wire2196/A vssd vssd vccd vccd _434_/B sky130_fd_sc_hd__buf_6
XFILLER_4_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1462 wire1463/X vssd vssd vccd vccd _330_/B sky130_fd_sc_hd__buf_8
XFILLER_21_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1473 wire1474/X vssd vssd vccd vccd wire1473/X sky130_fd_sc_hd__buf_6
XFILLER_1_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1484 wire1484/A vssd vssd vccd vccd wire1484/X sky130_fd_sc_hd__buf_6
XFILLER_46_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1495 wire1496/X vssd vssd vccd vccd wire1495/X sky130_fd_sc_hd__buf_6
Xpowergood_check vccd vssd vdda1_uq0 vssa1_uq0 vdda2_uq0 vssa2_uq0 output954/A output952/A
+ mgmt_protect_hv
XFILLER_19_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__455__C _455_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1106_A _407_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_319_ _319_/A _319_/B vssd vssd vccd vccd _319_/X sky130_fd_sc_hd__and2_2
XFILLER_50_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput11 la_data_out_mprj[106] vssd vssd vccd vccd _475_/C sky130_fd_sc_hd__clkbuf_4
Xinput22 la_data_out_mprj[116] vssd vssd vccd vccd input22/X sky130_fd_sc_hd__clkbuf_4
Xinput33 la_data_out_mprj[126] vssd vssd vccd vccd input33/X sky130_fd_sc_hd__buf_6
XANTENNA__471__B _471_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput44 la_data_out_mprj[20] vssd vssd vccd vccd _389_/C sky130_fd_sc_hd__clkbuf_4
Xinput55 la_data_out_mprj[30] vssd vssd vccd vccd _399_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output844_A _595_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput66 la_data_out_mprj[40] vssd vssd vccd vccd _409_/C sky130_fd_sc_hd__clkbuf_4
Xinput77 la_data_out_mprj[50] vssd vssd vccd vccd _419_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput88 la_data_out_mprj[60] vssd vssd vccd vccd _429_/C sky130_fd_sc_hd__clkbuf_4
Xinput99 la_data_out_mprj[70] vssd vssd vccd vccd input99/X sky130_fd_sc_hd__buf_6
XFILLER_28_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1475_A wire1476/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] wire1323/X vssd vssd vccd vccd wire966/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_48_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1642_A wire1642/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__199__A _199_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1907_A wire1907/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__381__B _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput404 mprj_adr_o_core[24] vssd vssd vccd vccd wire1471/A sky130_fd_sc_hd__buf_6
XFILLER_40_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput415 mprj_adr_o_core[5] vssd vssd vccd vccd wire1416/A sky130_fd_sc_hd__buf_6
XFILLER_44_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput426 mprj_dat_o_core[14] vssd vssd vccd vccd wire1382/A sky130_fd_sc_hd__buf_6
XFILLER_6_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput437 mprj_dat_o_core[24] vssd vssd vccd vccd wire1367/A sky130_fd_sc_hd__buf_6
XFILLER_40_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput448 mprj_dat_o_core[5] vssd vssd vccd vccd wire1353/A sky130_fd_sc_hd__buf_6
Xinput459 mprj_we_o_core vssd vssd vccd vccd wire1341/A sky130_fd_sc_hd__buf_6
XFILLER_29_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_798 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2123_A wire2123/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input206_A la_iena_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__572__A _572_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_104_ _104_/A vssd vssd vccd vccd _104_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_8_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__291__B _291_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_035_ _035_/A vssd vssd vccd vccd _035_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1056_A _479_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1270 _316_/X vssd vssd vccd vccd wire1270/X sky130_fd_sc_hd__buf_6
Xwire1281 wire1282/X vssd vssd vccd vccd wire1281/X sky130_fd_sc_hd__buf_6
XFILLER_19_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1292 wire1293/X vssd vssd vccd vccd wire1292/X sky130_fd_sc_hd__buf_6
XFILLER_19_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__466__B _466_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1223_A wire1224/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output794_A wire1007/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1857_A wire1857/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__376__B _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_B wire1318/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2073_A wire2074/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input156_A la_iena_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput201 la_iena_mprj[47] vssd vssd vccd vccd _210_/B sky130_fd_sc_hd__buf_4
XFILLER_27_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput212 la_iena_mprj[57] vssd vssd vccd vccd _220_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput223 la_iena_mprj[67] vssd vssd vccd vccd wire1610/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput234 la_iena_mprj[77] vssd vssd vccd vccd _240_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 la_iena_mprj[87] vssd vssd vccd vccd _250_/B sky130_fd_sc_hd__clkbuf_4
Xinput256 la_iena_mprj[97] vssd vssd vccd vccd _260_/B sky130_fd_sc_hd__buf_4
XFILLER_2_3453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput267 la_oenb_mprj[106] vssd vssd vccd vccd wire1601/A sky130_fd_sc_hd__buf_6
XANTENNA_input323_A la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput278 la_oenb_mprj[116] vssd vssd vccd vccd wire1590/A sky130_fd_sc_hd__buf_6
Xinput289 la_oenb_mprj[126] vssd vssd vccd vccd wire1580/A sky130_fd_sc_hd__buf_6
XANTENNA__567__A _567_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input17_A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__286__B _286_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_584_ _584_/A _584_/B vssd vssd vccd vccd _584_/X sky130_fd_sc_hd__and2_4
XFILLER_16_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[87\]_B wire1327/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput708 _073_/Y vssd vssd vccd vccd la_data_in_mprj[90] sky130_fd_sc_hd__buf_8
XFILLER_29_2823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput719 wire1053/X vssd vssd vccd vccd la_oenb_core[0] sky130_fd_sc_hd__buf_8
X_018_ _018_/A vssd vssd vccd vccd _018_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output542_A wire1085/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1173_A _362_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[11\]_B _174_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__442__A_N _570_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output807_A _561_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1438_A wire1439/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] _217_/X vssd vssd vccd vccd _037_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_B _241_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1974_A wire1974/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input9_A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_306 _565_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_317 wire1985/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_328 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_339 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3450 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input273_A la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__465__A_N _593_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input440_A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__297__A _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1870 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_567_ _567_/A _567_/B vssd vssd vccd vccd _567_/X sky130_fd_sc_hd__and2_4
XFILLER_53_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_498_ _498_/A _498_/B vssd vssd vccd vccd _498_/X sky130_fd_sc_hd__and2_4
XANTENNA_output492_A _495_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1019_A _536_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__463__C _463_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2194 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output757_A wire1033/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1290_A wire1291/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput505 wire1122/X vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__buf_8
Xoutput516 wire1112/X vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__buf_8
Xoutput527 wire1102/X vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__buf_8
XFILLER_29_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput538 wire1091/X vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__buf_8
XANTENNA_output924_A wire1249/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput549 wire1078/X vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__buf_8
XFILLER_42_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1722_A wire1722/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__000__A _000_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_4324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__488__A_N _616_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1803 wire1803/A vssd vssd vccd vccd _336_/A sky130_fd_sc_hd__buf_6
Xwire1814 wire1814/A vssd vssd vccd vccd _231_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1825 wire1825/A vssd vssd vccd vccd _194_/A sky130_fd_sc_hd__buf_6
Xwire1836 wire1836/A vssd vssd vccd vccd wire1836/X sky130_fd_sc_hd__buf_6
XFILLER_3_3570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1847 wire1848/X vssd vssd vccd vccd _178_/A sky130_fd_sc_hd__buf_6
XTAP_3103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1858 wire1858/A vssd vssd vccd vccd _171_/A sky130_fd_sc_hd__buf_6
XTAP_3114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1869 wire1870/X vssd vssd vccd vccd _164_/A sky130_fd_sc_hd__buf_6
XFILLER_18_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2036_A wire2036/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_125 _431_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_421_ _549_/A _421_/B _421_/C vssd vssd vccd vccd _421_/X sky130_fd_sc_hd__and3b_4
XANTENNA_136 _547_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_147 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _220_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__564__B _564_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_352_ _352_/A _352_/B vssd vssd vccd vccd _352_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[126\]_B _289_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2203_A wire2204/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_283_ _283_/A _283_/B vssd vssd vccd vccd _283_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input390_A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input84_A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__580__A _580_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3470 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput9 la_data_out_mprj[104] vssd vssd vccd vccd _473_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__458__C _458_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output505_A wire1122/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1136_A _378_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_619_ _619_/A _619_/B vssd vssd vccd vccd _619_/X sky130_fd_sc_hd__and2_4
XFILLER_17_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__474__B _474_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[117\]_B _280_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1303_A wire1304/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] _180_/X vssd vssd vccd vccd _000_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_11_3829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1672_A wire1673/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1937_A wire1938/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2494 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_A mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3008 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__384__B _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_B _271_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput880 wire1306/X vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__buf_8
Xoutput891 _133_/Y vssd vssd vccd vccd mprj_dat_i_core[19] sky130_fd_sc_hd__buf_8
XFILLER_5_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1600 wire1600/A vssd vssd vccd vccd _604_/A sky130_fd_sc_hd__buf_6
Xwire1611 input22/X vssd vssd vccd vccd _485_/C sky130_fd_sc_hd__buf_4
XFILLER_21_3446 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__559__B _559_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1622 wire1622/A vssd vssd vccd vccd _451_/C sky130_fd_sc_hd__buf_6
XANTENNA_input236_A la_iena_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2153_A wire2154/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[17\]_A mprj_dat_i_user[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1633 wire1633/A vssd vssd vccd vccd _440_/C sky130_fd_sc_hd__buf_4
XFILLER_4_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1644 wire1644/A vssd vssd vccd vccd wire1644/X sky130_fd_sc_hd__buf_6
XFILLER_41_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1655 wire1656/X vssd vssd vccd vccd _384_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1666 wire1667/X vssd vssd vccd vccd _379_/B sky130_fd_sc_hd__buf_6
XFILLER_19_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1677 wire1677/A vssd vssd vccd vccd wire1677/X sky130_fd_sc_hd__buf_6
Xwire1688 wire1689/X vssd vssd vccd vccd _369_/B sky130_fd_sc_hd__buf_6
XFILLER_41_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1699 wire1699/A vssd vssd vccd vccd wire1699/X sky130_fd_sc_hd__buf_6
XANTENNA_input403_A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__575__A _575_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_170 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__294__B _294_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_404_ _532_/A _404_/B _404_/C vssd vssd vccd vccd _404_/X sky130_fd_sc_hd__and3b_4
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_335_ _335_/A _335_/B vssd vssd vccd vccd _335_/X sky130_fd_sc_hd__and2_4
XFILLER_30_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_266_ _266_/A _266_/B vssd vssd vccd vccd _266_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3840 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire963 wire963/A vssd vssd vccd vccd _077_/A sky130_fd_sc_hd__buf_6
XFILLER_26_4003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_197_ _197_/A _197_/B vssd vssd vccd vccd _197_/X sky130_fd_sc_hd__and2_2
Xwire974 wire974/A vssd vssd vccd vccd _066_/A sky130_fd_sc_hd__buf_6
Xwire985 wire985/A vssd vssd vccd vccd _097_/A sky130_fd_sc_hd__buf_6
XFILLER_48_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire996 _558_/X vssd vssd vccd vccd wire996/X sky130_fd_sc_hd__buf_6
XFILLER_26_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__469__B _469_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1253_A _328_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_936 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1420_A wire1421/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1518_A wire1519/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_14 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_25 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1887_A wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_36 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_47 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_58 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_69 mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__379__B _379_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_120_ _120_/A vssd vssd vccd vccd _120_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_051_ _051_/A vssd vssd vccd vccd _051_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input186_A la_iena_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input353_A la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input47_A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2120 wire2120/A vssd vssd vccd vccd wire2120/X sky130_fd_sc_hd__buf_6
XFILLER_1_4027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2131 wire2131/A vssd vssd vccd vccd wire2131/X sky130_fd_sc_hd__buf_6
XANTENNA__289__B _289_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2142 wire2142/A vssd vssd vccd vccd _461_/B sky130_fd_sc_hd__buf_6
XFILLER_5_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2153 wire2154/X vssd vssd vccd vccd wire2153/X sky130_fd_sc_hd__buf_6
Xwire2164 wire2164/A vssd vssd vccd vccd wire2164/X sky130_fd_sc_hd__buf_6
Xwire1430 wire1431/X vssd vssd vccd vccd wire1430/X sky130_fd_sc_hd__buf_6
Xwire2175 wire2176/X vssd vssd vccd vccd _446_/B sky130_fd_sc_hd__buf_6
Xwire1441 wire1441/A vssd vssd vccd vccd wire1441/X sky130_fd_sc_hd__buf_6
XFILLER_1_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2186 wire2187/X vssd vssd vccd vccd _441_/B sky130_fd_sc_hd__buf_6
Xwire1452 wire1453/X vssd vssd vccd vccd _332_/B sky130_fd_sc_hd__buf_8
Xwire2197 wire2197/A vssd vssd vccd vccd _433_/B sky130_fd_sc_hd__buf_6
XFILLER_46_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1463 wire1464/X vssd vssd vccd vccd wire1463/X sky130_fd_sc_hd__buf_6
Xwire1474 wire1474/A vssd vssd vccd vccd wire1474/X sky130_fd_sc_hd__buf_6
Xwire1485 wire1486/X vssd vssd vccd vccd _306_/B sky130_fd_sc_hd__buf_6
XFILLER_47_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1496 wire1497/X vssd vssd vccd vccd wire1496/X sky130_fd_sc_hd__buf_6
XFILLER_46_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_318_ _318_/A _318_/B vssd vssd vccd vccd _318_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1001_A _555_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output572_A _452_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput12 la_data_out_mprj[107] vssd vssd vccd vccd _476_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_30_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput23 la_data_out_mprj[117] vssd vssd vccd vccd _486_/C sky130_fd_sc_hd__clkbuf_4
Xinput34 la_data_out_mprj[127] vssd vssd vccd vccd input34/X sky130_fd_sc_hd__clkbuf_4
Xinput45 la_data_out_mprj[21] vssd vssd vccd vccd _390_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__471__C _471_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_249_ _249_/A _249_/B vssd vssd vccd vccd _249_/X sky130_fd_sc_hd__and2_4
XFILLER_45_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput56 la_data_out_mprj[31] vssd vssd vccd vccd _400_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_7_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput67 la_data_out_mprj[41] vssd vssd vccd vccd _410_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput78 la_data_out_mprj[51] vssd vssd vccd vccd _420_/C sky130_fd_sc_hd__clkbuf_4
Xinput89 la_data_out_mprj[61] vssd vssd vccd vccd _430_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output837_A _588_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1370_A wire1370/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1468_A wire1469/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] wire1330/X vssd vssd vccd vccd wire973/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__199__B _199_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1635_A wire1636/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3846 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__381__C _381_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput405 mprj_adr_o_core[25] vssd vssd vccd vccd wire1466/A sky130_fd_sc_hd__buf_6
XFILLER_40_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput416 mprj_adr_o_core[6] vssd vssd vccd vccd wire1411/A sky130_fd_sc_hd__buf_6
XFILLER_2_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput427 mprj_dat_o_core[15] vssd vssd vccd vccd wire1380/A sky130_fd_sc_hd__buf_6
XFILLER_44_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput438 mprj_dat_o_core[25] vssd vssd vccd vccd wire1366/A sky130_fd_sc_hd__buf_6
Xinput449 mprj_dat_o_core[6] vssd vssd vccd vccd wire1351/A sky130_fd_sc_hd__buf_6
XFILLER_2_3657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input101_A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__572__B _572_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_103_ _103_/A vssd vssd vccd vccd _103_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_034_ _034_/A vssd vssd vccd vccd _034_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_4225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1260 _321_/X vssd vssd vccd vccd wire1260/X sky130_fd_sc_hd__buf_6
XFILLER_1_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1271 wire1272/X vssd vssd vccd vccd wire1271/X sky130_fd_sc_hd__buf_6
XFILLER_40_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1282 wire1283/X vssd vssd vccd vccd wire1282/X sky130_fd_sc_hd__buf_6
XFILLER_1_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1293 _302_/X vssd vssd vccd vccd wire1293/X sky130_fd_sc_hd__buf_6
XFILLER_47_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1049_A _501_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__466__C _466_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1216_A _350_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output787_A _543_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__371__A_N _499_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__B _482_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output954_A output954/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[12\] mprj_dat_i_user[12] max_length1311/X vssd vssd vccd vccd
+ _126_/A sky130_fd_sc_hd__nand2_2
XFILLER_12_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1752_A wire1752/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] _273_/X vssd vssd vccd vccd wire989/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_27_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__392__B _392_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_A mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput202 la_iena_mprj[48] vssd vssd vccd vccd _211_/B sky130_fd_sc_hd__clkbuf_4
Xinput213 la_iena_mprj[58] vssd vssd vccd vccd _221_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput224 la_iena_mprj[68] vssd vssd vccd vccd wire1609/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input149_A la_iena_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2066_A wire2067/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput235 la_iena_mprj[78] vssd vssd vccd vccd _241_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput246 la_iena_mprj[88] vssd vssd vccd vccd _251_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput257 la_iena_mprj[98] vssd vssd vccd vccd _261_/B sky130_fd_sc_hd__buf_4
Xinput268 la_oenb_mprj[107] vssd vssd vccd vccd wire1600/A sky130_fd_sc_hd__buf_6
XFILLER_40_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput279 la_oenb_mprj[117] vssd vssd vccd vccd wire1589/A sky130_fd_sc_hd__buf_6
XFILLER_18_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__567__B _567_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input316_A la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_583_ _583_/A _583_/B vssd vssd vccd vccd _583_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__394__A_N _522_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__583__A _583_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput709 _074_/Y vssd vssd vccd vccd la_data_in_mprj[91] sky130_fd_sc_hd__buf_8
XFILLER_7_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_017_ _017_/A vssd vssd vccd vccd _017_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output535_A wire1141/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1166_A wire1167/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__477__B _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1090 _422_/X vssd vssd vccd vccd wire1090/X sky130_fd_sc_hd__buf_6
XFILLER_47_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] _210_/X vssd vssd vccd vccd _030_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1967_A wire1968/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] _172_/X vssd vssd vccd vccd _156_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_28_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__387__B _387_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_307 wire2116/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_318 wire1985/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_329 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2183_A wire2183/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input266_A la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input433_A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__578__A _578_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_566_ _566_/A _566_/B vssd vssd vccd vccd _566_/X sky130_fd_sc_hd__and2_4
XFILLER_32_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_497_ _497_/A _497_/B vssd vssd vccd vccd _497_/X sky130_fd_sc_hd__and2_4
XFILLER_32_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output485_A wire1133/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput506 wire1121/X vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__buf_8
XFILLER_9_3427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput517 wire1111/X vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__buf_8
Xoutput528 wire1101/X vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__buf_8
XANTENNA_wire1283_A _304_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput539 wire1090/X vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__buf_8
XFILLER_10_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output917_A wire1214/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1450_A wire1451/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1715_A wire1715/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1804 wire1804/A vssd vssd vccd vccd _251_/A sky130_fd_sc_hd__buf_6
Xwire1815 wire1815/A vssd vssd vccd vccd _230_/A sky130_fd_sc_hd__buf_6
XFILLER_41_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1826 wire1826/A vssd vssd vccd vccd _193_/A sky130_fd_sc_hd__buf_6
XTAP_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1837 wire1838/X vssd vssd vccd vccd _186_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1848 wire1848/A vssd vssd vccd vccd wire1848/X sky130_fd_sc_hd__buf_6
XTAP_3104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1859 wire1860/X vssd vssd vccd vccd _170_/A sky130_fd_sc_hd__buf_6
XTAP_3115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_104 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _431_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_420_ _420_/A_N _420_/B _420_/C vssd vssd vccd vccd _420_/X sky130_fd_sc_hd__and3b_4
XANTENNA_137 _547_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _221_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2029_A wire2029/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_351_ _351_/A _351_/B vssd vssd vccd vccd _351_/X sky130_fd_sc_hd__and2_4
XFILLER_42_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_282_ _282_/A _282_/B vssd vssd vccd vccd _282_/X sky130_fd_sc_hd__and2_4
XANTENNA__432__A_N _560_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input383_A la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__580__B _580_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input77_A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4036 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__101__A _101_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_618_ _618_/A _618_/B vssd vssd vccd vccd _618_/X sky130_fd_sc_hd__and2_4
XTAP_3693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1031_A _518_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1129_A _384_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_549_ _549_/A _549_/B vssd vssd vccd vccd _549_/X sky130_fd_sc_hd__and2_2
XFILLER_32_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output867_A _332_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1498_A wire1499/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__B _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1832_A wire1832/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[26\]_B _294_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__455__A_N _583_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__384__C _384_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput870 _307_/X vssd vssd vccd vccd mprj_adr_o_user[2] sky130_fd_sc_hd__buf_8
XFILLER_5_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput881 _114_/Y vssd vssd vccd vccd mprj_dat_i_core[0] sky130_fd_sc_hd__buf_8
XFILLER_1_4209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput892 _115_/Y vssd vssd vccd vccd mprj_dat_i_core[1] sky130_fd_sc_hd__buf_8
XFILLER_21_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1601 wire1601/A vssd vssd vccd vccd _603_/A sky130_fd_sc_hd__buf_6
XFILLER_5_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1612 wire1612/A vssd vssd vccd vccd _189_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1623 wire1623/A vssd vssd vccd vccd _450_/C sky130_fd_sc_hd__buf_6
XFILLER_8_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[17\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1634 wire1634/A vssd vssd vccd vccd _304_/A sky130_fd_sc_hd__buf_6
XFILLER_41_2161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1645 wire1645/A vssd vssd vccd vccd _389_/B sky130_fd_sc_hd__buf_6
XANTENNA_input131_A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1656 wire1656/A vssd vssd vccd vccd wire1656/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2146_A wire2147/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1667 wire1667/A vssd vssd vccd vccd wire1667/X sky130_fd_sc_hd__buf_6
XANTENNA_input229_A la_iena_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1678 wire1679/X vssd vssd vccd vccd _374_/B sky130_fd_sc_hd__buf_6
Xwire1689 wire1689/A vssd vssd vccd vccd wire1689/X sky130_fd_sc_hd__buf_6
XFILLER_34_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__575__B _575_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _531_/A _403_/B _403_/C vssd vssd vccd vccd _403_/X sky130_fd_sc_hd__and3b_4
XFILLER_26_182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_334_ _334_/A _334_/B vssd vssd vccd vccd _334_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__591__A _591_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_265_ _265_/A _265_/B vssd vssd vccd vccd _265_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire964 wire964/A vssd vssd vccd vccd _076_/A sky130_fd_sc_hd__buf_6
X_196_ _196_/A _196_/B vssd vssd vccd vccd _196_/X sky130_fd_sc_hd__and2_4
Xwire975 wire975/A vssd vssd vccd vccd _064_/A sky130_fd_sc_hd__buf_6
XFILLER_41_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire986 wire986/A vssd vssd vccd vccd _096_/A sky130_fd_sc_hd__buf_6
Xwire997 wire998/X vssd vssd vccd vccd wire997/X sky130_fd_sc_hd__buf_6
XFILLER_48_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1079_A _430_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__469__C _469_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_gates\[2\]_A user_irq_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1246_A wire1247/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__478__A_N _478_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__485__B _485_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1413_A wire1414/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3763 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_15 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_26 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_37 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_48 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1782_A wire1783/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_59 mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__006__A _006_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__379__C _379_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__395__B _395_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_050_ _050_/A vssd vssd vccd vccd _050_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_49_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2096_A wire2096/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input179_A la_iena_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input346_A la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2110 wire2111/X vssd vssd vccd vccd _481_/B sky130_fd_sc_hd__buf_6
Xwire2121 wire2122/X vssd vssd vccd vccd _476_/B sky130_fd_sc_hd__buf_6
Xwire2132 wire2132/A vssd vssd vccd vccd _470_/B sky130_fd_sc_hd__buf_6
XFILLER_1_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2143 wire2143/A vssd vssd vccd vccd _460_/B sky130_fd_sc_hd__buf_6
XFILLER_1_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2154 wire2154/A vssd vssd vccd vccd wire2154/X sky130_fd_sc_hd__buf_6
Xwire1420 wire1421/X vssd vssd vccd vccd wire1420/X sky130_fd_sc_hd__buf_6
Xwire2165 wire2166/X vssd vssd vccd vccd _451_/B sky130_fd_sc_hd__buf_6
Xwire1431 wire1431/A vssd vssd vccd vccd wire1431/X sky130_fd_sc_hd__buf_6
Xwire2176 wire2176/A vssd vssd vccd vccd wire2176/X sky130_fd_sc_hd__buf_6
XFILLER_5_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1442 wire1443/X vssd vssd vccd vccd _334_/B sky130_fd_sc_hd__buf_8
Xwire2187 wire2187/A vssd vssd vccd vccd wire2187/X sky130_fd_sc_hd__buf_6
Xwire1453 wire1454/X vssd vssd vccd vccd wire1453/X sky130_fd_sc_hd__buf_6
Xwire2198 wire2198/A vssd vssd vccd vccd _432_/B sky130_fd_sc_hd__buf_6
XFILLER_4_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__586__A _586_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1464 wire1465/X vssd vssd vccd vccd wire1464/X sky130_fd_sc_hd__buf_6
XFILLER_46_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1475 wire1476/X vssd vssd vccd vccd _327_/B sky130_fd_sc_hd__buf_6
Xwire1486 wire1487/X vssd vssd vccd vccd wire1486/X sky130_fd_sc_hd__buf_6
Xwire1497 wire1497/A vssd vssd vccd vccd wire1497/X sky130_fd_sc_hd__buf_6
XFILLER_46_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_317_ _317_/A _317_/B vssd vssd vccd vccd _317_/X sky130_fd_sc_hd__and2_1
XFILLER_50_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput13 la_data_out_mprj[108] vssd vssd vccd vccd _477_/C sky130_fd_sc_hd__clkbuf_4
Xinput24 la_data_out_mprj[118] vssd vssd vccd vccd _487_/C sky130_fd_sc_hd__buf_4
XFILLER_10_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_248_ _248_/A _248_/B vssd vssd vccd vccd _248_/X sky130_fd_sc_hd__and2_4
XFILLER_7_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput35 la_data_out_mprj[12] vssd vssd vccd vccd _381_/C sky130_fd_sc_hd__clkbuf_4
Xinput46 la_data_out_mprj[22] vssd vssd vccd vccd _391_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_output565_A _446_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput57 la_data_out_mprj[32] vssd vssd vccd vccd _401_/C sky130_fd_sc_hd__clkbuf_4
Xinput68 la_data_out_mprj[42] vssd vssd vccd vccd _411_/C sky130_fd_sc_hd__clkbuf_4
Xinput79 la_data_out_mprj[52] vssd vssd vccd vccd _421_/C sky130_fd_sc_hd__clkbuf_4
X_179_ _179_/A _179_/B vssd vssd vccd vccd _179_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1196_A wire1197/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output732_A _608_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] _240_/X vssd vssd vccd vccd _060_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_38_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1530_A wire1530/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1628_A wire1628/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1997_A wire1997/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire983_A wire983/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput406 mprj_adr_o_core[26] vssd vssd vccd vccd wire1461/A sky130_fd_sc_hd__buf_6
XFILLER_22_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput417 mprj_adr_o_core[7] vssd vssd vccd vccd wire1408/A sky130_fd_sc_hd__buf_6
Xinput428 mprj_dat_o_core[16] vssd vssd vccd vccd wire1378/A sky130_fd_sc_hd__buf_6
XFILLER_2_4359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput439 mprj_dat_o_core[26] vssd vssd vccd vccd wire1365/A sky130_fd_sc_hd__buf_6
XFILLER_9_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2109_A wire2109/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input296_A la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_102_ _102_/A vssd vssd vccd vccd _102_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_033_ _033_/A vssd vssd vccd vccd _033_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_4_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1250 _338_/X vssd vssd vccd vccd wire1250/X sky130_fd_sc_hd__buf_6
Xwire1261 _320_/X vssd vssd vccd vccd wire1261/X sky130_fd_sc_hd__buf_6
XFILLER_47_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1272 wire1273/X vssd vssd vccd vccd wire1272/X sky130_fd_sc_hd__buf_6
XFILLER_47_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1283 _304_/X vssd vssd vccd vccd wire1283/X sky130_fd_sc_hd__buf_6
Xwire1294 wire1295/X vssd vssd vccd vccd wire1294/X sky130_fd_sc_hd__buf_8
XFILLER_38_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1209_A wire1210/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output682_A _050_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__C _482_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output947_A wire1284/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1480_A wire1481/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1912_A wire1913/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] wire1316/X vssd vssd vccd vccd
+ wire992/A sky130_fd_sc_hd__nand2_2
XFILLER_26_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__392__C _392_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_B _294_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput203 la_iena_mprj[49] vssd vssd vccd vccd _212_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_gates\[9\]_B _172_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput214 la_iena_mprj[59] vssd vssd vccd vccd _222_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput225 la_iena_mprj[69] vssd vssd vccd vccd _232_/B sky130_fd_sc_hd__buf_4
XTAP_4702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput236 la_iena_mprj[79] vssd vssd vccd vccd _242_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput247 la_iena_mprj[89] vssd vssd vccd vccd _252_/B sky130_fd_sc_hd__clkbuf_4
Xinput258 la_iena_mprj[99] vssd vssd vccd vccd _262_/B sky130_fd_sc_hd__buf_4
XFILLER_5_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput269 la_oenb_mprj[108] vssd vssd vccd vccd _477_/A_N sky130_fd_sc_hd__buf_6
XFILLER_2_2721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2059_A wire2059/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input211_A la_iena_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_582_ _582_/A _582_/B vssd vssd vccd vccd _582_/X sky130_fd_sc_hd__and2_4
XFILLER_29_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input309_A la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__583__B _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_016_ _016_/A vssd vssd vccd vccd _016_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__104__A _104_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output528_A wire1101/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1061_A _474_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1159_A wire1160/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1080 _429_/X vssd vssd vccd vccd wire1080/X sky130_fd_sc_hd__buf_6
XFILLER_53_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1091 _421_/X vssd vssd vccd vccd wire1091/X sky130_fd_sc_hd__buf_6
XFILLER_1_2264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1326_A _251_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__493__B _493_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_740 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1695_A wire1695/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1738 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1862_A wire1862/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_308 wire2209/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_319 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_length1562_A _416_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input161_A la_iena_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2176_A wire2176/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input259_A la_iena_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__578__B _578_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input426_A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input22_A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__594__A _594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_565_ _565_/A _565_/B vssd vssd vccd vccd _565_/X sky130_fd_sc_hd__and2_4
XFILLER_2_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_496_ _624_/A _496_/B _496_/C vssd vssd vccd vccd _496_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output478_A _482_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput507 wire1120/X vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__buf_8
XFILLER_29_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput518 wire1110/X vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__buf_8
XFILLER_9_3439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput529 wire1100/X vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__buf_8
XANTENNA_output645_A _016_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1276_A _313_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output812_A _566_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__488__B _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1443_A wire1444/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1708_A wire1708/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3940 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_max_length1310_A _294_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__384__A_N _512_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__398__B _398_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1805 wire1805/A vssd vssd vccd vccd _250_/A sky130_fd_sc_hd__buf_4
XTAP_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1816 wire1816/A vssd vssd vccd vccd _333_/A sky130_fd_sc_hd__buf_6
XFILLER_28_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1827 wire1827/A vssd vssd vccd vccd _330_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1838 wire1838/A vssd vssd vccd vccd wire1838/X sky130_fd_sc_hd__buf_6
XFILLER_41_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1849 wire1849/A vssd vssd vccd vccd _177_/A sky130_fd_sc_hd__buf_6
XTAP_3105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_105 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _431_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _556_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_149 _210_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _350_/A _350_/B vssd vssd vccd vccd _350_/X sky130_fd_sc_hd__and2_4
XTAP_1758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_281_ _281_/A _281_/B vssd vssd vccd vccd _281_/X sky130_fd_sc_hd__and2_4
XFILLER_14_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input376_A la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4048 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__589__A _589_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_617_ _617_/A _617_/B vssd vssd vccd vccd _617_/X sky130_fd_sc_hd__and2_4
XFILLER_45_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_548_ _548_/A _548_/B vssd vssd vccd vccd _548_/X sky130_fd_sc_hd__and2_4
XTAP_2993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1024_A _530_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output595_A _086_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_479_ _479_/A_N _479_/B _479_/C vssd vssd vccd vccd _479_/X sky130_fd_sc_hd__and3b_2
XFILLER_31_2501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output762_A wire1029/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__C _490_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1393_A wire1393/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2430 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1658_A wire1658/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__499__A _499_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput860 wire1256/X vssd vssd vccd vccd mprj_adr_o_user[20] sky130_fd_sc_hd__buf_8
Xoutput871 _335_/X vssd vssd vccd vccd mprj_adr_o_user[30] sky130_fd_sc_hd__buf_8
XFILLER_5_3623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput882 _124_/Y vssd vssd vccd vccd mprj_dat_i_core[10] sky130_fd_sc_hd__buf_8
XFILLER_8_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput893 _134_/Y vssd vssd vccd vccd mprj_dat_i_core[20] sky130_fd_sc_hd__buf_8
XANTENNA__202__A _202_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1602 wire1602/A vssd vssd vccd vccd _602_/A sky130_fd_sc_hd__buf_6
XFILLER_8_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1613 wire1613/A vssd vssd vccd vccd _188_/B sky130_fd_sc_hd__buf_6
Xwire1624 wire1624/A vssd vssd vccd vccd _449_/C sky130_fd_sc_hd__buf_6
XFILLER_5_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1635 wire1636/X vssd vssd vccd vccd _394_/B sky130_fd_sc_hd__buf_6
Xwire1646 wire1647/X vssd vssd vccd vccd _388_/B sky130_fd_sc_hd__buf_6
XFILLER_19_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1657 wire1658/X vssd vssd vccd vccd _383_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1668 wire1669/X vssd vssd vccd vccd _378_/B sky130_fd_sc_hd__buf_6
Xwire1679 wire1679/A vssd vssd vccd vccd wire1679/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2041_A wire2041/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input124_A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2139_A wire2139/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ _530_/A _402_/B _402_/C vssd vssd vccd vccd _402_/X sky130_fd_sc_hd__and3b_2
XTAP_1522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_333_ _333_/A _333_/B vssd vssd vccd vccd _333_/X sky130_fd_sc_hd__and2_4
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__591__B _591_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_264_ _264_/A _264_/B vssd vssd vccd vccd _264_/X sky130_fd_sc_hd__and2_2
XFILLER_10_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_195_ _195_/A _195_/B vssd vssd vccd vccd _195_/X sky130_fd_sc_hd__and2_4
XFILLER_6_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire965 wire965/A vssd vssd vccd vccd _075_/A sky130_fd_sc_hd__buf_6
XFILLER_10_3875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire976 wire976/A vssd vssd vccd vccd _063_/A sky130_fd_sc_hd__buf_6
Xuser_wb_dat_gates\[5\] mprj_dat_i_user[5] max_length1311/X vssd vssd vccd vccd _119_/A
+ sky130_fd_sc_hd__nand2_4
Xwire987 wire987/A vssd vssd vccd vccd _095_/A sky130_fd_sc_hd__buf_6
Xwire998 _557_/X vssd vssd vccd vccd wire998/X sky130_fd_sc_hd__buf_6
XFILLER_48_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output510_A wire1117/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output608_A _098_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1141_A _373_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1239_A wire1240/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4410 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__485__C _485_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1406_A wire1407/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] _185_/X vssd vssd vccd vccd _005_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_32_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_16 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_27 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_38 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_49 mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1775_A wire1776/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1942_A wire1942/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__422__A_N _550_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1686 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__395__C _395_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2089_A wire2090/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2100 wire2101/X vssd vssd vccd vccd wire2100/X sky130_fd_sc_hd__buf_6
Xoutput690 _057_/Y vssd vssd vccd vccd la_data_in_mprj[74] sky130_fd_sc_hd__buf_8
Xwire2111 wire2111/A vssd vssd vccd vccd wire2111/X sky130_fd_sc_hd__buf_6
XFILLER_40_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input241_A la_iena_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2122 wire2122/A vssd vssd vccd vccd wire2122/X sky130_fd_sc_hd__buf_6
XFILLER_8_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2133 wire2134/X vssd vssd vccd vccd _469_/B sky130_fd_sc_hd__buf_6
XANTENNA_input339_A la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2144 wire2144/A vssd vssd vccd vccd _459_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1410 wire1411/X vssd vssd vccd vccd wire1410/X sky130_fd_sc_hd__buf_6
Xwire2155 wire2155/A vssd vssd vccd vccd _310_/A sky130_fd_sc_hd__buf_6
Xwire1421 wire1421/A vssd vssd vccd vccd wire1421/X sky130_fd_sc_hd__buf_6
Xwire2166 wire2166/A vssd vssd vccd vccd wire2166/X sky130_fd_sc_hd__buf_6
XFILLER_4_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1432 wire1433/X vssd vssd vccd vccd _335_/B sky130_fd_sc_hd__buf_8
Xwire2177 wire2178/X vssd vssd vccd vccd _445_/B sky130_fd_sc_hd__buf_6
XFILLER_38_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1443 wire1444/X vssd vssd vccd vccd wire1443/X sky130_fd_sc_hd__buf_6
XFILLER_21_2544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2188 wire2188/A vssd vssd vccd vccd _440_/B sky130_fd_sc_hd__buf_6
Xwire1454 wire1455/X vssd vssd vccd vccd wire1454/X sky130_fd_sc_hd__buf_6
Xwire2199 wire2199/A vssd vssd vccd vccd _307_/A sky130_fd_sc_hd__buf_6
Xwire1465 wire1466/X vssd vssd vccd vccd wire1465/X sky130_fd_sc_hd__buf_6
XFILLER_1_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1476 wire1476/A vssd vssd vccd vccd wire1476/X sky130_fd_sc_hd__buf_6
XANTENNA__586__B _586_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1487 wire1488/X vssd vssd vccd vccd wire1487/X sky130_fd_sc_hd__buf_6
Xwire1498 wire1499/X vssd vssd vccd vccd _322_/B sky130_fd_sc_hd__buf_6
XTAP_2020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_316_ _316_/A _316_/B vssd vssd vccd vccd _316_/X sky130_fd_sc_hd__and2_2
XFILLER_10_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__107__A _107_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput14 la_data_out_mprj[109] vssd vssd vccd vccd _478_/C sky130_fd_sc_hd__clkbuf_4
X_247_ _247_/A _247_/B vssd vssd vccd vccd _247_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput25 la_data_out_mprj[119] vssd vssd vccd vccd input25/X sky130_fd_sc_hd__buf_6
Xinput36 la_data_out_mprj[13] vssd vssd vccd vccd _382_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput47 la_data_out_mprj[23] vssd vssd vccd vccd _392_/C sky130_fd_sc_hd__clkbuf_4
Xinput58 la_data_out_mprj[33] vssd vssd vccd vccd _402_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput69 la_data_out_mprj[43] vssd vssd vccd vccd _412_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_13_1360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_178_ _178_/A _178_/B vssd vssd vccd vccd _178_/X sky130_fd_sc_hd__and2_4
XFILLER_7_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output558_A _439_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1091_A _421_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__445__A_N _573_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output725_A _602_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1356_A wire1357/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__496__B _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1523_A wire1524/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1892_A wire1893/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire976_A wire976/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_B _195_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput407 mprj_adr_o_core[27] vssd vssd vccd vccd wire1456/A sky130_fd_sc_hd__buf_6
XFILLER_6_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput418 mprj_adr_o_core[8] vssd vssd vccd vccd wire1404/A sky130_fd_sc_hd__buf_6
Xinput429 mprj_dat_o_core[17] vssd vssd vccd vccd wire1377/A sky130_fd_sc_hd__buf_6
XFILLER_22_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[99\]_B wire1317/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2004_A wire2004/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_101_ _101_/A vssd vssd vccd vccd _101_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_1393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input191_A la_iena_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input289_A la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_032_ _032_/A vssd vssd vccd vccd _032_/Y sky130_fd_sc_hd__inv_2
XANTENNA__468__A_N _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input456_A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input52_A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__597__A _597_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1240 _342_/X vssd vssd vccd vccd wire1240/X sky130_fd_sc_hd__buf_6
Xwire1251 wire1252/X vssd vssd vccd vccd wire1251/X sky130_fd_sc_hd__buf_6
XFILLER_21_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1262 wire1263/X vssd vssd vccd vccd wire1262/X sky130_fd_sc_hd__buf_6
XFILLER_40_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1273 _315_/X vssd vssd vccd vccd wire1273/X sky130_fd_sc_hd__buf_6
Xwire1284 wire1285/X vssd vssd vccd vccd wire1284/X sky130_fd_sc_hd__buf_8
XFILLER_1_2446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1295 wire1296/X vssd vssd vccd vccd wire1295/X sky130_fd_sc_hd__buf_8
XFILLER_47_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1104_A _409_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output842_A _593_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1473_A wire1474/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_B _177_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1640_A wire1640/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1738_A wire1739/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__300__A _300_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1905_A wire1906/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3802 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput204 la_iena_mprj[4] vssd vssd vccd vccd _167_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput215 la_iena_mprj[5] vssd vssd vccd vccd _168_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput226 la_iena_mprj[6] vssd vssd vccd vccd _169_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 la_iena_mprj[7] vssd vssd vccd vccd _170_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput248 la_iena_mprj[8] vssd vssd vccd vccd _171_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput259 la_iena_mprj[9] vssd vssd vccd vccd _172_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__210__A _210_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_581_ _581_/A _581_/B vssd vssd vccd vccd _581_/X sky130_fd_sc_hd__and2_4
XFILLER_44_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input204_A la_iena_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2121_A wire2122/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_015_ _015_/A vssd vssd vccd vccd _015_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__120__A _120_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1070 _465_/X vssd vssd vccd vccd wire1070/X sky130_fd_sc_hd__buf_6
Xwire1081 _428_/X vssd vssd vccd vccd wire1081/X sky130_fd_sc_hd__buf_6
XFILLER_47_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1092 _420_/X vssd vssd vccd vccd wire1092/X sky130_fd_sc_hd__buf_6
XFILLER_53_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1221_A wire1222/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output792_A wire1009/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1319_A _258_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__493__C _493_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3586 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1688_A wire1689/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1855_A wire1855/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_309 _380_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__205__A _205_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input154_A la_iena_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2071_A wire2072/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2169_A wire2170/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input321_A la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input419_A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_95 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__594__B _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_564_ _564_/A _564_/B vssd vssd vccd vccd _564_/X sky130_fd_sc_hd__and2_4
XTAP_3898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_495_ _623_/A _495_/B _495_/C vssd vssd vccd vccd _495_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2874 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput508 wire1119/X vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__buf_8
XFILLER_5_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput519 wire1109/X vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__buf_8
XFILLER_49_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output540_A wire1089/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output638_A _010_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1171_A wire1172/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_ack_gate mprj_ack_i_user max_length1310/X vssd vssd vccd vccd _146_/A sky130_fd_sc_hd__nand2_1
XANTENNA_wire1269_A wire1270/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__488__C _488_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output805_A _559_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1436_A wire1436/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] _215_/X vssd vssd vccd vccd _035_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_48_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3784 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1972_A wire1972/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__025__A _025_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3952 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[29\]_A mprj_dat_i_user[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1806 wire1806/A vssd vssd vccd vccd _249_/A sky130_fd_sc_hd__buf_4
XFILLER_41_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input7_A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__398__C _398_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1817 wire1817/A vssd vssd vccd vccd _332_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1828 wire1828/A vssd vssd vccd vccd _192_/A sky130_fd_sc_hd__buf_6
XTAP_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1839 wire1839/A vssd vssd vccd vccd _185_/A sky130_fd_sc_hd__buf_6
XFILLER_41_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_128 _431_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_139 _556_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_280_ _280_/A _280_/B vssd vssd vccd vccd _280_/X sky130_fd_sc_hd__and2_4
XFILLER_30_4140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input271_A la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input369_A la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__589__B _589_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_616_ _616_/A _616_/B vssd vssd vccd vccd _616_/X sky130_fd_sc_hd__and2_4
XTAP_3673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_547_ _547_/A _547_/B vssd vssd vccd vccd _547_/X sky130_fd_sc_hd__and2_2
XFILLER_35_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_478_ _478_/A_N _478_/B _478_/C vssd vssd vccd vccd _478_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output490_A _493_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output588_A wire1068/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output755_A wire1035/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2442 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output922_A wire1198/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__499__B _499_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1720_A wire1721/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput850 wire1268/X vssd vssd vccd vccd mprj_adr_o_user[11] sky130_fd_sc_hd__buf_8
XFILLER_25_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput861 _326_/X vssd vssd vccd vccd mprj_adr_o_user[21] sky130_fd_sc_hd__buf_8
XFILLER_47_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput872 _336_/X vssd vssd vccd vccd mprj_adr_o_user[31] sky130_fd_sc_hd__buf_8
XFILLER_5_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput883 _125_/Y vssd vssd vccd vccd mprj_dat_i_core[11] sky130_fd_sc_hd__buf_8
XFILLER_5_2901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput894 _135_/Y vssd vssd vccd vccd mprj_dat_i_core[21] sky130_fd_sc_hd__buf_8
XFILLER_43_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1603 wire1603/A vssd vssd vccd vccd _601_/A sky130_fd_sc_hd__buf_6
XFILLER_3_4071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1614 wire1614/A vssd vssd vccd vccd _187_/B sky130_fd_sc_hd__buf_6
Xwire1625 wire1625/A vssd vssd vccd vccd _448_/C sky130_fd_sc_hd__buf_6
XFILLER_8_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1636 wire1636/A vssd vssd vccd vccd wire1636/X sky130_fd_sc_hd__buf_6
Xwire1647 wire1647/A vssd vssd vccd vccd wire1647/X sky130_fd_sc_hd__buf_6
XFILLER_41_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1658 wire1658/A vssd vssd vccd vccd wire1658/X sky130_fd_sc_hd__buf_6
Xwire1669 wire1669/A vssd vssd vccd vccd wire1669/X sky130_fd_sc_hd__buf_6
XFILLER_19_4046 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input117_A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2034_A wire2034/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_401_ _529_/A _401_/B _401_/C vssd vssd vccd vccd _401_/X sky130_fd_sc_hd__and3b_2
XFILLER_15_3209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_332_ _332_/A _332_/B vssd vssd vccd vccd _332_/X sky130_fd_sc_hd__and2_4
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2201_A wire2202/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_263_ _263_/A _263_/B vssd vssd vccd vccd _263_/X sky130_fd_sc_hd__and2_4
XFILLER_6_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input82_A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_194_ _194_/A _194_/B vssd vssd vccd vccd _194_/X sky130_fd_sc_hd__and2_4
XFILLER_10_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire966 wire966/A vssd vssd vccd vccd _074_/A sky130_fd_sc_hd__buf_6
XFILLER_6_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire977 wire977/A vssd vssd vccd vccd _062_/A sky130_fd_sc_hd__buf_6
XFILLER_48_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire988 wire988/A vssd vssd vccd vccd _094_/A sky130_fd_sc_hd__buf_6
Xwire999 _556_/X vssd vssd vccd vccd wire999/X sky130_fd_sc_hd__buf_6
XFILLER_6_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output503_A wire1124/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__374__A_N _502_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1301_A wire1302/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output872_A _336_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_17 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[28\] mprj_dat_i_user[28] max_length1310/X vssd vssd vccd vccd
+ _142_/A sky130_fd_sc_hd__nand2_8
XFILLER_33_1918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_28 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] _178_/X vssd vssd vccd vccd _162_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA_39 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1670_A wire1671/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1768_A wire1768/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__303__A _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1935_A wire1936/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] _289_/X vssd vssd vccd vccd wire980/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_4244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__213__A _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4166 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput680 _048_/Y vssd vssd vccd vccd la_data_in_mprj[65] sky130_fd_sc_hd__buf_8
Xwire2101 wire2101/A vssd vssd vccd vccd wire2101/X sky130_fd_sc_hd__buf_6
XFILLER_27_2979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2112 wire2113/X vssd vssd vccd vccd _480_/B sky130_fd_sc_hd__buf_6
Xoutput691 _058_/Y vssd vssd vccd vccd la_data_in_mprj[75] sky130_fd_sc_hd__buf_8
XFILLER_43_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2123 wire2123/A vssd vssd vccd vccd _475_/B sky130_fd_sc_hd__buf_6
XFILLER_5_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2134 wire2134/A vssd vssd vccd vccd wire2134/X sky130_fd_sc_hd__buf_6
XFILLER_47_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1400 wire1400/A vssd vssd vccd vccd wire1400/X sky130_fd_sc_hd__buf_6
Xwire2145 wire2145/A vssd vssd vccd vccd _458_/B sky130_fd_sc_hd__buf_6
Xwire1411 wire1411/A vssd vssd vccd vccd wire1411/X sky130_fd_sc_hd__buf_6
Xwire2156 wire2157/X vssd vssd vccd vccd _454_/B sky130_fd_sc_hd__buf_6
Xwire1422 wire1423/X vssd vssd vccd vccd _308_/B sky130_fd_sc_hd__buf_6
Xwire2167 wire2168/X vssd vssd vccd vccd _450_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input234_A la_iena_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1433 wire1434/X vssd vssd vccd vccd wire1433/X sky130_fd_sc_hd__buf_6
XFILLER_19_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2178 wire2178/A vssd vssd vccd vccd wire2178/X sky130_fd_sc_hd__buf_6
XFILLER_4_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1444 wire1445/X vssd vssd vccd vccd wire1444/X sky130_fd_sc_hd__buf_6
XFILLER_38_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2189 wire2190/X vssd vssd vccd vccd _439_/B sky130_fd_sc_hd__buf_6
Xwire1455 wire1456/X vssd vssd vccd vccd wire1455/X sky130_fd_sc_hd__buf_6
Xwire1466 wire1466/A vssd vssd vccd vccd wire1466/X sky130_fd_sc_hd__buf_6
XFILLER_1_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1477 wire1478/X vssd vssd vccd vccd _326_/B sky130_fd_sc_hd__buf_6
XFILLER_19_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__397__A_N _525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1488 wire1489/X vssd vssd vccd vccd wire1488/X sky130_fd_sc_hd__buf_6
XFILLER_41_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1499 wire1500/X vssd vssd vccd vccd wire1499/X sky130_fd_sc_hd__buf_6
XTAP_2010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input401_A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_315_ _315_/A _315_/B vssd vssd vccd vccd _315_/X sky130_fd_sc_hd__and2_2
XTAP_1397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_246_ _246_/A _246_/B vssd vssd vccd vccd _246_/X sky130_fd_sc_hd__and2_4
Xinput15 la_data_out_mprj[10] vssd vssd vccd vccd _379_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput26 la_data_out_mprj[11] vssd vssd vccd vccd _380_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput37 la_data_out_mprj[14] vssd vssd vccd vccd _383_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput48 la_data_out_mprj[24] vssd vssd vccd vccd _393_/C sky130_fd_sc_hd__clkbuf_4
Xinput59 la_data_out_mprj[34] vssd vssd vccd vccd _403_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_177_ _177_/A _177_/B vssd vssd vccd vccd _177_/X sky130_fd_sc_hd__and2_4
XFILLER_13_1372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1084_A _426_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2478 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1251_A wire1252/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1349_A wire1349/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__496__C _496_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1516_A wire1517/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1885_A wire1885/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire969_A wire969/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__033__A _033_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput408 mprj_adr_o_core[28] vssd vssd vccd vccd wire1451/A sky130_fd_sc_hd__buf_6
XFILLER_44_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput419 mprj_adr_o_core[9] vssd vssd vccd vccd wire1400/A sky130_fd_sc_hd__buf_6
XFILLER_6_3785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__208__A _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_100_ _100_/A vssd vssd vccd vccd _100_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_031_ _031_/A vssd vssd vccd vccd _031_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input184_A la_iena_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2199_A wire2199/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input351_A la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input449_A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input45_A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__597__B _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1230 wire1231/X vssd vssd vccd vccd wire1230/X sky130_fd_sc_hd__buf_6
XFILLER_1_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1241 wire1242/X vssd vssd vccd vccd wire1241/X sky130_fd_sc_hd__buf_6
XFILLER_40_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1252 _337_/X vssd vssd vccd vccd wire1252/X sky130_fd_sc_hd__buf_6
XFILLER_21_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1263 _319_/X vssd vssd vccd vccd wire1263/X sky130_fd_sc_hd__buf_6
XFILLER_19_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1274 wire1275/X vssd vssd vccd vccd wire1274/X sky130_fd_sc_hd__buf_6
Xwire1285 wire1286/X vssd vssd vccd vccd wire1285/X sky130_fd_sc_hd__buf_8
Xwire1296 wire1297/X vssd vssd vccd vccd wire1296/X sky130_fd_sc_hd__buf_6
XFILLER_1_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__118__A _118_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__A_N _412_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output570_A _450_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_229_ _229_/A _229_/B vssd vssd vccd vccd _229_/X sky130_fd_sc_hd__and2_2
XANTENNA_wire1299_A wire1300/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output835_A wire1045/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1466_A wire1466/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] _245_/X vssd vssd vccd vccd _065_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3875 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__300__B _300_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3814 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput205 la_iena_mprj[50] vssd vssd vccd vccd _213_/B sky130_fd_sc_hd__clkbuf_4
Xinput216 la_iena_mprj[60] vssd vssd vccd vccd _223_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput227 la_iena_mprj[70] vssd vssd vccd vccd _233_/B sky130_fd_sc_hd__buf_4
XTAP_4704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput238 la_iena_mprj[80] vssd vssd vccd vccd _243_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput249 la_iena_mprj[90] vssd vssd vccd vccd _253_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__210__B _210_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_580_ _580_/A _580_/B vssd vssd vccd vccd _580_/X sky130_fd_sc_hd__and2_4
XFILLER_44_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__435__A_N _563_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input399_A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_786 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_014_ _014_/A vssd vssd vccd vccd _014_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_29_2805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3230 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1060 _475_/X vssd vssd vccd vccd wire1060/X sky130_fd_sc_hd__buf_6
Xwire1071 _464_/X vssd vssd vccd vccd wire1071/X sky130_fd_sc_hd__buf_6
Xwire1082 wire1083/X vssd vssd vccd vccd wire1082/X sky130_fd_sc_hd__buf_6
XFILLER_35_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1093 wire1094/X vssd vssd vccd vccd wire1093/X sky130_fd_sc_hd__buf_6
XFILLER_1_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1047_A _503_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1214_A wire1215/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output785_A wire1015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output952_A output952/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[10\] mprj_dat_i_user[10] _294_/X vssd vssd vccd vccd _124_/A sky130_fd_sc_hd__nand2_2
XFILLER_12_3598 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1750_A wire1750/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__458__A_N _586_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__205__B _205_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2064_A wire2065/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input147_A la_iena_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input314_A la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_563_ _563_/A _563_/B vssd vssd vccd vccd _563_/X sky130_fd_sc_hd__and2_4
XTAP_3888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_494_ _622_/A _494_/B _494_/C vssd vssd vccd vccd _494_/X sky130_fd_sc_hd__and3b_4
XFILLER_38_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2110 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2886 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput509 wire1118/X vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__buf_8
XFILLER_29_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output533_A wire1096/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__131__A _131_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1164_A wire1165/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1331_A _246_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1429_A wire1430/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] _208_/X vssd vssd vccd vccd _028_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_4355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1798_A wire1798/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__306__A _306_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1965_A wire1966/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] _170_/X vssd vssd vccd vccd _154_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_25_3756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[29\]_B max_length1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1807 wire1807/A vssd vssd vccd vccd _245_/A sky130_fd_sc_hd__buf_6
XFILLER_41_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1818 wire1818/A vssd vssd vccd vccd _208_/A sky130_fd_sc_hd__buf_4
XTAP_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1829 wire1829/A vssd vssd vccd vccd _191_/A sky130_fd_sc_hd__buf_6
XTAP_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_118 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_129 _431_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__216__A _216_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2181_A wire2181/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input264_A la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input431_A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2598 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_615_ _615_/A _615_/B vssd vssd vccd vccd _615_/X sky130_fd_sc_hd__and2_4
XTAP_3663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_546_ _546_/A _546_/B vssd vssd vccd vccd _546_/X sky130_fd_sc_hd__and2_2
XFILLER_45_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_477_ _477_/A_N _477_/B _477_/C vssd vssd vccd vccd _477_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output483_A _487_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__126__A _126_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output650_A _021_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output748_A _623_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1281_A wire1282/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1379_A wire1380/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output915_A wire1220/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1713_A wire1713/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire999_A _556_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_678 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__036__A _036_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput840 _591_/X vssd vssd vccd vccd la_oenb_core[94] sky130_fd_sc_hd__buf_8
XFILLER_5_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput851 wire1266/X vssd vssd vccd vccd mprj_adr_o_user[12] sky130_fd_sc_hd__buf_8
XFILLER_43_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput862 wire1254/X vssd vssd vccd vccd mprj_adr_o_user[22] sky130_fd_sc_hd__buf_8
XFILLER_8_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput873 _308_/X vssd vssd vccd vccd mprj_adr_o_user[3] sky130_fd_sc_hd__buf_8
Xoutput884 _126_/Y vssd vssd vccd vccd mprj_dat_i_core[12] sky130_fd_sc_hd__buf_8
XFILLER_21_3406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput895 _136_/Y vssd vssd vccd vccd mprj_dat_i_core[22] sky130_fd_sc_hd__buf_8
XFILLER_43_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1604 _472_/A_N vssd vssd vccd vccd _600_/A sky130_fd_sc_hd__buf_6
XFILLER_28_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1615 wire1615/A vssd vssd vccd vccd _186_/B sky130_fd_sc_hd__buf_6
XFILLER_3_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1626 wire1626/A vssd vssd vccd vccd _447_/C sky130_fd_sc_hd__buf_6
XTAP_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1637 wire1638/X vssd vssd vccd vccd _393_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1648 wire1649/X vssd vssd vccd vccd _387_/B sky130_fd_sc_hd__buf_6
Xwire1659 wire1660/X vssd vssd vccd vccd _382_/B sky130_fd_sc_hd__buf_6
XFILLER_19_4036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_400_ _400_/A_N _400_/B _400_/C vssd vssd vccd vccd _400_/X sky130_fd_sc_hd__and3b_2
XTAP_2247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2027_A wire2027/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_331_ _331_/A _331_/B vssd vssd vccd vccd _331_/X sky130_fd_sc_hd__and2_4
XFILLER_19_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_262_ _262_/A _262_/B vssd vssd vccd vccd _262_/X sky130_fd_sc_hd__and2_1
XFILLER_52_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input381_A la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_193_ _193_/A _193_/B vssd vssd vccd vccd _193_/X sky130_fd_sc_hd__and2_4
XFILLER_6_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire967 wire967/A vssd vssd vccd vccd _073_/A sky130_fd_sc_hd__buf_6
XANTENNA_input75_A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire978 wire978/A vssd vssd vccd vccd _061_/A sky130_fd_sc_hd__buf_6
XFILLER_6_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire989 wire989/A vssd vssd vccd vccd _093_/A sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1127_A _386_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_529_ _529_/A _529_/B vssd vssd vccd vccd _529_/X sky130_fd_sc_hd__and2_4
XTAP_2792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_18 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_29 mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output865_A _330_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1496_A wire1497/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1663_A wire1664/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__303__B _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1830_A wire1830/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1928_A wire1929/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] _282_/X vssd vssd vccd vccd _102_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__213__B _213_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput670 _039_/Y vssd vssd vccd vccd la_data_in_mprj[56] sky130_fd_sc_hd__buf_8
XFILLER_27_2958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput681 _049_/Y vssd vssd vccd vccd la_data_in_mprj[66] sky130_fd_sc_hd__buf_8
XFILLER_5_4178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2102 wire2103/X vssd vssd vccd vccd _484_/B sky130_fd_sc_hd__buf_6
Xoutput692 _059_/Y vssd vssd vccd vccd la_data_in_mprj[76] sky130_fd_sc_hd__buf_8
XFILLER_21_3203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2113 wire2114/X vssd vssd vccd vccd wire2113/X sky130_fd_sc_hd__buf_6
Xwire2124 wire2125/X vssd vssd vccd vccd _474_/B sky130_fd_sc_hd__buf_6
XFILLER_25_3394 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2135 wire2135/A vssd vssd vccd vccd _468_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1401 wire1402/X vssd vssd vccd vccd _313_/B sky130_fd_sc_hd__buf_6
Xwire2146 wire2147/X vssd vssd vccd vccd _457_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1412 wire1413/X vssd vssd vccd vccd _310_/B sky130_fd_sc_hd__buf_6
Xwire2157 wire2158/X vssd vssd vccd vccd wire2157/X sky130_fd_sc_hd__buf_6
XFILLER_28_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1423 wire1424/X vssd vssd vccd vccd wire1423/X sky130_fd_sc_hd__buf_6
Xwire2168 wire2168/A vssd vssd vccd vccd wire2168/X sky130_fd_sc_hd__buf_6
XFILLER_43_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1434 wire1435/X vssd vssd vccd vccd wire1434/X sky130_fd_sc_hd__buf_6
Xwire2179 wire2179/A vssd vssd vccd vccd _309_/A sky130_fd_sc_hd__buf_6
Xwire1445 wire1446/X vssd vssd vccd vccd wire1445/X sky130_fd_sc_hd__buf_6
XFILLER_4_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1456 wire1456/A vssd vssd vccd vccd wire1456/X sky130_fd_sc_hd__buf_6
XFILLER_38_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1467 wire1468/X vssd vssd vccd vccd _329_/B sky130_fd_sc_hd__buf_8
XANTENNA_input227_A la_iena_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1478 wire1479/X vssd vssd vccd vccd wire1478/X sky130_fd_sc_hd__buf_6
Xwire1489 wire1489/A vssd vssd vccd vccd wire1489/X sky130_fd_sc_hd__buf_6
XFILLER_28_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_314_ _314_/A _314_/B vssd vssd vccd vccd _314_/X sky130_fd_sc_hd__and2_4
XTAP_1387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_245_ _245_/A _245_/B vssd vssd vccd vccd _245_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput16 la_data_out_mprj[110] vssd vssd vccd vccd _479_/C sky130_fd_sc_hd__clkbuf_4
Xinput27 la_data_out_mprj[120] vssd vssd vccd vccd input27/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput38 la_data_out_mprj[15] vssd vssd vccd vccd _384_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_6_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput49 la_data_out_mprj[25] vssd vssd vccd vccd _394_/C sky130_fd_sc_hd__clkbuf_4
X_176_ _176_/A _176_/B vssd vssd vccd vccd _176_/X sky130_fd_sc_hd__and2_2
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1077_A _458_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1244_A wire1245/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1990 wire1991/X vssd vssd vccd vccd _579_/B sky130_fd_sc_hd__buf_6
XFILLER_18_450 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1411_A wire1411/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_494 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__491__A_N _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1509_A wire1510/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_290 _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1780_A wire1781/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1878_A wire1878/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_1484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput409 mprj_adr_o_core[29] vssd vssd vccd vccd wire1446/A sky130_fd_sc_hd__buf_6
XFILLER_25_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__208__B _208_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_030_ _030_/A vssd vssd vccd vccd _030_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__224__A _224_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input177_A la_iena_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2094_A wire2095/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input344_A la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input38_A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1220 wire1221/X vssd vssd vccd vccd wire1220/X sky130_fd_sc_hd__buf_6
XFILLER_1_3127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1231 _345_/X vssd vssd vccd vccd wire1231/X sky130_fd_sc_hd__buf_6
Xwire1242 wire1243/X vssd vssd vccd vccd wire1242/X sky130_fd_sc_hd__buf_6
XFILLER_5_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1253 _328_/X vssd vssd vccd vccd wire1253/X sky130_fd_sc_hd__buf_6
XFILLER_43_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1264 wire1265/X vssd vssd vccd vccd wire1264/X sky130_fd_sc_hd__buf_6
XFILLER_21_2365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1275 _314_/X vssd vssd vccd vccd wire1275/X sky130_fd_sc_hd__buf_6
Xwire1286 wire1287/X vssd vssd vccd vccd wire1286/X sky130_fd_sc_hd__buf_6
XFILLER_1_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1297 wire1298/X vssd vssd vccd vccd wire1297/X sky130_fd_sc_hd__buf_6
XFILLER_35_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_228_ _228_/A _228_/B vssd vssd vccd vccd _228_/X sky130_fd_sc_hd__and2_2
XFILLER_7_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_159_ _159_/A vssd vssd vccd vccd _159_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1194_A wire1195/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output730_A wire1042/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output828_A _580_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1361_A wire1361/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1459_A wire1460/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] _238_/X vssd vssd vccd vccd _058_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3887 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1626_A wire1626/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1947 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__309__A _309_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1995_A wire1995/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__044__A _044_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__387__A_N _515_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput206 la_iena_mprj[51] vssd vssd vccd vccd _214_/B sky130_fd_sc_hd__clkbuf_4
Xinput217 la_iena_mprj[61] vssd vssd vccd vccd _224_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput228 la_iena_mprj[71] vssd vssd vccd vccd _234_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput239 la_iena_mprj[81] vssd vssd vccd vccd _244_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2107_A wire2107/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_798 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input294_A la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_013_ _013_/A vssd vssd vccd vccd _013_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_29_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input461_A user_irq_ena[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1050 _500_/X vssd vssd vccd vccd wire1050/X sky130_fd_sc_hd__buf_6
XFILLER_2_3981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1061 _474_/X vssd vssd vccd vccd wire1061/X sky130_fd_sc_hd__buf_6
XFILLER_40_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1072 _463_/X vssd vssd vccd vccd wire1072/X sky130_fd_sc_hd__buf_6
XFILLER_38_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1083 _427_/X vssd vssd vccd vccd wire1083/X sky130_fd_sc_hd__buf_6
Xwire1094 _419_/X vssd vssd vccd vccd wire1094/X sky130_fd_sc_hd__buf_6
XFILLER_53_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__129__A _129_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1207_A _353_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output778_A wire1020/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output945_A wire1294/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1576_A wire1577/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__311__B _311_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1910_A wire1910/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] _264_/X vssd vssd vccd vccd _084_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__502__A _502_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2057_A wire2057/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__402__A_N _530_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1831 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_562_ _562_/A _562_/B vssd vssd vccd vccd _562_/X sky130_fd_sc_hd__and2_4
XTAP_3878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input307_A la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_493_ _621_/A _493_/B _493_/C vssd vssd vccd vccd _493_/X sky130_fd_sc_hd__and3b_4
XFILLER_44_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2898 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output526_A wire1103/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1157_A _366_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1324_A _253_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4476 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output895_A _136_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] _201_/X vssd vssd vccd vccd _021_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1693_A wire1693/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__306__B _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1860_A wire1860/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1958_A wire1958/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3932 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__322__A _322_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__425__A_N _553_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1808 wire1808/A vssd vssd vccd vccd _244_/A sky130_fd_sc_hd__buf_6
XTAP_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1819 wire1819/A vssd vssd vccd vccd _207_/A sky130_fd_sc_hd__buf_4
XTAP_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_108 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_119 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__216__B _216_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_728 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_B wire1332/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__232__A _232_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input257_A la_iena_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2174_A wire2174/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input424_A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input20_A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_614_ _614_/A _614_/B vssd vssd vccd vccd _614_/X sky130_fd_sc_hd__and2_4
XTAP_4398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_545_ _545_/A _545_/B vssd vssd vccd vccd _545_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_476_ _604_/A _476_/B _476_/C vssd vssd vccd vccd _476_/X sky130_fd_sc_hd__and3b_4
XFILLER_53_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output476_A wire1055/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[71\]_B _234_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__448__A_N _576_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output643_A _014_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__142__A _142_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1274_A wire1275/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1826 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output810_A _564_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1441_A wire1441/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1539_A wire1539/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_4251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1706_A wire1707/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput830 _582_/X vssd vssd vccd vccd la_oenb_core[85] sky130_fd_sc_hd__buf_8
XANTENNA__052__A _052_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput841 _592_/X vssd vssd vccd vccd la_oenb_core[95] sky130_fd_sc_hd__buf_8
XFILLER_25_3521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput852 wire1264/X vssd vssd vccd vccd mprj_adr_o_user[13] sky130_fd_sc_hd__buf_8
XFILLER_47_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput863 wire1253/X vssd vssd vccd vccd mprj_adr_o_user[23] sky130_fd_sc_hd__buf_8
Xoutput874 _309_/X vssd vssd vccd vccd mprj_adr_o_user[4] sky130_fd_sc_hd__buf_8
XFILLER_28_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput885 _127_/Y vssd vssd vccd vccd mprj_dat_i_core[13] sky130_fd_sc_hd__buf_8
Xoutput896 _137_/Y vssd vssd vccd vccd mprj_dat_i_core[23] sky130_fd_sc_hd__buf_8
XFILLER_43_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1605 wire1605/A vssd vssd vccd vccd _599_/A sky130_fd_sc_hd__buf_6
XFILLER_8_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1616 wire1616/A vssd vssd vccd vccd _457_/C sky130_fd_sc_hd__buf_6
XFILLER_5_2958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1627 wire1627/A vssd vssd vccd vccd _446_/C sky130_fd_sc_hd__buf_6
XTAP_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1638 wire1638/A vssd vssd vccd vccd wire1638/X sky130_fd_sc_hd__buf_6
XFILLER_19_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1649 wire1649/A vssd vssd vccd vccd wire1649/X sky130_fd_sc_hd__buf_6
XFILLER_6_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_330_ _330_/A _330_/B vssd vssd vccd vccd _330_/X sky130_fd_sc_hd__and2_4
XFILLER_26_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__227__A _227_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_261_ _261_/A _261_/B vssd vssd vccd vccd _261_/X sky130_fd_sc_hd__and2_4
XFILLER_17_2370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_192_ _192_/A _192_/B vssd vssd vccd vccd _192_/X sky130_fd_sc_hd__and2_2
XFILLER_48_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_2289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire968 wire968/A vssd vssd vccd vccd _072_/A sky130_fd_sc_hd__buf_6
Xwire979 wire979/A vssd vssd vccd vccd _110_/A sky130_fd_sc_hd__buf_6
XANTENNA_input374_A la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input68_A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_528_ _528_/A _528_/B vssd vssd vccd vccd _528_/X sky130_fd_sc_hd__and2_4
XFILLER_50_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1022_A wire1023/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output593_A _084_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__137__A _137_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_459_ _587_/A _459_/B _459_/C vssd vssd vccd vccd _459_/X sky130_fd_sc_hd__and3b_4
XANTENNA_19 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output760_A wire1031/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output858_A wire1257/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1391_A wire1392/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1656_A wire1656/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__600__A _600_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1823_A wire1823/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__047__A _047_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[35\]_B _198_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput660 _030_/Y vssd vssd vccd vccd la_data_in_mprj[47] sky130_fd_sc_hd__buf_8
XFILLER_40_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput671 _040_/Y vssd vssd vccd vccd la_data_in_mprj[57] sky130_fd_sc_hd__buf_8
Xoutput682 _050_/Y vssd vssd vccd vccd la_data_in_mprj[67] sky130_fd_sc_hd__buf_8
Xwire2103 wire2104/X vssd vssd vccd vccd wire2103/X sky130_fd_sc_hd__buf_6
Xoutput693 _060_/Y vssd vssd vccd vccd la_data_in_mprj[77] sky130_fd_sc_hd__buf_8
XFILLER_8_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2114 wire2114/A vssd vssd vccd vccd wire2114/X sky130_fd_sc_hd__buf_6
Xwire2125 wire2125/A vssd vssd vccd vccd wire2125/X sky130_fd_sc_hd__buf_6
XANTENNA__510__A _510_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2136 wire2136/A vssd vssd vccd vccd _467_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1402 wire1403/X vssd vssd vccd vccd wire1402/X sky130_fd_sc_hd__buf_6
XFILLER_21_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2147 wire2148/X vssd vssd vccd vccd wire2147/X sky130_fd_sc_hd__buf_6
Xwire1413 wire1414/X vssd vssd vccd vccd wire1413/X sky130_fd_sc_hd__buf_6
Xwire2158 wire2158/A vssd vssd vccd vccd wire2158/X sky130_fd_sc_hd__buf_6
XFILLER_25_2683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1424 wire1425/X vssd vssd vccd vccd wire1424/X sky130_fd_sc_hd__buf_6
Xwire2169 wire2170/X vssd vssd vccd vccd _449_/B sky130_fd_sc_hd__buf_6
Xwire1435 wire1436/X vssd vssd vccd vccd wire1435/X sky130_fd_sc_hd__buf_6
XFILLER_47_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1446 wire1446/A vssd vssd vccd vccd wire1446/X sky130_fd_sc_hd__buf_6
Xwire1457 wire1458/X vssd vssd vccd vccd _331_/B sky130_fd_sc_hd__buf_8
Xwire1468 wire1469/X vssd vssd vccd vccd wire1468/X sky130_fd_sc_hd__buf_6
Xwire1479 wire1480/X vssd vssd vccd vccd wire1479/X sky130_fd_sc_hd__buf_6
XFILLER_38_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input122_A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2137_A wire2138/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2919 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_313_ _313_/A _313_/B vssd vssd vccd vccd _313_/X sky130_fd_sc_hd__and2_2
XFILLER_35_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_244_ _244_/A _244_/B vssd vssd vccd vccd _244_/X sky130_fd_sc_hd__and2_4
XFILLER_10_340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput17 la_data_out_mprj[111] vssd vssd vccd vccd _480_/C sky130_fd_sc_hd__clkbuf_4
Xinput28 la_data_out_mprj[121] vssd vssd vccd vccd _490_/C sky130_fd_sc_hd__buf_4
XFILLER_10_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput39 la_data_out_mprj[16] vssd vssd vccd vccd _385_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_175_ _175_/A _175_/B vssd vssd vccd vccd _175_/X sky130_fd_sc_hd__and2_1
XFILLER_6_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[3\] mprj_dat_i_user[3] max_length1311/X vssd vssd vccd vccd _117_/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_in_gates\[110\]_B _273_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output606_A _096_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1980 wire1980/A vssd vssd vccd vccd wire1980/X sky130_fd_sc_hd__buf_6
Xwire1991 wire1991/A vssd vssd vccd vccd wire1991/X sky130_fd_sc_hd__buf_6
XFILLER_4_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1404_A wire1404/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1831 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_280 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] _183_/X vssd vssd vccd vccd _003_/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA_291 _611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1773_A wire1774/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[17\]_B _180_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__314__B _314_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1940_A wire1940/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__330__A _330_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2580 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[10\]_A mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__505__A _505_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3446 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2087_A wire2087/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__240__A _240_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput490 _493_/X vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__buf_8
XFILLER_43_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input337_A la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1210 _352_/X vssd vssd vccd vccd wire1210/X sky130_fd_sc_hd__buf_6
XFILLER_43_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1221 wire1222/X vssd vssd vccd vccd wire1221/X sky130_fd_sc_hd__buf_6
Xwire1232 wire1233/X vssd vssd vccd vccd wire1232/X sky130_fd_sc_hd__buf_6
XFILLER_38_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1243 _341_/X vssd vssd vccd vccd wire1243/X sky130_fd_sc_hd__buf_6
Xwire1254 wire1255/X vssd vssd vccd vccd wire1254/X sky130_fd_sc_hd__buf_6
XFILLER_19_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1265 _318_/X vssd vssd vccd vccd wire1265/X sky130_fd_sc_hd__buf_6
XFILLER_5_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1276 _313_/X vssd vssd vccd vccd wire1276/X sky130_fd_sc_hd__buf_6
XFILLER_38_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1287 wire1288/X vssd vssd vccd vccd wire1287/X sky130_fd_sc_hd__buf_6
Xwire1298 _301_/X vssd vssd vccd vccd wire1298/X sky130_fd_sc_hd__buf_6
XFILLER_34_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_227_ _227_/A _227_/B vssd vssd vccd vccd _227_/X sky130_fd_sc_hd__and2_2
XFILLER_45_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_158_ _158_/A vssd vssd vccd vccd _158_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output556_A _438_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_089_ _089_/A vssd vssd vccd vccd _089_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_wire1187_A wire1188/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output723_A _600_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1354_A wire1355/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] _231_/X vssd vssd vccd vccd _051_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_22_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1521_A wire1521/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1619_A wire1619/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__309__B _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1890_A wire1891/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1988_A wire1989/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire974_A wire974/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3859 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__060__A _060_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4066 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput207 la_iena_mprj[52] vssd vssd vccd vccd _215_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput218 la_iena_mprj[62] vssd vssd vccd vccd _225_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_41_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput229 la_iena_mprj[72] vssd vssd vccd vccd _235_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2747 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_958 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2002_A wire2002/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__235__A _235_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input287_A la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_012_ _012_/A vssd vssd vccd vccd _012_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_4_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input454_A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input50_A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__481__A_N _609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__401__C _401_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1040 _509_/X vssd vssd vccd vccd wire1040/X sky130_fd_sc_hd__buf_6
Xwire1051 _499_/X vssd vssd vccd vccd wire1051/X sky130_fd_sc_hd__buf_6
Xwire1062 _473_/X vssd vssd vccd vccd wire1062/X sky130_fd_sc_hd__buf_6
Xwire1073 _462_/X vssd vssd vccd vccd wire1073/X sky130_fd_sc_hd__buf_6
XFILLER_40_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1084 _426_/X vssd vssd vccd vccd wire1084/X sky130_fd_sc_hd__buf_6
XFILLER_35_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1095 _418_/X vssd vssd vccd vccd wire1095/X sky130_fd_sc_hd__buf_6
XFILLER_18_3913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1102_A _411_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__145__A _145_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output840_A _591_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output938_A wire1244/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1471_A wire1471/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1736_A wire1737/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1903_A wire1904/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__055__A _055_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2988 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__502__B _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_561_ _561_/A _561_/B vssd vssd vccd vccd _561_/X sky130_fd_sc_hd__and2_4
XTAP_3868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1854 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input202_A la_iena_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_492_ _620_/A _492_/B _492_/C vssd vssd vccd vccd _492_/X sky130_fd_sc_hd__and3b_4
XFILLER_44_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input98_A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__B _412_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output519_A wire1109/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1052_A _498_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__377__A_N _505_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3754 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output790_A wire1011/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_828 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3618 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1686_A wire1687/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__603__A _603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1853_A wire1853/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__322__B _322_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4222 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[2\]_A mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1809 wire1809/A vssd vssd vccd vccd _335_/A sky130_fd_sc_hd__buf_6
XTAP_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_109 mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__513__A _513_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__232__B _232_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input152_A la_iena_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2167_A wire2168/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input417_A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_613_ _613_/A _613_/B vssd vssd vccd vccd _613_/X sky130_fd_sc_hd__and2_4
XTAP_4388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_544_ _544_/A _544_/B vssd vssd vccd vccd _544_/X sky130_fd_sc_hd__and2_4
XTAP_3698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_475_ _603_/A _475_/B _475_/C vssd vssd vccd vccd _475_/X sky130_fd_sc_hd__and3b_4
XFILLER_15_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__407__B _407_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output469_A wire1061/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output636_A _008_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output803_A wire997/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1434_A wire1435/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput390 mprj_adr_o_core[11] vssd vssd vccd vccd wire1519/A sky130_fd_sc_hd__buf_6
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] _213_/X vssd vssd vccd vccd _033_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__317__B _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1970_A wire1970/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__333__A _333_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput820 _573_/X vssd vssd vccd vccd la_oenb_core[76] sky130_fd_sc_hd__buf_8
XFILLER_47_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput831 _583_/X vssd vssd vccd vccd la_oenb_core[86] sky130_fd_sc_hd__buf_8
XFILLER_9_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput842 _593_/X vssd vssd vccd vccd la_oenb_core[96] sky130_fd_sc_hd__buf_8
XFILLER_8_2005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput853 wire1262/X vssd vssd vccd vccd mprj_adr_o_user[14] sky130_fd_sc_hd__buf_8
XFILLER_25_3533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput864 _329_/X vssd vssd vccd vccd mprj_adr_o_user[24] sky130_fd_sc_hd__buf_8
XFILLER_43_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput875 _310_/X vssd vssd vccd vccd mprj_adr_o_user[5] sky130_fd_sc_hd__buf_8
Xoutput886 _128_/Y vssd vssd vccd vccd mprj_dat_i_core[14] sky130_fd_sc_hd__buf_8
Xoutput897 _138_/Y vssd vssd vccd vccd mprj_dat_i_core[24] sky130_fd_sc_hd__buf_8
XFILLER_25_3577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1606 wire1606/A vssd vssd vccd vccd _598_/A sky130_fd_sc_hd__buf_6
XANTENNA_input5_A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1617 wire1617/A vssd vssd vccd vccd _456_/C sky130_fd_sc_hd__buf_6
XTAP_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1628 wire1628/A vssd vssd vccd vccd _445_/C sky130_fd_sc_hd__buf_6
XTAP_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1639 wire1640/X vssd vssd vccd vccd _392_/B sky130_fd_sc_hd__buf_6
XFILLER_3_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__508__A _508_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__227__B _227_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_260_ _260_/A _260_/B vssd vssd vccd vccd _260_/X sky130_fd_sc_hd__and2_4
XFILLER_23_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_191_ _191_/A _191_/B vssd vssd vccd vccd _191_/X sky130_fd_sc_hd__and2_2
XFILLER_32_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire969 wire969/A vssd vssd vccd vccd _071_/A sky130_fd_sc_hd__buf_6
XFILLER_10_3879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__243__A _243_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input367_A la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_irq_gates\[2\] user_irq_core[2] _293_/X vssd vssd vccd vccd _113_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_527_ _527_/A _527_/B vssd vssd vccd vccd _527_/X sky130_fd_sc_hd__and2_2
XFILLER_15_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_458_ _586_/A _458_/B _458_/C vssd vssd vccd vccd _458_/X sky130_fd_sc_hd__and3b_4
XANTENNA__415__A_N _415_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output586_A wire1070/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_389_ _517_/A _389_/B _389_/C vssd vssd vccd vccd _389_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output753_A wire1037/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output920_A wire1205/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] _261_/X vssd vssd vccd vccd _081_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_29_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1649_A wire1649/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__600__B _600_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1816_A wire1816/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__063__A _063_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput650 _021_/Y vssd vssd vccd vccd la_data_in_mprj[38] sky130_fd_sc_hd__buf_8
Xoutput661 _031_/Y vssd vssd vccd vccd la_data_in_mprj[48] sky130_fd_sc_hd__buf_8
XFILLER_9_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput672 _041_/Y vssd vssd vccd vccd la_data_in_mprj[58] sky130_fd_sc_hd__buf_8
XFILLER_40_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput683 _051_/Y vssd vssd vccd vccd la_data_in_mprj[68] sky130_fd_sc_hd__buf_8
XFILLER_44_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2104 wire2104/A vssd vssd vccd vccd wire2104/X sky130_fd_sc_hd__buf_6
Xwire2115 wire2116/X vssd vssd vccd vccd _479_/B sky130_fd_sc_hd__buf_6
Xoutput694 _061_/Y vssd vssd vccd vccd la_data_in_mprj[78] sky130_fd_sc_hd__buf_8
XFILLER_8_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2126 wire2127/X vssd vssd vccd vccd _473_/B sky130_fd_sc_hd__buf_6
XANTENNA__510__B _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2137 wire2138/X vssd vssd vccd vccd _466_/B sky130_fd_sc_hd__buf_6
Xwire1403 wire1404/X vssd vssd vccd vccd wire1403/X sky130_fd_sc_hd__buf_6
Xwire2148 wire2148/A vssd vssd vccd vccd wire2148/X sky130_fd_sc_hd__buf_6
XFILLER_5_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1414 wire1415/X vssd vssd vccd vccd wire1414/X sky130_fd_sc_hd__buf_6
Xwire2159 wire2160/X vssd vssd vccd vccd _453_/B sky130_fd_sc_hd__buf_6
Xwire1425 wire1426/X vssd vssd vccd vccd wire1425/X sky130_fd_sc_hd__buf_6
XFILLER_25_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1436 wire1436/A vssd vssd vccd vccd wire1436/X sky130_fd_sc_hd__buf_6
Xwire1447 wire1448/X vssd vssd vccd vccd _333_/B sky130_fd_sc_hd__buf_8
XFILLER_3_3181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1458 wire1459/X vssd vssd vccd vccd wire1458/X sky130_fd_sc_hd__buf_6
Xwire1469 wire1470/X vssd vssd vccd vccd wire1469/X sky130_fd_sc_hd__buf_6
XFILLER_28_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2032_A wire2032/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input115_A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__438__A_N _566_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__238__A _238_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ _312_/A _312_/B vssd vssd vccd vccd _312_/X sky130_fd_sc_hd__and2_2
XFILLER_51_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_2488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_243_ _243_/A _243_/B vssd vssd vccd vccd _243_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput18 la_data_out_mprj[112] vssd vssd vccd vccd _481_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_input80_A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput29 la_data_out_mprj[122] vssd vssd vccd vccd _491_/C sky130_fd_sc_hd__clkbuf_4
X_174_ _174_/A _174_/B vssd vssd vccd vccd _174_/X sky130_fd_sc_hd__and2_2
XFILLER_6_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__404__C _404_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__420__B _420_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1690 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1970 wire1970/A vssd vssd vccd vccd wire1970/X sky130_fd_sc_hd__buf_6
XFILLER_19_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output501_A wire1125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1981 wire1982/X vssd vssd vccd vccd _583_/B sky130_fd_sc_hd__buf_6
XFILLER_37_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1992 wire1993/X vssd vssd vccd vccd _578_/B sky130_fd_sc_hd__buf_6
XFILLER_15_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1132_A _381_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_270 _215_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_281 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_292 wire1707/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] _176_/X vssd vssd vccd vccd _160_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[26\] mprj_dat_i_user[26] _294_/X vssd vssd vccd vccd _140_/A sky130_fd_sc_hd__nand2_4
XFILLER_14_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1599_A _477_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1766_A wire1766/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__611__A _611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__330__B _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] wire1312/X vssd vssd vccd vccd
+ _107_/A sky130_fd_sc_hd__nand2_8
XFILLER_42_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__058__A _058_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[10\]_B _294_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__505__B _505_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__521__A _521_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput480 _484_/X vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__buf_8
Xoutput491 _494_/X vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__buf_8
XFILLER_40_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__240__B _240_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1200 wire1201/X vssd vssd vccd vccd wire1200/X sky130_fd_sc_hd__buf_6
Xwire1211 wire1212/X vssd vssd vccd vccd wire1211/X sky130_fd_sc_hd__buf_6
XFILLER_43_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1222 _348_/X vssd vssd vccd vccd wire1222/X sky130_fd_sc_hd__buf_6
Xwire1233 wire1234/X vssd vssd vccd vccd wire1233/X sky130_fd_sc_hd__buf_6
XANTENNA_input232_A la_iena_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1244 wire1245/X vssd vssd vccd vccd wire1244/X sky130_fd_sc_hd__buf_6
XFILLER_5_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1255 _327_/X vssd vssd vccd vccd wire1255/X sky130_fd_sc_hd__buf_6
Xwire1266 wire1267/X vssd vssd vccd vccd wire1266/X sky130_fd_sc_hd__buf_6
Xwire1277 _312_/X vssd vssd vccd vccd wire1277/X sky130_fd_sc_hd__buf_6
XFILLER_35_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1288 _303_/X vssd vssd vccd vccd wire1288/X sky130_fd_sc_hd__buf_6
Xwire1299 wire1300/X vssd vssd vccd vccd wire1299/X sky130_fd_sc_hd__buf_8
XFILLER_38_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_226_ _226_/A _226_/B vssd vssd vccd vccd _226_/X sky130_fd_sc_hd__and2_2
XANTENNA__415__B _415_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_157_ _157_/A vssd vssd vccd vccd _157_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_6_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_088_ _088_/A vssd vssd vccd vccd _088_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output549_A wire1078/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1082_A wire1083/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output716_A _081_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1347_A wire1347/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__606__A _606_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1883_A wire1884/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__325__B _325_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire967_A wire967/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__341__A _341_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4034 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput208 la_iena_mprj[53] vssd vssd vccd vccd _216_/B sky130_fd_sc_hd__clkbuf_4
Xinput219 la_iena_mprj[63] vssd vssd vccd vccd _226_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1251 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__516__A _516_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__235__B _235_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_011_ _011_/A vssd vssd vccd vccd _011_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_46_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input182_A la_iena_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2197_A wire2197/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__251__A _251_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3266 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input447_A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input43_A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1030 _519_/X vssd vssd vccd vccd wire1030/X sky130_fd_sc_hd__buf_6
XFILLER_7_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1041 _508_/X vssd vssd vccd vccd wire1041/X sky130_fd_sc_hd__buf_6
XFILLER_2_3961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_856 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1052 _498_/X vssd vssd vccd vccd wire1052/X sky130_fd_sc_hd__buf_6
XFILLER_38_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1063 _472_/X vssd vssd vccd vccd wire1063/X sky130_fd_sc_hd__buf_6
Xwire1074 _461_/X vssd vssd vccd vccd wire1074/X sky130_fd_sc_hd__buf_6
Xwire1085 wire1086/X vssd vssd vccd vccd wire1085/X sky130_fd_sc_hd__buf_6
XFILLER_1_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1096 _417_/X vssd vssd vccd vccd wire1096/X sky130_fd_sc_hd__buf_6
XFILLER_1_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output499_A wire1127/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_209_ _209_/A _209_/B vssd vssd vccd vccd _209_/X sky130_fd_sc_hd__and2_1
XFILLER_32_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1297_A wire1298/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output833_A _585_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__161__A _161_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1464_A wire1465/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] wire1332/X vssd vssd vccd vccd wire976/A
+ sky130_fd_sc_hd__nand2_4
XTAP_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1806 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1631_A wire1631/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1729_A wire1730/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__336__A _336_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__071__A _071_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1070 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_560_ _560_/A _560_/B vssd vssd vccd vccd _560_/X sky130_fd_sc_hd__and2_4
XTAP_3858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_491_ _619_/A _491_/B _491_/C vssd vssd vccd vccd _491_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2112_A wire2113/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__246__A _246_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input397_A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__C _412_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4470 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1045_A _505_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3766 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1212_A wire1213/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output783_A wire1016/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__156__A _156_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output950_A wire1299/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1679_A wire1679/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__603__B _603_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1846_A wire1846/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[2\]_B max_length1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__471__A_N _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__066__A _066_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__513__B _513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2062_A wire2063/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input145_A la_iena_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_612_ _612_/A _612_/B vssd vssd vccd vccd _612_/X sky130_fd_sc_hd__and2_4
XTAP_4378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input312_A la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_543_ _543_/A _543_/B vssd vssd vccd vccd _543_/X sky130_fd_sc_hd__and2_4
XTAP_2932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_474_ _602_/A _474_/B _474_/C vssd vssd vccd vccd _474_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_4320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__423__B _423_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output531_A wire1098/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1162_A wire1163/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput380 la_oenb_mprj[93] vssd vssd vccd vccd _590_/A sky130_fd_sc_hd__buf_8
XFILLER_42_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput391 mprj_adr_o_core[12] vssd vssd vccd vccd wire1517/A sky130_fd_sc_hd__buf_6
XFILLER_36_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1427_A wire1428/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__494__A_N _622_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] _206_/X vssd vssd vccd vccd _026_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_3530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1090 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__614__A _614_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1963_A wire1964/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__333__B _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput810 _564_/X vssd vssd vccd vccd la_oenb_core[67] sky130_fd_sc_hd__buf_8
Xoutput821 _574_/X vssd vssd vccd vccd la_oenb_core[77] sky130_fd_sc_hd__buf_8
Xoutput832 _584_/X vssd vssd vccd vccd la_oenb_core[87] sky130_fd_sc_hd__buf_8
XFILLER_47_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput843 _594_/X vssd vssd vccd vccd la_oenb_core[97] sky130_fd_sc_hd__buf_8
XFILLER_9_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput854 wire1261/X vssd vssd vccd vccd mprj_adr_o_user[15] sky130_fd_sc_hd__buf_8
Xoutput865 _330_/X vssd vssd vccd vccd mprj_adr_o_user[25] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] _168_/X vssd vssd vccd vccd _152_/A
+ sky130_fd_sc_hd__nand2_2
Xoutput876 wire1278/X vssd vssd vccd vccd mprj_adr_o_user[6] sky130_fd_sc_hd__buf_8
XFILLER_8_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput887 _129_/Y vssd vssd vccd vccd mprj_dat_i_core[15] sky130_fd_sc_hd__buf_8
XFILLER_28_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput898 _139_/Y vssd vssd vccd vccd mprj_dat_i_core[25] sky130_fd_sc_hd__buf_8
XFILLER_25_3589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1607 wire1607/A vssd vssd vccd vccd _597_/A sky130_fd_sc_hd__buf_6
XTAP_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1618 wire1618/A vssd vssd vccd vccd _455_/C sky130_fd_sc_hd__buf_6
XFILLER_3_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1629 wire1629/A vssd vssd vccd vccd _444_/C sky130_fd_sc_hd__buf_6
XTAP_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__508__B _508_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_190_ _190_/A _190_/B vssd vssd vccd vccd _190_/X sky130_fd_sc_hd__and2_1
XFILLER_10_3836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_394 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__524__A _524_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_41_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__243__B _243_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input262_A la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__418__B _418_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_526_ _526_/A _526_/B vssd vssd vccd vccd _526_/X sky130_fd_sc_hd__and2_4
XFILLER_50_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_457_ _585_/A _457_/B _457_/C vssd vssd vccd vccd _457_/X sky130_fd_sc_hd__and3b_4
XFILLER_53_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_388_ _516_/A _388_/B _388_/C vssd vssd vccd vccd _388_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output481_A _485_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output579_A wire1137/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output746_A _621_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1377_A wire1377/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output913_A wire1251/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1544_A wire1544/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1711_A wire1711/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1809_A wire1809/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__609__A _609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__328__B _328_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire997_A wire998/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__344__A _344_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_10_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput640 _012_/Y vssd vssd vccd vccd la_data_in_mprj[29] sky130_fd_sc_hd__buf_8
XFILLER_5_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput651 _022_/Y vssd vssd vccd vccd la_data_in_mprj[39] sky130_fd_sc_hd__buf_8
XFILLER_25_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput662 _032_/Y vssd vssd vccd vccd la_data_in_mprj[49] sky130_fd_sc_hd__buf_8
XFILLER_25_3353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput673 _042_/Y vssd vssd vccd vccd la_data_in_mprj[59] sky130_fd_sc_hd__buf_8
Xoutput684 _052_/Y vssd vssd vccd vccd la_data_in_mprj[69] sky130_fd_sc_hd__buf_8
Xwire2105 wire2106/X vssd vssd vccd vccd _483_/B sky130_fd_sc_hd__buf_6
XFILLER_40_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput695 _062_/Y vssd vssd vccd vccd la_data_in_mprj[79] sky130_fd_sc_hd__buf_8
Xwire2116 wire2116/A vssd vssd vccd vccd wire2116/X sky130_fd_sc_hd__buf_6
XFILLER_47_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2127 wire2127/A vssd vssd vccd vccd wire2127/X sky130_fd_sc_hd__buf_6
Xwire2138 wire2138/A vssd vssd vccd vccd wire2138/X sky130_fd_sc_hd__buf_6
Xwire1404 wire1404/A vssd vssd vccd vccd wire1404/X sky130_fd_sc_hd__buf_6
XFILLER_21_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2149 wire2150/X vssd vssd vccd vccd _456_/B sky130_fd_sc_hd__buf_6
Xwire1415 wire1416/X vssd vssd vccd vccd wire1415/X sky130_fd_sc_hd__buf_6
Xwire1426 wire1426/A vssd vssd vccd vccd wire1426/X sky130_fd_sc_hd__buf_6
XFILLER_8_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1437 wire1438/X vssd vssd vccd vccd _307_/B sky130_fd_sc_hd__buf_8
XFILLER_47_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1448 wire1449/X vssd vssd vccd vccd wire1448/X sky130_fd_sc_hd__buf_6
Xwire1459 wire1460/X vssd vssd vccd vccd wire1459/X sky130_fd_sc_hd__buf_6
XFILLER_28_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__519__A _519_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__238__B _238_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input108_A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_311_ _311_/A _311_/B vssd vssd vccd vccd _311_/X sky130_fd_sc_hd__and2_4
XTAP_1368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_242_ _242_/A _242_/B vssd vssd vccd vccd _242_/X sky130_fd_sc_hd__and2_2
XFILLER_52_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__254__A _254_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput19 la_data_out_mprj[113] vssd vssd vccd vccd _482_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_7_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_173_ _173_/A _173_/B vssd vssd vccd vccd _173_/X sky130_fd_sc_hd__and2_1
XFILLER_32_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input73_A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__420__C _420_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1960 wire1961/X vssd vssd vccd vccd wire1960/X sky130_fd_sc_hd__buf_6
Xwire1971 wire1971/A vssd vssd vccd vccd _590_/B sky130_fd_sc_hd__buf_6
XFILLER_20_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1982 wire1983/X vssd vssd vccd vccd wire1982/X sky130_fd_sc_hd__buf_6
XFILLER_4_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1993 wire1993/A vssd vssd vccd vccd wire1993/X sky130_fd_sc_hd__buf_6
XTAP_3260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1125_A _388_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_260 _470_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_271 _216_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_282 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_509_ _509_/A _509_/B vssd vssd vccd vccd _509_/X sky130_fd_sc_hd__and2_4
XFILLER_37_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_293 wire1754/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output863_A wire1253/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__164__A _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[19\] mprj_dat_i_user[19] max_length1311/X vssd vssd vccd vccd
+ _133_/A sky130_fd_sc_hd__nand2_4
XFILLER_31_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1494_A wire1495/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1661_A wire1662/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1759_A wire1760/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__611__B _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1926_A wire1927/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] _280_/X vssd vssd vccd vccd wire983/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__074__A _074_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3986 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__521__B _521_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput470 wire1060/X vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__buf_8
XFILLER_44_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput481 _485_/X vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__buf_8
XFILLER_47_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput492 _495_/X vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__buf_8
XFILLER_40_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__405__A_N _405_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1201 _355_/X vssd vssd vccd vccd wire1201/X sky130_fd_sc_hd__buf_6
XFILLER_25_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1212 wire1213/X vssd vssd vccd vccd wire1212/X sky130_fd_sc_hd__buf_6
Xwire1223 wire1224/X vssd vssd vccd vccd wire1223/X sky130_fd_sc_hd__buf_6
XFILLER_43_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1234 _344_/X vssd vssd vccd vccd wire1234/X sky130_fd_sc_hd__buf_6
Xwire1245 _340_/X vssd vssd vccd vccd wire1245/X sky130_fd_sc_hd__buf_6
XFILLER_1_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1256 _325_/X vssd vssd vccd vccd wire1256/X sky130_fd_sc_hd__buf_6
XFILLER_21_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2142_A wire2142/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input225_A la_iena_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1267 _317_/X vssd vssd vccd vccd wire1267/X sky130_fd_sc_hd__buf_6
XFILLER_47_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1278 wire1279/X vssd vssd vccd vccd wire1278/X sky130_fd_sc_hd__buf_6
XFILLER_21_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1289 wire1290/X vssd vssd vccd vccd wire1289/X sky130_fd_sc_hd__buf_8
XFILLER_34_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__249__A _249_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_225_ _225_/A _225_/B vssd vssd vccd vccd _225_/X sky130_fd_sc_hd__and2_2
XFILLER_11_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__415__C _415_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_156_ _156_/A vssd vssd vccd vccd _156_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_087_ _087_/A vssd vssd vccd vccd _087_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_49_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__B _431_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1075_A _460_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output611_A _101_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output709_A _074_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1242_A wire1243/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1790 wire1790/A vssd vssd vccd vccd wire1790/X sky130_fd_sc_hd__buf_6
XFILLER_0_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1507_A wire1508/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4064 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__606__B _606_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1876_A wire1877/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__622__A _622_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__341__B _341_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__428__A_N _556_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4046 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput209 la_iena_mprj[54] vssd vssd vccd vccd _217_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__069__A _069_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__516__B _516_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_010_ _010_/A vssd vssd vccd vccd _010_/Y sky130_fd_sc_hd__inv_4
XFILLER_10_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__532__A _532_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2092_A wire2093/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input175_A la_iena_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3278 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input342_A la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input36_A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1020 wire1021/X vssd vssd vccd vccd wire1020/X sky130_fd_sc_hd__buf_6
XFILLER_0_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1031 _518_/X vssd vssd vccd vccd wire1031/X sky130_fd_sc_hd__buf_6
XFILLER_1_2204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1042 wire1043/X vssd vssd vccd vccd wire1042/X sky130_fd_sc_hd__buf_6
Xwire1053 _497_/X vssd vssd vccd vccd wire1053/X sky130_fd_sc_hd__buf_6
XFILLER_5_2395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1064 _471_/X vssd vssd vccd vccd wire1064/X sky130_fd_sc_hd__buf_6
XFILLER_53_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1075 _460_/X vssd vssd vccd vccd wire1075/X sky130_fd_sc_hd__buf_6
Xwire1086 _425_/X vssd vssd vccd vccd wire1086/X sky130_fd_sc_hd__buf_6
Xwire1097 _416_/X vssd vssd vccd vccd wire1097/X sky130_fd_sc_hd__buf_6
XFILLER_35_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_208_ _208_/A _208_/B vssd vssd vccd vccd _208_/X sky130_fd_sc_hd__and2_1
XFILLER_45_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output561_A _442_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output659_A _029_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_139_ _139_/A vssd vssd vccd vccd _139_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1192_A wire1193/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output826_A _578_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3790 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1457_A wire1458/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] _236_/X vssd vssd vccd vccd _056_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1624_A wire1624/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1046 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__617__A _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1993_A wire1993/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__336__B _336_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2924 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[92\]_B wire1322/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__352__A _352_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2430 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_490_ _618_/A _490_/B _490_/C vssd vssd vccd vccd _490_/X sky130_fd_sc_hd__and3b_4
XANTENNA__527__A _527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2105_A wire2106/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input292_A la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[83\]_B wire1331/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__262__A _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xmax_length1562 _416_/A_N vssd vssd vccd vccd wire1561/A sky130_fd_sc_hd__buf_6
XFILLER_4_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1038_A _511_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_562 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1205_A wire1206/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output776_A _533_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[74\]_B _237_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output943_A wire1229/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__172__A _172_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1741_A wire1741/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1839_A wire1839/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1058 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__347__A _347_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__082__A _082_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input138_A la_iena_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2055_A wire2056/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_611_ _611_/A _611_/B vssd vssd vccd vccd _611_/X sky130_fd_sc_hd__and2_4
XFILLER_29_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_542_ _542_/A _542_/B vssd vssd vccd vccd _542_/X sky130_fd_sc_hd__and2_2
XTAP_3678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input305_A la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__257__A _257_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_473_ _601_/A _473_/B _473_/C vssd vssd vccd vccd _473_/X sky130_fd_sc_hd__and3b_4
XFILLER_44_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__423__C _423_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3810 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output524_A wire1142/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3854 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1155_A wire1156/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput370 la_oenb_mprj[84] vssd vssd vccd vccd wire1533/A sky130_fd_sc_hd__buf_6
Xinput381 la_oenb_mprj[94] vssd vssd vccd vccd _591_/A sky130_fd_sc_hd__buf_6
XFILLER_7_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput392 mprj_adr_o_core[13] vssd vssd vccd vccd wire1514/A sky130_fd_sc_hd__buf_6
XFILLER_40_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1322_A _255_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__167__A _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] _199_/X vssd vssd vccd vccd _019_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_36_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1691_A wire1691/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1789_A wire1790/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__614__B _614_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1956_A wire1956/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput800 wire1000/X vssd vssd vccd vccd la_oenb_core[58] sky130_fd_sc_hd__buf_8
Xoutput811 _565_/X vssd vssd vccd vccd la_oenb_core[68] sky130_fd_sc_hd__buf_8
XFILLER_9_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput822 _575_/X vssd vssd vccd vccd la_oenb_core[78] sky130_fd_sc_hd__buf_8
Xoutput833 _585_/X vssd vssd vccd vccd la_oenb_core[88] sky130_fd_sc_hd__buf_8
Xoutput844 _595_/X vssd vssd vccd vccd la_oenb_core[98] sky130_fd_sc_hd__buf_8
Xoutput855 wire1260/X vssd vssd vccd vccd mprj_adr_o_user[16] sky130_fd_sc_hd__buf_8
XFILLER_47_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput866 _331_/X vssd vssd vccd vccd mprj_adr_o_user[26] sky130_fd_sc_hd__buf_8
XFILLER_25_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput877 wire1277/X vssd vssd vccd vccd mprj_adr_o_user[7] sky130_fd_sc_hd__buf_8
XFILLER_5_3629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput888 _130_/Y vssd vssd vccd vccd mprj_dat_i_core[16] sky130_fd_sc_hd__buf_8
XFILLER_28_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput899 _140_/Y vssd vssd vccd vccd mprj_dat_i_core[26] sky130_fd_sc_hd__buf_8
XFILLER_25_2834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1608 input25/X vssd vssd vccd vccd _488_/C sky130_fd_sc_hd__buf_6
XTAP_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1619 wire1619/A vssd vssd vccd vccd _454_/C sky130_fd_sc_hd__buf_6
XFILLER_3_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__077__A _077_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_B _201_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__524__B _524_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_B _285_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__540__A _540_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2172_A wire2172/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input255_A la_iena_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input422_A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[31\]_A mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_525_ _525_/A _525_/B vssd vssd vccd vccd _525_/X sky130_fd_sc_hd__and2_4
XTAP_2752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__418__C _418_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_456_ _584_/A _456_/B _456_/C vssd vssd vccd vccd _456_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_387_ _515_/A _387_/B _387_/C vssd vssd vccd vccd _387_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[29\]_B _192_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__434__B _434_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_B _276_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output474_A wire1135/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output739_A _615_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1272_A wire1273/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__461__A_N _589_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1537_A wire1537/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__609__B _609_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1704_A wire1705/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[22\]_A mprj_dat_i_user[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__625__A _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__344__B _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[104\]_B _267_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput630 _148_/Y vssd vssd vccd vccd la_data_in_mprj[1] sky130_fd_sc_hd__buf_8
XANTENNA__360__A _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput641 _149_/Y vssd vssd vccd vccd la_data_in_mprj[2] sky130_fd_sc_hd__buf_8
Xoutput652 _150_/Y vssd vssd vccd vccd la_data_in_mprj[3] sky130_fd_sc_hd__buf_8
XFILLER_47_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput663 _151_/Y vssd vssd vccd vccd la_data_in_mprj[4] sky130_fd_sc_hd__buf_8
XFILLER_9_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput674 _152_/Y vssd vssd vccd vccd la_data_in_mprj[5] sky130_fd_sc_hd__buf_8
XFILLER_25_3365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput685 _153_/Y vssd vssd vccd vccd la_data_in_mprj[6] sky130_fd_sc_hd__buf_8
Xwire2106 wire2107/X vssd vssd vccd vccd wire2106/X sky130_fd_sc_hd__buf_6
Xoutput696 _154_/Y vssd vssd vccd vccd la_data_in_mprj[7] sky130_fd_sc_hd__buf_8
Xwire2117 wire2118/X vssd vssd vccd vccd _478_/B sky130_fd_sc_hd__buf_6
Xwire2128 wire2129/X vssd vssd vccd vccd _472_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2139 wire2139/A vssd vssd vccd vccd _465_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1405 wire1406/X vssd vssd vccd vccd _312_/B sky130_fd_sc_hd__buf_6
Xwire1416 wire1416/A vssd vssd vccd vccd wire1416/X sky130_fd_sc_hd__buf_6
Xwire1427 wire1428/X vssd vssd vccd vccd _336_/B sky130_fd_sc_hd__buf_6
XFILLER_3_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1438 wire1439/X vssd vssd vccd vccd wire1438/X sky130_fd_sc_hd__buf_6
XFILLER_41_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1449 wire1450/X vssd vssd vccd vccd wire1449/X sky130_fd_sc_hd__buf_6
XFILLER_39_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__519__B _519_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[13\]_A mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ _310_/A _310_/B vssd vssd vccd vccd _310_/X sky130_fd_sc_hd__and2_4
XFILLER_42_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2018_A wire2018/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__535__A _535_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_241_ _241_/A _241_/B vssd vssd vccd vccd _241_/X sky130_fd_sc_hd__and2_4
XFILLER_51_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__254__B _254_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_172_ _172_/A _172_/B vssd vssd vccd vccd _172_/X sky130_fd_sc_hd__and2_4
XFILLER_49_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input372_A la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__484__A_N _612_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input66_A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__270__A _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1950 wire1951/X vssd vssd vccd vccd _598_/B sky130_fd_sc_hd__buf_6
Xwire1961 wire1962/X vssd vssd vccd vccd wire1961/X sky130_fd_sc_hd__buf_6
Xwire1972 wire1972/A vssd vssd vccd vccd _589_/B sky130_fd_sc_hd__buf_6
XFILLER_18_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1983 wire1983/A vssd vssd vccd vccd wire1983/X sky130_fd_sc_hd__buf_6
XFILLER_18_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1994 wire1995/X vssd vssd vccd vccd _577_/B sky130_fd_sc_hd__buf_6
XTAP_3250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_250 _539_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_261 _469_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_508_ _508_/A _508_/B vssd vssd vccd vccd _508_/X sky130_fd_sc_hd__and2_4
XANTENNA_272 wire1667/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1020_A wire1021/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_283 _352_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1118_A _395_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_294 wire1756/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output689_A _056_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_439_ _567_/A _439_/B _439_/C vssd vssd vccd vccd _439_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output856_A wire1258/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1487_A wire1488/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__180__A _180_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1654_A wire1654/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1919_A wire1920/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__339__B _339_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__355__A _355_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__090__A _090_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput471 wire1059/X vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__buf_8
XFILLER_9_3392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput482 _486_/X vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__buf_8
Xoutput493 _496_/X vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__buf_8
XFILLER_5_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1202 wire1203/X vssd vssd vccd vccd wire1202/X sky130_fd_sc_hd__buf_6
XFILLER_43_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1213 _351_/X vssd vssd vccd vccd wire1213/X sky130_fd_sc_hd__buf_6
XFILLER_47_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1224 wire1225/X vssd vssd vccd vccd wire1224/X sky130_fd_sc_hd__buf_6
Xwire1235 wire1236/X vssd vssd vccd vccd wire1235/X sky130_fd_sc_hd__buf_6
Xwire1246 wire1247/X vssd vssd vccd vccd wire1246/X sky130_fd_sc_hd__buf_6
XFILLER_5_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1257 _324_/X vssd vssd vccd vccd wire1257/X sky130_fd_sc_hd__buf_6
Xwire1268 wire1269/X vssd vssd vccd vccd wire1268/X sky130_fd_sc_hd__buf_6
XFILLER_38_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1279 _311_/X vssd vssd vccd vccd wire1279/X sky130_fd_sc_hd__buf_6
XFILLER_1_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input120_A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2135_A wire2135/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input218_A la_iena_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__265__A _265_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_224_ _224_/A _224_/B vssd vssd vccd vccd _224_/X sky130_fd_sc_hd__and2_2
XFILLER_7_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_155_ _155_/A vssd vssd vccd vccd _155_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[1\] mprj_dat_i_user[1] max_length1310/X vssd vssd vccd vccd _115_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_45_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_086_ _086_/A vssd vssd vccd vccd _086_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__C _431_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1068_A _467_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output604_A _094_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1780 wire1781/X vssd vssd vccd vccd _268_/A sky130_fd_sc_hd__buf_6
XANTENNA_wire1235_A wire1236/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1791 wire1792/X vssd vssd vccd vccd _262_/A sky130_fd_sc_hd__buf_6
XFILLER_18_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1402_A wire1403/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1642 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__175__A _175_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[31\] mprj_dat_i_user[31] max_length1310/X vssd vssd vccd vccd
+ _145_/A sky130_fd_sc_hd__nand2_8
XFILLER_37_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1771_A wire1772/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1869_A wire1870/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__622__B _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__085__A _085_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2730 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2085_A wire2086/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input168_A la_iena_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input335_A la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1010 _547_/X vssd vssd vccd vccd wire1010/X sky130_fd_sc_hd__buf_6
Xwire1021 _535_/X vssd vssd vccd vccd wire1021/X sky130_fd_sc_hd__buf_6
Xwire1032 _517_/X vssd vssd vccd vccd wire1032/X sky130_fd_sc_hd__buf_6
Xwire1043 _507_/X vssd vssd vccd vccd wire1043/X sky130_fd_sc_hd__buf_6
XFILLER_47_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input29_A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1054 _481_/X vssd vssd vccd vccd wire1054/X sky130_fd_sc_hd__buf_6
Xwire1065 _470_/X vssd vssd vccd vccd wire1065/X sky130_fd_sc_hd__buf_6
XFILLER_1_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1076 _459_/X vssd vssd vccd vccd wire1076/X sky130_fd_sc_hd__buf_6
Xwire1087 wire1088/X vssd vssd vccd vccd wire1087/X sky130_fd_sc_hd__buf_6
XFILLER_5_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1098 _415_/X vssd vssd vccd vccd wire1098/X sky130_fd_sc_hd__buf_6
XFILLER_18_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__426__C _426_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_207_ _207_/A _207_/B vssd vssd vccd vccd _207_/X sky130_fd_sc_hd__and2_1
XFILLER_50_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_138_ _138_/A vssd vssd vccd vccd _138_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__442__B _442_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output554_A _436_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_069_ _069_/A vssd vssd vccd vccd _069_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output721_A _598_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output819_A _572_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1352_A wire1353/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] _229_/X vssd vssd vccd vccd _049_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_1_3440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1617_A wire1617/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__617__B _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1986_A wire1987/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire972_A wire972/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__352__B _352_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[5\]_A mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__543__A _543_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input285_A la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__262__B _262_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input452_A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4494 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__437__B _437_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_574 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__418__A_N _546_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1100_A _413_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output769_A wire1051/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4418 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output936_A wire1150/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3936 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1567_A _406_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1734_A wire1734/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1901_A wire1901/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_828 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__347__B _347_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__363__A _363_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_4169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_610_ _610_/A _610_/B vssd vssd vccd vccd _610_/X sky130_fd_sc_hd__and2_4
XTAP_4358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2048_A wire2048/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__538__A _538_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_541_ _541_/A _541_/B vssd vssd vccd vccd _541_/X sky130_fd_sc_hd__and2_2
XTAP_2912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input200_A la_iena_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__257__B _257_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_472_ _472_/A_N _472_/B _472_/C vssd vssd vccd vccd _472_/X sky130_fd_sc_hd__and3b_4
XTAP_2978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input96_A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__273__A _273_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3866 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output517_A wire1111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput360 la_oenb_mprj[75] vssd vssd vccd vccd wire1542/A sky130_fd_sc_hd__buf_6
XFILLER_42_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput371 la_oenb_mprj[85] vssd vssd vccd vccd wire1532/A sky130_fd_sc_hd__buf_6
XFILLER_23_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput382 la_oenb_mprj[95] vssd vssd vccd vccd _592_/A sky130_fd_sc_hd__buf_8
XANTENNA_wire1050_A _500_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1148_A wire1149/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput393 mprj_adr_o_core[14] vssd vssd vccd vccd wire1511/A sky130_fd_sc_hd__buf_6
XFILLER_36_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] _192_/X vssd vssd vccd vccd _012_/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA__390__A_N _518_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__183__A _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1684_A wire1685/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput801 wire999/X vssd vssd vccd vccd la_oenb_core[59] sky130_fd_sc_hd__buf_8
XFILLER_25_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput812 _566_/X vssd vssd vccd vccd la_oenb_core[69] sky130_fd_sc_hd__buf_8
XANTENNA_wire1851_A wire1851/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput823 _576_/X vssd vssd vccd vccd la_oenb_core[79] sky130_fd_sc_hd__buf_8
XFILLER_9_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1949_A wire1949/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput834 wire995/X vssd vssd vccd vccd la_oenb_core[89] sky130_fd_sc_hd__buf_8
Xoutput845 _596_/X vssd vssd vccd vccd la_oenb_core[99] sky130_fd_sc_hd__buf_8
XFILLER_8_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput856 wire1258/X vssd vssd vccd vccd mprj_adr_o_user[17] sky130_fd_sc_hd__buf_8
Xoutput867 _332_/X vssd vssd vccd vccd mprj_adr_o_user[27] sky130_fd_sc_hd__buf_8
XFILLER_9_3788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput878 wire1276/X vssd vssd vccd vccd mprj_adr_o_user[8] sky130_fd_sc_hd__buf_8
XFILLER_47_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput889 _131_/Y vssd vssd vccd vccd mprj_dat_i_core[17] sky130_fd_sc_hd__buf_8
XFILLER_3_4033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1609 wire1609/A vssd vssd vccd vccd _231_/B sky130_fd_sc_hd__buf_4
XTAP_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__358__A _358_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3930 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__093__A _093_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input150_A la_iena_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2165_A wire2166/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input248_A la_iena_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input415_A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input11_A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__268__A _268_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[31\]_B max_length1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_524_ _524_/A _524_/B vssd vssd vccd vccd _524_/X sky130_fd_sc_hd__and2_4
XTAP_2742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_455_ _583_/A _455_/B _455_/C vssd vssd vccd vccd _455_/X sky130_fd_sc_hd__and3b_4
XTAP_2797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_386_ _514_/A _386_/B _386_/C vssd vssd vccd vccd _386_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__434__C _434_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output467_A wire1063/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1098_A _415_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__450__B _450_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output634_A _006_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1265_A _318_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2052 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output801_A wire999/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1432_A wire1433/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput190 la_iena_mprj[37] vssd vssd vccd vccd _200_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_37_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__178__A _178_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_B max_length1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1899_A wire1900/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1294 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput620 _109_/Y vssd vssd vccd vccd la_data_in_mprj[126] sky130_fd_sc_hd__buf_8
XFILLER_47_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput631 _003_/Y vssd vssd vccd vccd la_data_in_mprj[20] sky130_fd_sc_hd__buf_8
XFILLER_9_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__360__B _360_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput642 _013_/Y vssd vssd vccd vccd la_data_in_mprj[30] sky130_fd_sc_hd__buf_8
XFILLER_47_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput653 _023_/Y vssd vssd vccd vccd la_data_in_mprj[40] sky130_fd_sc_hd__buf_8
XFILLER_47_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput664 _033_/Y vssd vssd vccd vccd la_data_in_mprj[50] sky130_fd_sc_hd__buf_8
XFILLER_28_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput675 _043_/Y vssd vssd vccd vccd la_data_in_mprj[60] sky130_fd_sc_hd__buf_8
XFILLER_9_3596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput686 _053_/Y vssd vssd vccd vccd la_data_in_mprj[70] sky130_fd_sc_hd__buf_8
Xwire2107 wire2107/A vssd vssd vccd vccd wire2107/X sky130_fd_sc_hd__buf_6
Xoutput697 _063_/Y vssd vssd vccd vccd la_data_in_mprj[80] sky130_fd_sc_hd__buf_8
Xwire2118 wire2118/A vssd vssd vccd vccd wire2118/X sky130_fd_sc_hd__buf_6
XFILLER_25_2643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2129 wire2129/A vssd vssd vccd vccd wire2129/X sky130_fd_sc_hd__buf_6
XFILLER_28_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input3_A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1406 wire1407/X vssd vssd vccd vccd wire1406/X sky130_fd_sc_hd__buf_6
Xwire1417 wire1418/X vssd vssd vccd vccd _309_/B sky130_fd_sc_hd__buf_8
XFILLER_47_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1428 wire1429/X vssd vssd vccd vccd wire1428/X sky130_fd_sc_hd__buf_6
Xwire1439 wire1440/X vssd vssd vccd vccd wire1439/X sky130_fd_sc_hd__buf_6
XFILLER_3_3173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__088__A _088_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[13\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_240_ _240_/A _240_/B vssd vssd vccd vccd _240_/X sky130_fd_sc_hd__and2_4
XANTENNA__535__B _535_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_171_ _171_/A _171_/B vssd vssd vccd vccd _171_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input198_A la_iena_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__551__A _551_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input365_A la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_510 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_irq_gates\[0\] user_irq_core[0] _291_/X vssd vssd vccd vccd _111_/A sky130_fd_sc_hd__nand2_1
XANTENNA_input59_A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4410 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1940 wire1940/A vssd vssd vccd vccd wire1940/X sky130_fd_sc_hd__buf_6
XFILLER_4_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1951 wire1952/X vssd vssd vccd vccd wire1951/X sky130_fd_sc_hd__buf_6
XFILLER_19_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1962 wire1962/A vssd vssd vccd vccd wire1962/X sky130_fd_sc_hd__buf_6
Xwire1973 wire1974/X vssd vssd vccd vccd _588_/B sky130_fd_sc_hd__buf_6
Xwire1984 wire1985/X vssd vssd vccd vccd _582_/B sky130_fd_sc_hd__buf_6
XTAP_3240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__429__C _429_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1995 wire1995/A vssd vssd vccd vccd wire1995/X sky130_fd_sc_hd__buf_6
XFILLER_19_967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_240 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 _539_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_262 wire2134/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_507_ _507_/A _507_/B vssd vssd vccd vccd _507_/X sky130_fd_sc_hd__and2_2
XFILLER_19_3693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_273 wire1645/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_284 _351_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_295 _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__445__B _445_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1013_A wire1014/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_438_ _566_/A _438_/B _438_/C vssd vssd vccd vccd _438_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output584_A wire1072/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_369_ _497_/A _369_/B _369_/C vssd vssd vccd vccd _369_/X sky130_fd_sc_hd__and3b_4
XFILLER_18_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output751_A wire1039/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output849_A wire1271/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] wire1318/X vssd vssd vccd vccd _079_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_4387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1647_A wire1647/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__355__B _355_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput472 wire1058/X vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__buf_8
XFILLER_47_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput483 _487_/X vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__buf_8
Xoutput494 wire1132/X vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__buf_8
XFILLER_5_3257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1203 wire1204/X vssd vssd vccd vccd wire1203/X sky130_fd_sc_hd__buf_6
Xwire1214 wire1215/X vssd vssd vccd vccd wire1214/X sky130_fd_sc_hd__buf_6
XFILLER_5_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1225 _347_/X vssd vssd vccd vccd wire1225/X sky130_fd_sc_hd__buf_6
XFILLER_47_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1236 wire1237/X vssd vssd vccd vccd wire1236/X sky130_fd_sc_hd__buf_6
XFILLER_1_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1247 wire1248/X vssd vssd vccd vccd wire1247/X sky130_fd_sc_hd__buf_6
XFILLER_5_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1258 wire1259/X vssd vssd vccd vccd wire1258/X sky130_fd_sc_hd__buf_6
XFILLER_21_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1269 wire1270/X vssd vssd vccd vccd wire1269/X sky130_fd_sc_hd__buf_6
XFILLER_38_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2030_A wire2030/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input113_A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2128_A wire2129/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__546__A _546_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__265__B _265_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__451__A_N _579_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_223_ _223_/A _223_/B vssd vssd vccd vccd _223_/X sky130_fd_sc_hd__and2_2
XFILLER_50_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_154_ _154_/A vssd vssd vccd vccd _154_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__281__A _281_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_085_ _085_/A vssd vssd vccd vccd _085_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1770 wire1770/A vssd vssd vccd vccd wire1770/X sky130_fd_sc_hd__buf_6
XFILLER_4_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1781 wire1781/A vssd vssd vccd vccd wire1781/X sky130_fd_sc_hd__buf_6
XFILLER_53_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1792 wire1792/A vssd vssd vccd vccd wire1792/X sky130_fd_sc_hd__buf_6
XFILLER_15_4000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1130_A _383_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1228_A _346_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output799_A _554_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] _174_/X vssd vssd vccd vccd _158_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_15_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_gates\[24\] mprj_dat_i_user[24] _294_/X vssd vssd vccd vccd _138_/A sky130_fd_sc_hd__nand2_4
XFILLER_50_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1597_A _478_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__191__A _191_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1764_A wire1764/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1931_A wire1932/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1046 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] _285_/X vssd vssd vccd vccd wire982/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_6_2876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__474__A_N _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__366__A _366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2078_A wire2078/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1000 wire1001/X vssd vssd vccd vccd wire1000/X sky130_fd_sc_hd__buf_6
Xwire1011 wire1012/X vssd vssd vccd vccd wire1011/X sky130_fd_sc_hd__buf_6
XFILLER_40_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1022 wire1023/X vssd vssd vccd vccd wire1022/X sky130_fd_sc_hd__buf_6
XANTENNA_input230_A la_iena_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1033 _516_/X vssd vssd vccd vccd wire1033/X sky130_fd_sc_hd__buf_6
XANTENNA_input328_A la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1044 _506_/X vssd vssd vccd vccd wire1044/X sky130_fd_sc_hd__buf_6
XFILLER_2_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1055 _480_/X vssd vssd vccd vccd wire1055/X sky130_fd_sc_hd__buf_6
XFILLER_53_4509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1066 _469_/X vssd vssd vccd vccd wire1066/X sky130_fd_sc_hd__buf_6
XFILLER_2_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1077 _458_/X vssd vssd vccd vccd wire1077/X sky130_fd_sc_hd__buf_6
Xwire1088 _424_/X vssd vssd vccd vccd wire1088/X sky130_fd_sc_hd__buf_6
Xwire1099 _414_/X vssd vssd vccd vccd wire1099/X sky130_fd_sc_hd__buf_6
XFILLER_28_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__276__A _276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_206_ _206_/A _206_/B vssd vssd vccd vccd _206_/X sky130_fd_sc_hd__and2_1
XFILLER_10_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_137_ _137_/A vssd vssd vccd vccd _137_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_8_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2550 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__442__C _442_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_068_ _068_/A vssd vssd vccd vccd _068_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output547_A wire1080/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1080_A _429_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1178_A wire1179/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output714_A _079_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1345_A wire1345/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] _222_/X vssd vssd vccd vccd _042_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_2740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1512_A wire1513/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1716 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__186__A _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1881_A wire1882/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1979_A wire1980/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[5\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__096__A _096_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__543__B _543_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input180_A la_iena_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2195_A wire2195/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input278_A la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input445_A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input41_A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__437__C _437_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output497_A wire1129/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__453__B _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1295_A wire1296/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output831_A _583_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output929_A wire1174/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1462_A wire1463/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1727_A wire1728/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__363__B _363_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__538__B _538_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_540_ _540_/A _540_/B vssd vssd vccd vccd _540_/X sky130_fd_sc_hd__and2_4
XTAP_2913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_471_ _599_/A _471_/B _471_/C vssd vssd vccd vccd _471_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2110_A wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2208_A wire2209/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__554__A _554_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input395_A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__273__B _273_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input89_A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput350 la_oenb_mprj[66] vssd vssd vccd vccd wire1551/A sky130_fd_sc_hd__buf_6
Xinput361 la_oenb_mprj[76] vssd vssd vccd vccd wire1541/A sky130_fd_sc_hd__buf_6
Xinput372 la_oenb_mprj[86] vssd vssd vccd vccd wire1531/A sky130_fd_sc_hd__buf_6
XFILLER_40_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput383 la_oenb_mprj[96] vssd vssd vccd vccd _593_/A sky130_fd_sc_hd__buf_6
XFILLER_48_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput394 mprj_adr_o_core[15] vssd vssd vccd vccd wire1508/A sky130_fd_sc_hd__buf_6
XFILLER_53_4103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__448__B _448_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1210_A _352_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output781_A _537_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1308_A wire1309/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output879_A wire1274/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3198 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput802 wire1048/X vssd vssd vccd vccd la_oenb_core[5] sky130_fd_sc_hd__buf_8
Xoutput813 wire1047/X vssd vssd vccd vccd la_oenb_core[6] sky130_fd_sc_hd__buf_8
Xoutput824 wire1046/X vssd vssd vccd vccd la_oenb_core[7] sky130_fd_sc_hd__buf_8
XFILLER_25_4249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput835 wire1045/X vssd vssd vccd vccd la_oenb_core[8] sky130_fd_sc_hd__buf_8
XFILLER_6_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput846 wire1044/X vssd vssd vccd vccd la_oenb_core[9] sky130_fd_sc_hd__buf_8
XFILLER_29_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput857 _323_/X vssd vssd vccd vccd mprj_adr_o_user[18] sky130_fd_sc_hd__buf_8
XFILLER_5_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1844_A wire1844/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput868 _333_/X vssd vssd vccd vccd mprj_adr_o_user[28] sky130_fd_sc_hd__buf_8
XFILLER_42_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput879 wire1274/X vssd vssd vccd vccd mprj_adr_o_user[9] sky130_fd_sc_hd__buf_8
XTAP_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2104 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__358__B _358_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_52_2244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input143_A la_iena_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2060_A wire2061/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2158_A wire2158/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1886 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__549__A _549_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__268__B _268_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input310_A la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input408_A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_523_ _523_/A _523_/B vssd vssd vccd vccd _523_/X sky130_fd_sc_hd__and2_4
XFILLER_22_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_454_ _582_/A _454_/B _454_/C vssd vssd vccd vccd _454_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__284__A _284_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_385_ _513_/A _385_/B _385_/C vssd vssd vccd vccd _385_/X sky130_fd_sc_hd__and3b_4
XFILLER_9_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__450__C _450_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3879 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1160_A wire1161/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_4229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1258_A wire1259/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput180 la_iena_mprj[28] vssd vssd vccd vccd _191_/B sky130_fd_sc_hd__buf_4
XFILLER_42_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput191 la_iena_mprj[38] vssd vssd vccd vccd _201_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__178__B _178_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1425_A wire1426/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] _204_/X vssd vssd vccd vccd _024_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__194__A _194_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1961_A wire1962/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput610 _100_/Y vssd vssd vccd vccd la_data_in_mprj[117] sky130_fd_sc_hd__buf_8
Xoutput621 _110_/Y vssd vssd vccd vccd la_data_in_mprj[127] sky130_fd_sc_hd__buf_8
Xoutput632 _004_/Y vssd vssd vccd vccd la_data_in_mprj[21] sky130_fd_sc_hd__buf_8
Xoutput643 _014_/Y vssd vssd vccd vccd la_data_in_mprj[31] sky130_fd_sc_hd__buf_8
XFILLER_9_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput654 _024_/Y vssd vssd vccd vccd la_data_in_mprj[41] sky130_fd_sc_hd__buf_8
XFILLER_5_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput665 _034_/Y vssd vssd vccd vccd la_data_in_mprj[51] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] _166_/X vssd vssd vccd vccd _150_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_47_1656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput676 _044_/Y vssd vssd vccd vccd la_data_in_mprj[61] sky130_fd_sc_hd__buf_8
XFILLER_28_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2108 wire2109/X vssd vssd vccd vccd _482_/B sky130_fd_sc_hd__buf_6
Xoutput687 _054_/Y vssd vssd vccd vccd la_data_in_mprj[71] sky130_fd_sc_hd__buf_8
Xoutput698 _064_/Y vssd vssd vccd vccd la_data_in_mprj[81] sky130_fd_sc_hd__buf_8
Xwire2119 wire2120/X vssd vssd vccd vccd _477_/B sky130_fd_sc_hd__buf_6
XFILLER_42_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1407 wire1408/X vssd vssd vccd vccd wire1407/X sky130_fd_sc_hd__buf_6
XFILLER_25_2677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1418 wire1419/X vssd vssd vccd vccd wire1418/X sky130_fd_sc_hd__buf_6
Xwire1429 wire1430/X vssd vssd vccd vccd wire1429/X sky130_fd_sc_hd__buf_6
XTAP_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_170_ _170_/A _170_/B vssd vssd vccd vccd _170_/X sky130_fd_sc_hd__and2_2
XFILLER_32_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__551__B _551_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input260_A la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input358_A la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_566 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__380__A_N _508_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__279__A _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1930 wire1930/A vssd vssd vccd vccd wire1930/X sky130_fd_sc_hd__buf_6
Xwire1941 wire1942/X vssd vssd vccd vccd _602_/B sky130_fd_sc_hd__buf_6
XFILLER_4_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1952 wire1952/A vssd vssd vccd vccd wire1952/X sky130_fd_sc_hd__buf_6
XFILLER_19_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1963 wire1964/X vssd vssd vccd vccd _594_/B sky130_fd_sc_hd__buf_6
Xwire1974 wire1974/A vssd vssd vccd vccd wire1974/X sky130_fd_sc_hd__buf_6
XFILLER_20_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1985 wire1985/A vssd vssd vccd vccd wire1985/X sky130_fd_sc_hd__buf_6
XFILLER_19_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1996 wire1997/X vssd vssd vccd vccd _576_/B sky130_fd_sc_hd__buf_6
XFILLER_34_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_230 _191_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_241 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_506_ _506_/A _506_/B vssd vssd vccd vccd _506_/X sky130_fd_sc_hd__and2_4
XANTENNA_252 _521_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_263 _467_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 _380_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 wire1428/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3558 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_296 wire1781/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_437_ _565_/A _437_/B _437_/C vssd vssd vccd vccd _437_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__445__C _445_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_368_ _368_/A _368_/B vssd vssd vccd vccd _368_/X sky130_fd_sc_hd__and2_2
XFILLER_31_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output577_A _457_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_299_ _299_/A _299_/B vssd vssd vccd vccd _299_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__461__B _461_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output744_A _619_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1375_A wire1375/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] wire1325/X vssd vssd vccd vccd wire968/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_29_2098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1542_A wire1542/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__189__A _189_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1807_A wire1807/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire995_A _586_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_2470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__371__B _371_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput473 wire1057/X vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__buf_8
Xoutput484 _488_/X vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__buf_8
XFILLER_47_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput495 wire1131/X vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__buf_8
XFILLER_5_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1204 _354_/X vssd vssd vccd vccd wire1204/X sky130_fd_sc_hd__buf_6
XFILLER_9_1970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1215 wire1216/X vssd vssd vccd vccd wire1215/X sky130_fd_sc_hd__buf_6
XFILLER_9_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__099__A _099_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1226 wire1227/X vssd vssd vccd vccd wire1226/X sky130_fd_sc_hd__buf_6
XFILLER_19_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1237 _343_/X vssd vssd vccd vccd wire1237/X sky130_fd_sc_hd__buf_6
XFILLER_47_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1248 _339_/X vssd vssd vccd vccd wire1248/X sky130_fd_sc_hd__buf_6
XFILLER_47_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1259 _322_/X vssd vssd vccd vccd wire1259/X sky130_fd_sc_hd__buf_6
XFILLER_41_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__546__B _546_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4270 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_222_ _222_/A _222_/B vssd vssd vccd vccd _222_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3422 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__562__A _562_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_153_ _153_/A vssd vssd vccd vccd _153_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input71_A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_084_ _084_/A vssd vssd vccd vccd _084_/Y sky130_fd_sc_hd__inv_4
XFILLER_45_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1760 wire1760/A vssd vssd vccd vccd wire1760/X sky130_fd_sc_hd__buf_6
XFILLER_20_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1771 wire1772/X vssd vssd vccd vccd _273_/A sky130_fd_sc_hd__buf_6
XFILLER_19_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1782 wire1783/X vssd vssd vccd vccd _267_/A sky130_fd_sc_hd__buf_6
Xwire1793 wire1794/X vssd vssd vccd vccd _261_/A sky130_fd_sc_hd__buf_6
XFILLER_19_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__456__B _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1123_A _390_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output861_A _326_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[17\] mprj_dat_i_user[17] max_length1311/X vssd vssd vccd vccd
+ _131_/A sky130_fd_sc_hd__nand2_4
XANTENNA_wire1492_A wire1493/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__191__B _191_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1757_A wire1758/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1924_A wire1924/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] _278_/X vssd vssd vccd vccd wire984/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_39_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__366__B _366_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_B wire1319/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1001 _555_/X vssd vssd vccd vccd wire1001/X sky130_fd_sc_hd__buf_6
XFILLER_5_2332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1012 _546_/X vssd vssd vccd vccd wire1012/X sky130_fd_sc_hd__buf_6
Xwire1023 _531_/X vssd vssd vccd vccd wire1023/X sky130_fd_sc_hd__buf_6
XFILLER_25_2282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1034 _515_/X vssd vssd vccd vccd wire1034/X sky130_fd_sc_hd__buf_6
XFILLER_43_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1045 _505_/X vssd vssd vccd vccd wire1045/X sky130_fd_sc_hd__buf_6
XFILLER_47_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1056 _479_/X vssd vssd vccd vccd wire1056/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2140_A wire2140/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1067 _468_/X vssd vssd vccd vccd wire1067/X sky130_fd_sc_hd__buf_6
XANTENNA_input223_A la_iena_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1078 _431_/X vssd vssd vccd vccd wire1078/X sky130_fd_sc_hd__buf_6
XFILLER_38_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1089 _423_/X vssd vssd vccd vccd wire1089/X sky130_fd_sc_hd__buf_6
XANTENNA__557__A _557_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__276__B _276_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[86\]_B wire1328/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__292__A _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_205_ _205_/A _205_/B vssd vssd vccd vccd _205_/X sky130_fd_sc_hd__and2_1
XFILLER_11_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_136_ _136_/A vssd vssd vccd vccd _136_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_2540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1574 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_067_ _067_/A vssd vssd vccd vccd _067_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1073_A _462_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_4071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1590 wire1590/A vssd vssd vccd vccd _613_/A sky130_fd_sc_hd__buf_8
XFILLER_0_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__186__B _186_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1505_A wire1506/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[77\]_B _240_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1874_A wire1875/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_4225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__441__A_N _569_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input173_A la_iena_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2188_A wire2188/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input340_A la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input438_A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input34_A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__287__A _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1614 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__453__C _453_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output657_A _027_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_119_ _119_/A vssd vssd vccd vccd _119_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1190_A wire1191/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__A_N _592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output824_A wire1046/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1455_A wire1456/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] _234_/X vssd vssd vccd vccd _054_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1622_A wire1622/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__197__A _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1991_A wire1991/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_470_ _598_/A _470_/B _470_/C vssd vssd vccd vccd _470_/X sky130_fd_sc_hd__and3b_4
XTAP_2958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[125\]_B _288_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__554__B _554_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2103_A wire2104/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input290_A la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input388_A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__487__A_N _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__570__A _570_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3982 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3616 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput340 la_oenb_mprj[57] vssd vssd vccd vccd _554_/A sky130_fd_sc_hd__buf_6
XFILLER_2_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput351 la_oenb_mprj[67] vssd vssd vccd vccd wire1550/A sky130_fd_sc_hd__buf_6
Xinput362 la_oenb_mprj[77] vssd vssd vccd vccd wire1540/A sky130_fd_sc_hd__buf_6
XFILLER_3_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput373 la_oenb_mprj[87] vssd vssd vccd vccd wire1530/A sky130_fd_sc_hd__buf_6
Xinput384 la_oenb_mprj[97] vssd vssd vccd vccd _594_/A sky130_fd_sc_hd__buf_4
Xinput395 mprj_adr_o_core[16] vssd vssd vccd vccd wire1504/A sky130_fd_sc_hd__buf_6
XFILLER_53_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__448__C _448_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1036_A _513_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_599_ _599_/A _599_/B vssd vssd vccd vccd _599_/X sky130_fd_sc_hd__and2_4
XFILLER_43_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__B _464_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_B _279_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1203_A wire1204/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output774_A wire1022/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output941_A wire1235/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput803 wire997/X vssd vssd vccd vccd la_oenb_core[60] sky130_fd_sc_hd__buf_8
Xoutput814 _567_/X vssd vssd vccd vccd la_oenb_core[70] sky130_fd_sc_hd__buf_8
Xoutput825 _577_/X vssd vssd vccd vccd la_oenb_core[80] sky130_fd_sc_hd__buf_8
XFILLER_47_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput836 wire994/X vssd vssd vccd vccd la_oenb_core[90] sky130_fd_sc_hd__buf_8
Xoutput847 _146_/Y vssd vssd vccd vccd mprj_ack_i_core sky130_fd_sc_hd__buf_8
Xoutput858 wire1257/X vssd vssd vccd vccd mprj_adr_o_user[19] sky130_fd_sc_hd__buf_8
XFILLER_3_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput869 _334_/X vssd vssd vccd vccd mprj_adr_o_user[29] sky130_fd_sc_hd__buf_8
XFILLER_47_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1837_A wire1838/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[25\]_A mprj_dat_i_user[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1366 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[107\]_B wire1315/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__374__B _374_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2522 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__549__B _549_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2053_A wire2054/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input136_A la_iena_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[16\]_A mprj_dat_i_user[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_522_ _522_/A _522_/B vssd vssd vccd vccd _522_/X sky130_fd_sc_hd__and2_1
XFILLER_22_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input303_A la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__565__A _565_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_453_ _581_/A _453_/B _453_/C vssd vssd vccd vccd _453_/X sky130_fd_sc_hd__and3b_4
XTAP_2777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_384_ _512_/A _384_/B _384_/C vssd vssd vccd vccd _384_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output522_A wire1106/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__459__B _459_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1153_A _367_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput170 la_iena_mprj[19] vssd vssd vccd vccd _182_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput181 la_iena_mprj[29] vssd vssd vccd vccd _192_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_36_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput192 la_iena_mprj[39] vssd vssd vccd vccd _202_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1320_A _257_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1418_A wire1419/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] _197_/X vssd vssd vccd vccd _017_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_53_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__194__B _194_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1787_A wire1788/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1954_A wire1954/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput600 _091_/Y vssd vssd vccd vccd la_data_in_mprj[108] sky130_fd_sc_hd__buf_8
Xoutput611 _101_/Y vssd vssd vccd vccd la_data_in_mprj[118] sky130_fd_sc_hd__buf_8
Xoutput622 _159_/Y vssd vssd vccd vccd la_data_in_mprj[12] sky130_fd_sc_hd__buf_8
XFILLER_29_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput633 _005_/Y vssd vssd vccd vccd la_data_in_mprj[22] sky130_fd_sc_hd__buf_8
XFILLER_44_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput644 _015_/Y vssd vssd vccd vccd la_data_in_mprj[32] sky130_fd_sc_hd__buf_8
Xoutput655 _025_/Y vssd vssd vccd vccd la_data_in_mprj[42] sky130_fd_sc_hd__buf_8
XFILLER_9_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput666 _035_/Y vssd vssd vccd vccd la_data_in_mprj[52] sky130_fd_sc_hd__buf_8
XFILLER_29_2770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput677 _045_/Y vssd vssd vccd vccd la_data_in_mprj[62] sky130_fd_sc_hd__buf_8
Xoutput688 _055_/Y vssd vssd vccd vccd la_data_in_mprj[72] sky130_fd_sc_hd__buf_8
Xwire2109 wire2109/A vssd vssd vccd vccd wire2109/X sky130_fd_sc_hd__buf_6
XFILLER_47_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput699 _065_/Y vssd vssd vccd vccd la_data_in_mprj[82] sky130_fd_sc_hd__buf_8
Xwire1408 wire1408/A vssd vssd vccd vccd wire1408/X sky130_fd_sc_hd__buf_6
XFILLER_42_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1419 wire1420/X vssd vssd vccd vccd wire1419/X sky130_fd_sc_hd__buf_6
XFILLER_25_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__369__B _369_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2170_A wire2170/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input253_A la_iena_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input420_A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__279__B _279_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1920 wire1921/X vssd vssd vccd vccd wire1920/X sky130_fd_sc_hd__buf_6
XFILLER_19_903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1931 wire1932/X vssd vssd vccd vccd _606_/B sky130_fd_sc_hd__buf_6
XFILLER_1_3849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1942 wire1942/A vssd vssd vccd vccd wire1942/X sky130_fd_sc_hd__buf_6
Xwire1953 wire1954/X vssd vssd vccd vccd _597_/B sky130_fd_sc_hd__buf_6
XFILLER_19_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1964 wire1964/A vssd vssd vccd vccd wire1964/X sky130_fd_sc_hd__buf_6
XTAP_3220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1975 wire1975/A vssd vssd vccd vccd _587_/B sky130_fd_sc_hd__buf_6
XFILLER_19_4330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1986 wire1987/X vssd vssd vccd vccd _581_/B sky130_fd_sc_hd__buf_6
XFILLER_46_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1997 wire1997/A vssd vssd vccd vccd wire1997/X sky130_fd_sc_hd__buf_6
XFILLER_19_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_220 _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 _191_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_505_ _505_/A _505_/B vssd vssd vccd vccd _505_/X sky130_fd_sc_hd__and2_2
XTAP_2552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_242 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 _521_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_264 _466_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_275 _522_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 _319_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_436_ _564_/A _436_/B _436_/C vssd vssd vccd vccd _436_/X sky130_fd_sc_hd__and3b_4
XTAP_1862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_297 wire1790/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_367_ _367_/A _367_/B vssd vssd vccd vccd _367_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_298_ _298_/A _298_/B vssd vssd vccd vccd _298_/X sky130_fd_sc_hd__and2_2
XANTENNA_output472_A wire1058/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__461__C _461_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output737_A _613_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1270_A _316_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1368_A wire1368/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__189__B _189_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1535_A wire1535/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1702_A wire1703/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__371__C _371_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput463 wire1145/X vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__buf_8
Xoutput474 wire1135/X vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__buf_8
Xoutput485 wire1133/X vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__buf_8
Xoutput496 wire1130/X vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__buf_8
XFILLER_9_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1205 wire1206/X vssd vssd vccd vccd wire1205/X sky130_fd_sc_hd__buf_6
XFILLER_9_1960 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2475 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1216 _350_/X vssd vssd vccd vccd wire1216/X sky130_fd_sc_hd__buf_6
Xwire1227 wire1228/X vssd vssd vccd vccd wire1227/X sky130_fd_sc_hd__buf_6
XFILLER_21_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1238 wire1239/X vssd vssd vccd vccd wire1238/X sky130_fd_sc_hd__buf_6
Xwire1249 wire1250/X vssd vssd vccd vccd wire1249/X sky130_fd_sc_hd__buf_6
XFILLER_38_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2016_A wire2016/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_221_ _221_/A _221_/B vssd vssd vccd vccd _221_/X sky130_fd_sc_hd__and2_1
XFILLER_10_4146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_152_ _152_/A vssd vssd vccd vccd _152_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__562__B _562_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_083_ _083_/A vssd vssd vccd vccd _083_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_input370_A la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input64_A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_342 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1750 wire1750/A vssd vssd vccd vccd wire1750/X sky130_fd_sc_hd__buf_6
Xwire1761 wire1762/X vssd vssd vccd vccd _278_/A sky130_fd_sc_hd__buf_6
Xwire1772 wire1772/A vssd vssd vccd vccd wire1772/X sky130_fd_sc_hd__buf_6
XFILLER_18_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1783 wire1783/A vssd vssd vccd vccd wire1783/X sky130_fd_sc_hd__buf_6
XFILLER_37_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1794 wire1794/A vssd vssd vccd vccd wire1794/X sky130_fd_sc_hd__buf_6
XTAP_3050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__456__C _456_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1116_A _397_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output687_A _054_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_419_ _547_/A _419_/B _419_/C vssd vssd vccd vccd _419_/X sky130_fd_sc_hd__and3b_2
XFILLER_50_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__472__B _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output854_A wire1261/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1485_A wire1486/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1652_A wire1653/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_2615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1917_A wire1918/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] _271_/X vssd vssd vccd vccd wire990/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_17_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__370__A_N _498_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__382__B _382_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[8\]_A mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1002 wire1003/X vssd vssd vccd vccd wire1002/X sky130_fd_sc_hd__buf_6
XFILLER_40_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1013 wire1014/X vssd vssd vccd vccd wire1013/X sky130_fd_sc_hd__buf_6
XFILLER_2_3933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1024 _530_/X vssd vssd vccd vccd wire1024/X sky130_fd_sc_hd__buf_6
Xwire1035 _514_/X vssd vssd vccd vccd wire1035/X sky130_fd_sc_hd__buf_6
XFILLER_5_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1046 _504_/X vssd vssd vccd vccd wire1046/X sky130_fd_sc_hd__buf_6
XFILLER_38_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1057 _478_/X vssd vssd vccd vccd wire1057/X sky130_fd_sc_hd__buf_6
XFILLER_47_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1068 _467_/X vssd vssd vccd vccd wire1068/X sky130_fd_sc_hd__buf_6
XFILLER_0_4391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1079 _430_/X vssd vssd vccd vccd wire1079/X sky130_fd_sc_hd__buf_6
XFILLER_38_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2133_A wire2134/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input216_A la_iena_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__573__A _573_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_204_ _204_/A _204_/B vssd vssd vccd vccd _204_/X sky130_fd_sc_hd__and2_1
XFILLER_12_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__292__B _292_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_135_ _135_/A vssd vssd vccd vccd _135_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_066_ _066_/A vssd vssd vccd vccd _066_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4050 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__467__B _467_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1580 wire1580/A vssd vssd vccd vccd _623_/A sky130_fd_sc_hd__buf_6
XFILLER_21_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1591 wire1591/A vssd vssd vccd vccd _612_/A sky130_fd_sc_hd__buf_8
XANTENNA_wire1233_A wire1234/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__393__A_N _521_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1400_A wire1400/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1867_A wire1868/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__377__B _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input166_A la_iena_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2083_A wire2084/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input333_A la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__568__A _568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input27_A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__287__B _287_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1751 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_118_ _118_/A vssd vssd vccd vccd _118_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output552_A _434_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_049_ _049_/A vssd vssd vccd vccd _049_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1183_A wire1184/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output817_A _570_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1350_A wire1351/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1448_A wire1449/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] _227_/X vssd vssd vccd vccd _047_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_1_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1984_A wire1985/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire970_A wire970/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3050 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input283_A la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__570__B _570_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input450_A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput330 la_oenb_mprj[48] vssd vssd vccd vccd _417_/A_N sky130_fd_sc_hd__buf_6
XFILLER_2_4261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__298__A _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput341 la_oenb_mprj[58] vssd vssd vccd vccd wire1556/A sky130_fd_sc_hd__buf_6
XFILLER_48_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput352 la_oenb_mprj[68] vssd vssd vccd vccd wire1549/A sky130_fd_sc_hd__buf_6
Xinput363 la_oenb_mprj[78] vssd vssd vccd vccd wire1539/A sky130_fd_sc_hd__buf_6
Xinput374 la_oenb_mprj[88] vssd vssd vccd vccd wire1529/A sky130_fd_sc_hd__buf_6
XFILLER_29_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput385 la_oenb_mprj[98] vssd vssd vccd vccd wire1528/A sky130_fd_sc_hd__buf_6
XFILLER_48_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput396 mprj_adr_o_core[17] vssd vssd vccd vccd wire1500/A sky130_fd_sc_hd__buf_6
XFILLER_18_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1029_A _520_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_598_ _598_/A _598_/B vssd vssd vccd vccd _598_/X sky130_fd_sc_hd__and2_4
XFILLER_38_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__C _464_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__A_N _559_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output767_A wire1025/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1398_A wire1399/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__480__B _480_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1 la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput804 wire996/X vssd vssd vccd vccd la_oenb_core[61] sky130_fd_sc_hd__buf_8
XANTENNA_output934_A wire1154/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput815 _568_/X vssd vssd vccd vccd la_oenb_core[71] sky130_fd_sc_hd__buf_8
Xoutput826 _578_/X vssd vssd vccd vccd la_oenb_core[81] sky130_fd_sc_hd__buf_8
XFILLER_42_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput837 _588_/X vssd vssd vccd vccd la_oenb_core[91] sky130_fd_sc_hd__buf_8
XFILLER_6_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1565_A _409_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput848 _305_/X vssd vssd vccd vccd mprj_adr_o_user[0] sky130_fd_sc_hd__buf_8
XFILLER_28_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput859 _306_/X vssd vssd vccd vccd mprj_adr_o_user[1] sky130_fd_sc_hd__buf_8
XFILLER_42_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1732_A wire1733/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[25\]_B _294_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__390__B _390_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[16\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2046_A wire2046/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input129_A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1994 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_521_ _521_/A _521_/B vssd vssd vccd vccd _521_/X sky130_fd_sc_hd__and2_2
XTAP_2723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__565__B _565_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3708 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_452_ _580_/A _452_/B _452_/C vssd vssd vccd vccd _452_/X sky130_fd_sc_hd__and3b_4
XFILLER_17_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__454__A_N _582_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_383_ _511_/A _383_/B _383_/C vssd vssd vccd vccd _383_/X sky130_fd_sc_hd__and3b_4
XFILLER_25_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input94_A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__581__A _581_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__459__C _459_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output515_A wire1113/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_irq_gates\[1\]_A user_irq_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput160 la_iena_mprj[125] vssd vssd vccd vccd _288_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput171 la_iena_mprj[1] vssd vssd vccd vccd _164_/B sky130_fd_sc_hd__clkbuf_4
Xinput182 la_iena_mprj[2] vssd vssd vccd vccd _165_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput193 la_iena_mprj[3] vssd vssd vccd vccd _166_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1146_A wire1147/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__475__B _475_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1313_A _286_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] _190_/X vssd vssd vccd vccd _010_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1682_A wire1683/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput601 _092_/Y vssd vssd vccd vccd la_data_in_mprj[109] sky130_fd_sc_hd__buf_8
XFILLER_25_4037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput612 _102_/Y vssd vssd vccd vccd la_data_in_mprj[119] sky130_fd_sc_hd__buf_8
XFILLER_47_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput623 _160_/Y vssd vssd vccd vccd la_data_in_mprj[13] sky130_fd_sc_hd__buf_8
Xoutput634 _006_/Y vssd vssd vccd vccd la_data_in_mprj[23] sky130_fd_sc_hd__buf_8
Xoutput645 _016_/Y vssd vssd vccd vccd la_data_in_mprj[33] sky130_fd_sc_hd__buf_8
XFILLER_47_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput656 _026_/Y vssd vssd vccd vccd la_data_in_mprj[43] sky130_fd_sc_hd__buf_8
XFILLER_25_3336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput667 _036_/Y vssd vssd vccd vccd la_data_in_mprj[53] sky130_fd_sc_hd__buf_8
XFILLER_29_2782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput678 _046_/Y vssd vssd vccd vccd la_data_in_mprj[63] sky130_fd_sc_hd__buf_8
Xoutput689 _056_/Y vssd vssd vccd vccd la_data_in_mprj[73] sky130_fd_sc_hd__buf_8
XFILLER_42_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1409 wire1410/X vssd vssd vccd vccd _311_/B sky130_fd_sc_hd__buf_6
XFILLER_41_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__369__C _369_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__477__A_N _477_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__385__B _385_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input246_A la_iena_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2163_A wire2164/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1910 wire1910/A vssd vssd vccd vccd wire1910/X sky130_fd_sc_hd__buf_6
Xwire1921 wire1921/A vssd vssd vccd vccd wire1921/X sky130_fd_sc_hd__buf_6
XFILLER_41_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1932 wire1933/X vssd vssd vccd vccd wire1932/X sky130_fd_sc_hd__buf_6
XFILLER_46_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1943 wire1944/X vssd vssd vccd vccd _601_/B sky130_fd_sc_hd__buf_6
Xwire1954 wire1954/A vssd vssd vccd vccd wire1954/X sky130_fd_sc_hd__buf_6
XTAP_3210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1965 wire1966/X vssd vssd vccd vccd _593_/B sky130_fd_sc_hd__buf_6
XFILLER_20_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1976 wire1976/A vssd vssd vccd vccd _586_/B sky130_fd_sc_hd__buf_6
XANTENNA_input413_A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1987 wire1987/A vssd vssd vccd vccd wire1987/X sky130_fd_sc_hd__buf_6
XANTENNA__576__A _576_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1998 wire1999/X vssd vssd vccd vccd _575_/B sky130_fd_sc_hd__buf_6
XFILLER_41_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _232_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 _205_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_504_ _504_/A _504_/B vssd vssd vccd vccd _504_/X sky130_fd_sc_hd__and2_4
XANTENNA_232 _191_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__295__B _295_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_243 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 _521_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 _557_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_287 _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_435_ _563_/A _435_/B _435_/C vssd vssd vccd vccd _435_/X sky130_fd_sc_hd__and3b_4
XFILLER_37_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_298 wire1888/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_366_ _366_/A _366_/B vssd vssd vccd vccd _366_/X sky130_fd_sc_hd__and2_2
XFILLER_31_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_297_ _297_/A _297_/B vssd vssd vccd vccd _297_/X sky130_fd_sc_hd__and2_2
XFILLER_35_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output465_A wire1065/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1096_A _417_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1263_A _319_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1430_A wire1431/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1897_A wire1897/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput464 wire1066/X vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput475 wire1056/X vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__buf_8
XFILLER_9_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3166 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput486 _489_/X vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__buf_8
Xoutput497 wire1129/X vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__buf_8
XFILLER_5_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1206 wire1207/X vssd vssd vccd vccd wire1206/X sky130_fd_sc_hd__buf_6
XANTENNA_input1_A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1217 wire1218/X vssd vssd vccd vccd wire1217/X sky130_fd_sc_hd__buf_6
XFILLER_47_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1228 _346_/X vssd vssd vccd vccd wire1228/X sky130_fd_sc_hd__buf_6
XFILLER_41_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1239 wire1240/X vssd vssd vccd vccd wire1239/X sky130_fd_sc_hd__buf_6
XFILLER_28_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_220_ _220_/A _220_/B vssd vssd vccd vccd _220_/X sky130_fd_sc_hd__and2_2
XFILLER_10_4125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2009_A wire2009/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_151_ _151_/A vssd vssd vccd vccd _151_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input196_A la_iena_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_082_ _082_/A vssd vssd vccd vccd _082_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_49_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input363_A la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input57_A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4298 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1740 wire1741/X vssd vssd vccd vccd _288_/A sky130_fd_sc_hd__buf_6
XFILLER_1_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1751 wire1752/X vssd vssd vccd vccd _283_/A sky130_fd_sc_hd__buf_6
XFILLER_43_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1762 wire1762/A vssd vssd vccd vccd wire1762/X sky130_fd_sc_hd__buf_6
XFILLER_46_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1773 wire1774/X vssd vssd vccd vccd _272_/A sky130_fd_sc_hd__buf_6
XFILLER_1_2946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1784 wire1784/A vssd vssd vccd vccd _266_/A sky130_fd_sc_hd__buf_6
XTAP_3040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1795 wire1796/X vssd vssd vccd vccd _260_/A sky130_fd_sc_hd__buf_6
XTAP_3051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_266 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_418_ _546_/A _418_/B _418_/C vssd vssd vccd vccd _418_/X sky130_fd_sc_hd__and3b_4
XFILLER_42_792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1011_A wire1012/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output582_A wire1074/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1109_A _404_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_349_ _349_/A _349_/B vssd vssd vccd vccd _349_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1478_A wire1479/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] wire1320/X vssd vssd vccd vccd wire963/A
+ sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3306 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3475 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1645_A wire1645/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1812_A wire1812/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__382__C _382_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[8\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1003 _553_/X vssd vssd vccd vccd wire1003/X sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[8\]_B _171_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1014 _542_/X vssd vssd vccd vccd wire1014/X sky130_fd_sc_hd__buf_6
XFILLER_38_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1025 _525_/X vssd vssd vccd vccd wire1025/X sky130_fd_sc_hd__buf_6
XFILLER_9_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1036 _513_/X vssd vssd vccd vccd wire1036/X sky130_fd_sc_hd__buf_6
Xwire1047 _503_/X vssd vssd vccd vccd wire1047/X sky130_fd_sc_hd__buf_6
Xwire1058 _477_/X vssd vssd vccd vccd wire1058/X sky130_fd_sc_hd__buf_6
Xwire1069 _466_/X vssd vssd vccd vccd wire1069/X sky130_fd_sc_hd__buf_6
XFILLER_38_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input111_A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input209_A la_iena_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2126_A wire2127/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__573__B _573_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_203_ _203_/A _203_/B vssd vssd vccd vccd _203_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_134_ _134_/A vssd vssd vccd vccd _134_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_065_ _065_/A vssd vssd vccd vccd _065_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_49_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1059_A _476_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1570 wire1570/A vssd vssd vccd vccd _529_/A sky130_fd_sc_hd__buf_6
XFILLER_39_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1581 wire1581/A vssd vssd vccd vccd _622_/A sky130_fd_sc_hd__buf_6
Xwire1592 wire1592/A vssd vssd vccd vccd _611_/A sky130_fd_sc_hd__buf_8
XFILLER_0_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1226_A wire1227/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output797_A wire1004/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__483__B _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[22\] mprj_dat_i_user[22] max_length1310/X vssd vssd vccd vccd
+ _136_/A sky130_fd_sc_hd__nand2_4
XFILLER_50_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1762_A wire1762/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3250 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] _283_/X vssd vssd vccd vccd _103_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_6_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__377__C _377_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__393__B _393_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2076_A wire2077/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input159_A la_iena_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__568__B _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input326_A la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__584__A _584_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4066 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_117_ _117_/A vssd vssd vccd vccd _117_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_3846 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_048_ _048_/A vssd vssd vccd vccd _048_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_4_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output545_A wire1081/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1176_A wire1177/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output712_A _077_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__478__B _478_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1343_A wire1343/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2090 wire2090/A vssd vssd vccd vccd wire2090/X sky130_fd_sc_hd__buf_6
XFILLER_26_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] _220_/X vssd vssd vccd vccd _040_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1510_A wire1511/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_39_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1977_A wire1978/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__388__B _388_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1048 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2962 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1346 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2193_A wire2193/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input276_A la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__383__A_N _511_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input443_A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__579__A _579_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput320 la_oenb_mprj[39] vssd vssd vccd vccd _536_/A sky130_fd_sc_hd__clkbuf_4
Xinput331 la_oenb_mprj[49] vssd vssd vccd vccd _546_/A sky130_fd_sc_hd__buf_4
XFILLER_0_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput342 la_oenb_mprj[59] vssd vssd vccd vccd _556_/A sky130_fd_sc_hd__buf_4
XANTENNA__298__B _298_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput353 la_oenb_mprj[69] vssd vssd vccd vccd wire1548/A sky130_fd_sc_hd__buf_6
XFILLER_48_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput364 la_oenb_mprj[79] vssd vssd vccd vccd wire1538/A sky130_fd_sc_hd__buf_6
Xinput375 la_oenb_mprj[89] vssd vssd vccd vccd _586_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput386 la_oenb_mprj[99] vssd vssd vccd vccd wire1527/A sky130_fd_sc_hd__buf_6
Xinput397 mprj_adr_o_core[18] vssd vssd vccd vccd wire1497/A sky130_fd_sc_hd__buf_6
XFILLER_48_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_597_ _597_/A _597_/B vssd vssd vccd vccd _597_/X sky130_fd_sc_hd__and2_4
XFILLER_43_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output495_A wire1131/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output662_A _032_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__480__C _480_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2 la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput805 _559_/X vssd vssd vccd vccd la_oenb_core[62] sky130_fd_sc_hd__buf_8
XFILLER_47_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput816 _569_/X vssd vssd vccd vccd la_oenb_core[72] sky130_fd_sc_hd__buf_8
Xoutput827 _579_/X vssd vssd vccd vccd la_oenb_core[82] sky130_fd_sc_hd__buf_8
Xoutput838 _589_/X vssd vssd vccd vccd la_oenb_core[92] sky130_fd_sc_hd__buf_8
XFILLER_42_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output927_A wire1182/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput849 wire1271/X vssd vssd vccd vccd mprj_adr_o_user[10] sky130_fd_sc_hd__buf_8
XFILLER_6_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1460_A wire1461/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1558_A _420_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1725_A wire1725/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_520_ _520_/A _520_/B vssd vssd vccd vccd _520_/X sky130_fd_sc_hd__and2_4
XTAP_2702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2039_A wire2039/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_451_ _579_/A _451_/B _451_/C vssd vssd vccd vccd _451_/X sky130_fd_sc_hd__and3b_4
XTAP_2757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_382_ _510_/A _382_/B _382_/C vssd vssd vccd vccd _382_/X sky130_fd_sc_hd__and3b_4
XFILLER_15_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2206_A wire2207/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input393_A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__581__B _581_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input87_A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__102__A _102_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput150 la_iena_mprj[116] vssd vssd vccd vccd _279_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput161 la_iena_mprj[126] vssd vssd vccd vccd _289_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput172 la_iena_mprj[20] vssd vssd vccd vccd _183_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput183 la_iena_mprj[30] vssd vssd vccd vccd _193_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output508_A wire1119/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput194 la_iena_mprj[40] vssd vssd vccd vccd _203_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1041_A _508_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1139_A _375_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output877_A wire1277/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__491__B _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1675_A wire1675/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput602 _157_/Y vssd vssd vccd vccd la_data_in_mprj[10] sky130_fd_sc_hd__buf_8
XFILLER_9_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput613 _158_/Y vssd vssd vccd vccd la_data_in_mprj[11] sky130_fd_sc_hd__buf_8
Xoutput624 _161_/Y vssd vssd vccd vccd la_data_in_mprj[14] sky130_fd_sc_hd__buf_8
XFILLER_29_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput635 _007_/Y vssd vssd vccd vccd la_data_in_mprj[24] sky130_fd_sc_hd__buf_8
Xoutput646 _017_/Y vssd vssd vccd vccd la_data_in_mprj[34] sky130_fd_sc_hd__buf_8
Xoutput657 _027_/Y vssd vssd vccd vccd la_data_in_mprj[44] sky130_fd_sc_hd__buf_8
XANTENNA_wire1842_A wire1842/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput668 _037_/Y vssd vssd vccd vccd la_data_in_mprj[54] sky130_fd_sc_hd__buf_8
XFILLER_47_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput679 _047_/Y vssd vssd vccd vccd la_data_in_mprj[64] sky130_fd_sc_hd__buf_8
XFILLER_29_2794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1900 wire1901/X vssd vssd vccd vccd wire1900/X sky130_fd_sc_hd__buf_6
XANTENNA_input141_A la_iena_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1911 wire1912/X vssd vssd vccd vccd _612_/B sky130_fd_sc_hd__buf_6
XFILLER_3_4390 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1922 wire1923/X vssd vssd vccd vccd _609_/B sky130_fd_sc_hd__buf_6
XANTENNA_wire2156_A wire2157/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input239_A la_iena_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1933 wire1933/A vssd vssd vccd vccd wire1933/X sky130_fd_sc_hd__buf_6
XANTENNA__421__A_N _549_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1944 wire1944/A vssd vssd vccd vccd wire1944/X sky130_fd_sc_hd__buf_6
XTAP_3200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1955 wire1956/X vssd vssd vccd vccd _596_/B sky130_fd_sc_hd__buf_6
XTAP_3211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1966 wire1966/A vssd vssd vccd vccd wire1966/X sky130_fd_sc_hd__buf_6
XFILLER_19_4321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1977 wire1978/X vssd vssd vccd vccd _585_/B sky130_fd_sc_hd__buf_6
XTAP_3233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1988 wire1989/X vssd vssd vccd vccd _580_/B sky130_fd_sc_hd__buf_6
XFILLER_45_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1999 wire2000/X vssd vssd vccd vccd wire1999/X sky130_fd_sc_hd__buf_6
XANTENNA__576__B _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input406_A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_200 _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 _232_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_503_ _503_/A _503_/B vssd vssd vccd vccd _503_/X sky130_fd_sc_hd__and2_4
XANTENNA_222 _205_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_255 wire2071/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_266 mprj_dat_i_user[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_434_ _562_/A _434_/B _434_/C vssd vssd vccd vccd _434_/X sky130_fd_sc_hd__and3b_4
XANTENNA_277 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_288 _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_299 wire1904/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__592__A _592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1238 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_365_ _365_/A _365_/B vssd vssd vccd vccd _365_/X sky130_fd_sc_hd__and2_2
XFILLER_9_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_296_ _296_/A _296_/B vssd vssd vccd vccd _296_/X sky130_fd_sc_hd__and2_4
XFILLER_13_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1089_A _423_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[40\]_B _203_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1256_A _325_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__486__B _486_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1423_A wire1424/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1792_A wire1792/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1062 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__007__A _007_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] _164_/X vssd vssd vccd vccd _148_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput465 wire1065/X vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__buf_8
XFILLER_5_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[31\]_B _194_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput476 wire1055/X vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__buf_8
XFILLER_44_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__444__A_N _572_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput487 _490_/X vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__buf_8
XFILLER_9_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput498 wire1128/X vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__buf_8
XFILLER_25_3178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1207 _353_/X vssd vssd vccd vccd wire1207/X sky130_fd_sc_hd__buf_6
Xwire1218 wire1219/X vssd vssd vccd vccd wire1218/X sky130_fd_sc_hd__buf_6
XFILLER_47_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1229 wire1230/X vssd vssd vccd vccd wire1229/X sky130_fd_sc_hd__buf_6
XFILLER_9_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__396__B _396_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_B _261_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_150_ _150_/A vssd vssd vccd vccd _150_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_081_ _081_/A vssd vssd vccd vccd _081_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_12_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input189_A la_iena_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input356_A la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[22\]_B _185_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__587__A _587_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1730 wire1731/X vssd vssd vccd vccd wire1730/X sky130_fd_sc_hd__buf_6
Xwire1741 wire1741/A vssd vssd vccd vccd wire1741/X sky130_fd_sc_hd__buf_6
Xwire1752 wire1752/A vssd vssd vccd vccd wire1752/X sky130_fd_sc_hd__buf_6
Xwire1763 wire1764/X vssd vssd vccd vccd _277_/A sky130_fd_sc_hd__buf_6
XFILLER_1_2936 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1774 wire1774/A vssd vssd vccd vccd wire1774/X sky130_fd_sc_hd__buf_6
XTAP_3030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1785 wire1786/X vssd vssd vccd vccd _265_/A sky130_fd_sc_hd__buf_6
XTAP_3041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1796 wire1796/A vssd vssd vccd vccd wire1796/X sky130_fd_sc_hd__buf_6
XTAP_3052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[89\]_B wire1325/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_417_ _417_/A_N _417_/B _417_/C vssd vssd vccd vccd _417_/X sky130_fd_sc_hd__and3b_4
XTAP_1672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_348_ _348_/A _348_/B vssd vssd vccd vccd _348_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1004_A _552_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output575_A _455_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_279_ _279_/A _279_/B vssd vssd vccd vccd _279_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__467__A_N _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output742_A _617_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1373_A wire1374/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] wire1327/X vssd vssd vccd vccd wire970/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_22_3318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1540_A wire1540/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1638_A wire1638/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__497__A _497_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1004 _552_/X vssd vssd vccd vccd wire1004/X sky130_fd_sc_hd__buf_6
Xwire1015 _541_/X vssd vssd vccd vccd wire1015/X sky130_fd_sc_hd__buf_6
Xwire1026 _523_/X vssd vssd vccd vccd wire1026/X sky130_fd_sc_hd__buf_6
XFILLER_2_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1037 _512_/X vssd vssd vccd vccd wire1037/X sky130_fd_sc_hd__buf_6
XFILLER_47_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1048 _502_/X vssd vssd vccd vccd wire1048/X sky130_fd_sc_hd__buf_6
XANTENNA__200__A _200_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1059 _476_/X vssd vssd vccd vccd wire1059/X sky130_fd_sc_hd__buf_6
XFILLER_21_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input104_A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2119_A wire2120/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_202_ _202_/A _202_/B vssd vssd vccd vccd _202_/X sky130_fd_sc_hd__and2_4
XFILLER_51_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_133_ _133_/A vssd vssd vccd vccd _133_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_064_ _064_/A vssd vssd vccd vccd _064_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__110__A _110_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2650 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1560 input33/X vssd vssd vccd vccd _495_/C sky130_fd_sc_hd__buf_6
Xwire1571 _400_/A_N vssd vssd vccd vccd _528_/A sky130_fd_sc_hd__buf_6
Xwire1582 wire1582/A vssd vssd vccd vccd _621_/A sky130_fd_sc_hd__buf_6
XFILLER_19_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1593 wire1593/A vssd vssd vccd vccd _610_/A sky130_fd_sc_hd__buf_8
XFILLER_1_2788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1121_A _392_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output692_A _059_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1219_A _349_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__483__C _483_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[15\] mprj_dat_i_user[15] max_length1311/X vssd vssd vccd vccd
+ _129_/A sky130_fd_sc_hd__nand2_4
XFILLER_31_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1490_A wire1491/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1755_A wire1756/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1922_A wire1923/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2414 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__020__A _020_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1807 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] _276_/X vssd vssd vccd vccd wire986/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_6_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__393__C _393_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2069_A wire2070/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input221_A la_iena_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input319_A la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__584__B _584_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_116_ _116_/A vssd vssd vccd vccd _116_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__105__A _105_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_047_ _047_/A vssd vssd vccd vccd _047_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output538_A wire1091/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1071_A _464_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2080 wire2081/X vssd vssd vccd vccd wire2080/X sky130_fd_sc_hd__buf_6
XFILLER_43_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2091 wire2092/X vssd vssd vccd vccd _488_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1336_A input96/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1390 wire1390/A vssd vssd vccd vccd wire1390/X sky130_fd_sc_hd__buf_6
XFILLER_36_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__494__B _494_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[119\]_B _282_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1503_A wire1504/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1872_A wire1873/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[28\]_A mprj_dat_i_user[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__388__C _388_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_800 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmax_length1310 _294_/X vssd vssd vccd vccd max_length1310/X sky130_fd_sc_hd__buf_8
XFILLER_29_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input171_A la_iena_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input269_A la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2186_A wire2187/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__579__B _579_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input436_A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[19\]_A mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput310 la_oenb_mprj[2] vssd vssd vccd vccd _499_/A sky130_fd_sc_hd__buf_4
XFILLER_22_4180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput321 la_oenb_mprj[3] vssd vssd vccd vccd _500_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input32_A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput332 la_oenb_mprj[4] vssd vssd vccd vccd _501_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput343 la_oenb_mprj[5] vssd vssd vccd vccd _502_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput354 la_oenb_mprj[6] vssd vssd vccd vccd _503_/A sky130_fd_sc_hd__clkbuf_4
Xinput365 la_oenb_mprj[7] vssd vssd vccd vccd _504_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput376 la_oenb_mprj[8] vssd vssd vccd vccd _505_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput387 la_oenb_mprj[9] vssd vssd vccd vccd _506_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput398 mprj_adr_o_core[19] vssd vssd vccd vccd wire1493/A sky130_fd_sc_hd__buf_6
XANTENNA__595__A _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_596_ _596_/A _596_/B vssd vssd vccd vccd _596_/X sky130_fd_sc_hd__and2_4
XFILLER_32_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output488_A _491_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output655_A _025_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_3 la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput806 _560_/X vssd vssd vccd vccd la_oenb_core[63] sky130_fd_sc_hd__buf_8
Xoutput817 _570_/X vssd vssd vccd vccd la_oenb_core[73] sky130_fd_sc_hd__buf_8
XFILLER_6_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput828 _580_/X vssd vssd vccd vccd la_oenb_core[83] sky130_fd_sc_hd__buf_8
XFILLER_29_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1286_A wire1287/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput839 _590_/X vssd vssd vccd vccd la_oenb_core[93] sky130_fd_sc_hd__buf_8
XFILLER_42_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output822_A _575_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__489__B _489_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1453_A wire1454/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1620_A wire1620/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__399__B _399_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_450_ _578_/A _450_/B _450_/C vssd vssd vccd vccd _450_/X sky130_fd_sc_hd__and3b_4
XTAP_2747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_381_ _509_/A _381_/B _381_/C vssd vssd vccd vccd _381_/X sky130_fd_sc_hd__and3b_4
XFILLER_40_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2101_A wire2101/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input386_A la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput140 la_iena_mprj[107] vssd vssd vccd vccd _270_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput151 la_iena_mprj[117] vssd vssd vccd vccd _280_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput162 la_iena_mprj[127] vssd vssd vccd vccd _290_/B sky130_fd_sc_hd__clkbuf_4
Xinput173 la_iena_mprj[21] vssd vssd vccd vccd _184_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput184 la_iena_mprj[31] vssd vssd vccd vccd _194_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput195 la_iena_mprj[41] vssd vssd vccd vccd _204_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_4068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_579_ _579_/A _579_/B vssd vssd vccd vccd _579_/X sky130_fd_sc_hd__and2_4
XFILLER_53_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output772_A _529_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__491__C _491_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput603 _093_/Y vssd vssd vccd vccd la_data_in_mprj[110] sky130_fd_sc_hd__buf_8
Xoutput614 _103_/Y vssd vssd vccd vccd la_data_in_mprj[120] sky130_fd_sc_hd__buf_8
XANTENNA_wire1668_A wire1669/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput625 _162_/Y vssd vssd vccd vccd la_data_in_mprj[15] sky130_fd_sc_hd__buf_8
XFILLER_25_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput636 _008_/Y vssd vssd vccd vccd la_data_in_mprj[25] sky130_fd_sc_hd__buf_8
XFILLER_29_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput647 _018_/Y vssd vssd vccd vccd la_data_in_mprj[35] sky130_fd_sc_hd__buf_8
XFILLER_42_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput658 _028_/Y vssd vssd vccd vccd la_data_in_mprj[45] sky130_fd_sc_hd__buf_8
XFILLER_45_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput669 _038_/Y vssd vssd vccd vccd la_data_in_mprj[55] sky130_fd_sc_hd__buf_8
XFILLER_28_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1835_A wire1836/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4422 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__373__A_N _501_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__203__A _203_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_4459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1901 wire1901/A vssd vssd vccd vccd wire1901/X sky130_fd_sc_hd__buf_6
XFILLER_41_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1912 wire1913/X vssd vssd vccd vccd wire1912/X sky130_fd_sc_hd__buf_6
Xwire1923 wire1924/X vssd vssd vccd vccd wire1923/X sky130_fd_sc_hd__buf_6
Xwire1934 wire1935/X vssd vssd vccd vccd _605_/B sky130_fd_sc_hd__buf_6
Xwire1945 wire1946/X vssd vssd vccd vccd _600_/B sky130_fd_sc_hd__buf_6
XFILLER_19_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input134_A la_iena_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1956 wire1956/A vssd vssd vccd vccd wire1956/X sky130_fd_sc_hd__buf_6
XFILLER_18_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2051_A wire2051/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1967 wire1968/X vssd vssd vccd vccd _592_/B sky130_fd_sc_hd__buf_6
XANTENNA_wire2149_A wire2150/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1978 wire1978/A vssd vssd vccd vccd wire1978/X sky130_fd_sc_hd__buf_6
XTAP_3234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1989 wire1989/A vssd vssd vccd vccd wire1989/X sky130_fd_sc_hd__buf_6
XFILLER_18_438 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_502_ _502_/A _502_/B vssd vssd vccd vccd _502_/X sky130_fd_sc_hd__and2_4
XFILLER_19_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_212 _230_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input301_A la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_223 _205_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_245 _570_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 wire2111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_433_ _561_/A _433_/B _433_/C vssd vssd vccd vccd _433_/X sky130_fd_sc_hd__and3b_4
XTAP_1843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 wire2192/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_278 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_289 _570_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__592__B _592_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_364_ _364_/A _364_/B vssd vssd vccd vccd _364_/X sky130_fd_sc_hd__and2_2
XFILLER_35_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_295_ _295_/A_N _295_/B vssd vssd vccd vccd _295_/X sky130_fd_sc_hd__and2b_2
XFILLER_9_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output520_A wire1108/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output618_A _107_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1151_A wire1152/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1249_A wire1250/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__486__C _486_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__396__A_N _524_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1416_A wire1416/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] _195_/X vssd vssd vccd vccd _015_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_18_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1785_A wire1786/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1074 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__023__A _023_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput466 wire1064/X vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__buf_8
XFILLER_25_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput477 wire1054/X vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__buf_8
XFILLER_47_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput488 _491_/X vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__buf_8
Xoutput499 wire1127/X vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__buf_8
XFILLER_47_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1208 wire1209/X vssd vssd vccd vccd wire1208/X sky130_fd_sc_hd__buf_6
XFILLER_5_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1219 _349_/X vssd vssd vccd vccd wire1219/X sky130_fd_sc_hd__buf_6
XFILLER_45_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__396__C _396_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_080_ _080_/A vssd vssd vccd vccd _080_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_17_1294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2099_A wire2100/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input251_A la_iena_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input349_A la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1720 wire1721/X vssd vssd vccd vccd _294_/A sky130_fd_sc_hd__buf_6
XANTENNA__587__B _587_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1731 wire1731/A vssd vssd vccd vccd wire1731/X sky130_fd_sc_hd__buf_6
XFILLER_4_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1742 wire1743/X vssd vssd vccd vccd _287_/A sky130_fd_sc_hd__buf_6
Xwire1753 wire1754/X vssd vssd vccd vccd _282_/A sky130_fd_sc_hd__buf_6
Xwire1764 wire1764/A vssd vssd vccd vccd wire1764/X sky130_fd_sc_hd__buf_6
XFILLER_46_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1775 wire1776/X vssd vssd vccd vccd _271_/A sky130_fd_sc_hd__buf_6
XTAP_3031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1786 wire1786/A vssd vssd vccd vccd wire1786/X sky130_fd_sc_hd__buf_6
XFILLER_37_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1797 wire1797/A vssd vssd vccd vccd _259_/A sky130_fd_sc_hd__buf_6
XTAP_3053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_416_ _416_/A_N _416_/B _416_/C vssd vssd vccd vccd _416_/X sky130_fd_sc_hd__and3b_4
XTAP_1673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__108__A _108_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_347_ _347_/A _347_/B vssd vssd vccd vccd _347_/X sky130_fd_sc_hd__and2_4
X_278_ _278_/A _278_/B vssd vssd vccd vccd _278_/X sky130_fd_sc_hd__and2_4
XANTENNA_output470_A wire1060/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output568_A wire1138/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1199_A wire1200/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output735_A _611_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1366_A wire1366/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__497__B _497_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1533_A wire1533/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1700_A wire1701/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire986_A wire986/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__411__A_N _539_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1005 wire1006/X vssd vssd vccd vccd wire1005/X sky130_fd_sc_hd__buf_6
XFILLER_40_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1016 wire1017/X vssd vssd vccd vccd wire1016/X sky130_fd_sc_hd__buf_6
XFILLER_25_2286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1027 _522_/X vssd vssd vccd vccd wire1027/X sky130_fd_sc_hd__buf_6
Xwire1038 _511_/X vssd vssd vccd vccd wire1038/X sky130_fd_sc_hd__buf_6
Xwire1049 _501_/X vssd vssd vccd vccd wire1049/X sky130_fd_sc_hd__buf_6
XFILLER_0_4383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2014_A wire2014/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_201_ _201_/A _201_/B vssd vssd vccd vccd _201_/X sky130_fd_sc_hd__and2_4
XFILLER_11_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input299_A la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_132_ _132_/A vssd vssd vccd vccd _132_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_063_ _063_/A vssd vssd vccd vccd _063_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_3289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input62_A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__598__A _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1550 wire1550/A vssd vssd vccd vccd _564_/A sky130_fd_sc_hd__buf_6
XFILLER_19_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1561 wire1561/A vssd vssd vccd vccd _544_/A sky130_fd_sc_hd__buf_6
XFILLER_21_2662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1572 wire1572/A vssd vssd vccd vccd _527_/A sky130_fd_sc_hd__buf_8
Xwire1583 wire1583/A vssd vssd vccd vccd _620_/A sky130_fd_sc_hd__buf_6
XFILLER_19_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1594 wire1594/A vssd vssd vccd vccd _609_/A sky130_fd_sc_hd__buf_6
XFILLER_1_2756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__434__A_N _562_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output852_A wire1264/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1483_A wire1484/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1650_A wire1651/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__301__A _301_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1915_A wire1916/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] _269_/X vssd vssd vccd vccd _089_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_0_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__211__A _211_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input214_A la_iena_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__457__A_N _585_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_115_ _115_/A vssd vssd vccd vccd _115_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_046_ _046_/A vssd vssd vccd vccd _046_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__121__A _121_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1064_A _471_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2070 wire2071/X vssd vssd vccd vccd wire2070/X sky130_fd_sc_hd__buf_6
Xwire2081 wire2081/A vssd vssd vccd vccd wire2081/X sky130_fd_sc_hd__buf_6
XFILLER_36_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output600_A _091_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2092 wire2093/X vssd vssd vccd vccd wire2092/X sky130_fd_sc_hd__buf_6
XFILLER_43_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1380 wire1380/A vssd vssd vccd vccd wire1380/X sky130_fd_sc_hd__buf_6
XFILLER_19_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1391 wire1392/X vssd vssd vccd vccd _337_/B sky130_fd_sc_hd__buf_6
XANTENNA_wire1231_A _345_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1329_A _248_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__494__C _494_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1698_A wire1699/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3896 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1865_A wire1866/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[28\]_B max_length1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__206__A _206_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xmax_length1311 _294_/X vssd vssd vccd vccd max_length1311/X sky130_fd_sc_hd__buf_8
XFILLER_11_2683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2081_A wire2081/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input164_A la_iena_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2179_A wire2179/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput300 la_oenb_mprj[20] vssd vssd vccd vccd _517_/A sky130_fd_sc_hd__buf_4
XFILLER_1_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[19\]_B max_length1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput311 la_oenb_mprj[30] vssd vssd vccd vccd wire1572/A sky130_fd_sc_hd__buf_6
Xinput322 la_oenb_mprj[40] vssd vssd vccd vccd _409_/A_N sky130_fd_sc_hd__buf_6
XFILLER_22_4192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput333 la_oenb_mprj[50] vssd vssd vccd vccd _547_/A sky130_fd_sc_hd__buf_4
XANTENNA_input331_A la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput344 la_oenb_mprj[60] vssd vssd vccd vccd _557_/A sky130_fd_sc_hd__buf_4
XFILLER_29_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input429_A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput355 la_oenb_mprj[70] vssd vssd vccd vccd wire1547/A sky130_fd_sc_hd__buf_6
XFILLER_2_4297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput366 la_oenb_mprj[80] vssd vssd vccd vccd wire1537/A sky130_fd_sc_hd__buf_6
XANTENNA_input25_A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput377 la_oenb_mprj[90] vssd vssd vccd vccd _587_/A sky130_fd_sc_hd__buf_4
XFILLER_48_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput388 mprj_adr_o_core[0] vssd vssd vccd vccd wire1526/A sky130_fd_sc_hd__buf_6
Xinput399 mprj_adr_o_core[1] vssd vssd vccd vccd wire1489/A sky130_fd_sc_hd__buf_6
XFILLER_18_4217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__595__B _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_595_ _595_/A _595_/B vssd vssd vccd vccd _595_/X sky130_fd_sc_hd__and2_4
XFILLER_31_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_4 mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput807 _561_/X vssd vssd vccd vccd la_oenb_core[64] sky130_fd_sc_hd__buf_8
Xoutput818 _571_/X vssd vssd vccd vccd la_oenb_core[74] sky130_fd_sc_hd__buf_8
XFILLER_49_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output550_A _432_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput829 _581_/X vssd vssd vccd vccd la_oenb_core[84] sky130_fd_sc_hd__buf_8
XFILLER_6_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_029_ _029_/A vssd vssd vccd vccd _029_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1279_A _311_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3222 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__489__C _489_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output815_A _568_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1446_A wire1446/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] _225_/X vssd vssd vccd vccd _045_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_3_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_826 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1982_A wire1983/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__026__A _026_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__399__C _399_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_380_ _508_/A _380_/B _380_/C vssd vssd vccd vccd _380_/X sky130_fd_sc_hd__and3b_1
XFILLER_13_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_97 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input281_A la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input379_A la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_4061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput130 la_data_out_mprj[99] vssd vssd vccd vccd _468_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput141 la_iena_mprj[108] vssd vssd vccd vccd _271_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput152 la_iena_mprj[118] vssd vssd vccd vccd _281_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput163 la_iena_mprj[12] vssd vssd vccd vccd _175_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput174 la_iena_mprj[22] vssd vssd vccd vccd _185_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput185 la_iena_mprj[32] vssd vssd vccd vccd _195_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput196 la_iena_mprj[42] vssd vssd vccd vccd _205_/B sky130_fd_sc_hd__buf_4
XTAP_4673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3302 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_578_ _578_/A _578_/B vssd vssd vccd vccd _578_/X sky130_fd_sc_hd__and2_4
XFILLER_16_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output598_A _089_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output765_A wire1026/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1396_A wire1397/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output932_A wire1162/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput604 _094_/Y vssd vssd vccd vccd la_data_in_mprj[111] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput615 _104_/Y vssd vssd vccd vccd la_data_in_mprj[121] sky130_fd_sc_hd__buf_8
XFILLER_44_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput626 _163_/Y vssd vssd vccd vccd la_data_in_mprj[16] sky130_fd_sc_hd__buf_8
Xoutput637 _009_/Y vssd vssd vccd vccd la_data_in_mprj[26] sky130_fd_sc_hd__buf_8
XANTENNA_wire1563_A _415_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput648 _019_/Y vssd vssd vccd vccd la_data_in_mprj[36] sky130_fd_sc_hd__buf_8
XFILLER_28_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput659 _029_/Y vssd vssd vccd vccd la_data_in_mprj[46] sky130_fd_sc_hd__buf_8
XFILLER_42_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1730_A wire1731/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
.ends

