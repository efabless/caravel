VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM256
  CLASS BLOCK ;
  FOREIGN RAM256 ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 550.000 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 14.320 800.000 14.920 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 25.880 800.000 26.480 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 37.440 800.000 38.040 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 49.000 800.000 49.600 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 60.560 800.000 61.160 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 72.120 800.000 72.720 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 83.680 800.000 84.280 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 95.240 800.000 95.840 ;
    END
  END A0[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 349.560 800.000 350.160 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 164.600 800.000 165.200 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 280.200 800.000 280.800 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 291.760 800.000 292.360 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 303.320 800.000 303.920 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 314.880 800.000 315.480 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 326.440 800.000 327.040 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 338.000 800.000 338.600 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 361.120 800.000 361.720 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 372.680 800.000 373.280 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 384.240 800.000 384.840 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 395.800 800.000 396.400 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 176.160 800.000 176.760 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 407.360 800.000 407.960 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 418.920 800.000 419.520 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 430.480 800.000 431.080 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 442.040 800.000 442.640 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 453.600 800.000 454.200 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 465.160 800.000 465.760 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 476.720 800.000 477.320 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 488.280 800.000 488.880 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 499.840 800.000 500.440 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 511.400 800.000 512.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 187.720 800.000 188.320 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 522.960 800.000 523.560 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 534.520 800.000 535.120 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 199.280 800.000 199.880 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 210.840 800.000 211.440 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 222.400 800.000 223.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 233.960 800.000 234.560 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 245.520 800.000 246.120 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 257.080 800.000 257.680 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 268.640 800.000 269.240 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 546.000 15.090 550.000 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 546.000 263.490 550.000 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 546.000 288.330 550.000 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 546.000 313.170 550.000 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 546.000 338.010 550.000 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 546.000 362.850 550.000 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 546.000 387.690 550.000 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 546.000 412.530 550.000 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 546.000 437.370 550.000 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 546.000 462.210 550.000 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 546.000 487.050 550.000 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 546.000 39.930 550.000 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 546.000 511.890 550.000 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 546.000 536.730 550.000 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 546.000 561.570 550.000 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 546.000 586.410 550.000 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 546.000 611.250 550.000 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 546.000 636.090 550.000 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 546.000 660.930 550.000 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 546.000 685.770 550.000 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 546.000 710.610 550.000 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 546.000 735.450 550.000 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 546.000 64.770 550.000 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 546.000 760.290 550.000 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 546.000 785.130 550.000 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 546.000 89.610 550.000 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 546.000 114.450 550.000 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 546.000 139.290 550.000 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 546.000 164.130 550.000 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 546.000 188.970 550.000 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 546.000 213.810 550.000 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 546.000 238.650 550.000 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 153.040 800.000 153.640 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.920 10.640 98.520 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.520 10.640 252.120 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 10.640 405.720 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 557.720 10.640 559.320 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.320 10.640 712.920 538.800 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.120 10.640 21.720 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 173.720 10.640 175.320 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.320 10.640 328.920 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 480.920 10.640 482.520 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 634.520 10.640 636.120 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 788.120 10.640 789.720 538.800 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 106.800 800.000 107.400 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 118.360 800.000 118.960 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 129.920 800.000 130.520 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 141.480 800.000 142.080 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 4.600 10.795 795.340 538.645 ;
      LAYER met1 ;
        RECT 4.300 9.220 795.340 539.200 ;
      LAYER met2 ;
        RECT 6.080 545.720 14.530 546.450 ;
        RECT 15.370 545.720 39.370 546.450 ;
        RECT 40.210 545.720 64.210 546.450 ;
        RECT 65.050 545.720 89.050 546.450 ;
        RECT 89.890 545.720 113.890 546.450 ;
        RECT 114.730 545.720 138.730 546.450 ;
        RECT 139.570 545.720 163.570 546.450 ;
        RECT 164.410 545.720 188.410 546.450 ;
        RECT 189.250 545.720 213.250 546.450 ;
        RECT 214.090 545.720 238.090 546.450 ;
        RECT 238.930 545.720 262.930 546.450 ;
        RECT 263.770 545.720 287.770 546.450 ;
        RECT 288.610 545.720 312.610 546.450 ;
        RECT 313.450 545.720 337.450 546.450 ;
        RECT 338.290 545.720 362.290 546.450 ;
        RECT 363.130 545.720 387.130 546.450 ;
        RECT 387.970 545.720 411.970 546.450 ;
        RECT 412.810 545.720 436.810 546.450 ;
        RECT 437.650 545.720 461.650 546.450 ;
        RECT 462.490 545.720 486.490 546.450 ;
        RECT 487.330 545.720 511.330 546.450 ;
        RECT 512.170 545.720 536.170 546.450 ;
        RECT 537.010 545.720 561.010 546.450 ;
        RECT 561.850 545.720 585.850 546.450 ;
        RECT 586.690 545.720 610.690 546.450 ;
        RECT 611.530 545.720 635.530 546.450 ;
        RECT 636.370 545.720 660.370 546.450 ;
        RECT 661.210 545.720 685.210 546.450 ;
        RECT 686.050 545.720 710.050 546.450 ;
        RECT 710.890 545.720 734.890 546.450 ;
        RECT 735.730 545.720 759.730 546.450 ;
        RECT 760.570 545.720 784.570 546.450 ;
        RECT 785.410 545.720 794.320 546.450 ;
        RECT 6.080 9.190 794.320 545.720 ;
      LAYER met3 ;
        RECT 10.645 535.520 796.410 538.725 ;
        RECT 10.645 534.120 795.600 535.520 ;
        RECT 10.645 523.960 796.410 534.120 ;
        RECT 10.645 522.560 795.600 523.960 ;
        RECT 10.645 512.400 796.410 522.560 ;
        RECT 10.645 511.000 795.600 512.400 ;
        RECT 10.645 500.840 796.410 511.000 ;
        RECT 10.645 499.440 795.600 500.840 ;
        RECT 10.645 489.280 796.410 499.440 ;
        RECT 10.645 487.880 795.600 489.280 ;
        RECT 10.645 477.720 796.410 487.880 ;
        RECT 10.645 476.320 795.600 477.720 ;
        RECT 10.645 466.160 796.410 476.320 ;
        RECT 10.645 464.760 795.600 466.160 ;
        RECT 10.645 454.600 796.410 464.760 ;
        RECT 10.645 453.200 795.600 454.600 ;
        RECT 10.645 443.040 796.410 453.200 ;
        RECT 10.645 441.640 795.600 443.040 ;
        RECT 10.645 431.480 796.410 441.640 ;
        RECT 10.645 430.080 795.600 431.480 ;
        RECT 10.645 419.920 796.410 430.080 ;
        RECT 10.645 418.520 795.600 419.920 ;
        RECT 10.645 408.360 796.410 418.520 ;
        RECT 10.645 406.960 795.600 408.360 ;
        RECT 10.645 396.800 796.410 406.960 ;
        RECT 10.645 395.400 795.600 396.800 ;
        RECT 10.645 385.240 796.410 395.400 ;
        RECT 10.645 383.840 795.600 385.240 ;
        RECT 10.645 373.680 796.410 383.840 ;
        RECT 10.645 372.280 795.600 373.680 ;
        RECT 10.645 362.120 796.410 372.280 ;
        RECT 10.645 360.720 795.600 362.120 ;
        RECT 10.645 350.560 796.410 360.720 ;
        RECT 10.645 349.160 795.600 350.560 ;
        RECT 10.645 339.000 796.410 349.160 ;
        RECT 10.645 337.600 795.600 339.000 ;
        RECT 10.645 327.440 796.410 337.600 ;
        RECT 10.645 326.040 795.600 327.440 ;
        RECT 10.645 315.880 796.410 326.040 ;
        RECT 10.645 314.480 795.600 315.880 ;
        RECT 10.645 304.320 796.410 314.480 ;
        RECT 10.645 302.920 795.600 304.320 ;
        RECT 10.645 292.760 796.410 302.920 ;
        RECT 10.645 291.360 795.600 292.760 ;
        RECT 10.645 281.200 796.410 291.360 ;
        RECT 10.645 279.800 795.600 281.200 ;
        RECT 10.645 269.640 796.410 279.800 ;
        RECT 10.645 268.240 795.600 269.640 ;
        RECT 10.645 258.080 796.410 268.240 ;
        RECT 10.645 256.680 795.600 258.080 ;
        RECT 10.645 246.520 796.410 256.680 ;
        RECT 10.645 245.120 795.600 246.520 ;
        RECT 10.645 234.960 796.410 245.120 ;
        RECT 10.645 233.560 795.600 234.960 ;
        RECT 10.645 223.400 796.410 233.560 ;
        RECT 10.645 222.000 795.600 223.400 ;
        RECT 10.645 211.840 796.410 222.000 ;
        RECT 10.645 210.440 795.600 211.840 ;
        RECT 10.645 200.280 796.410 210.440 ;
        RECT 10.645 198.880 795.600 200.280 ;
        RECT 10.645 188.720 796.410 198.880 ;
        RECT 10.645 187.320 795.600 188.720 ;
        RECT 10.645 177.160 796.410 187.320 ;
        RECT 10.645 175.760 795.600 177.160 ;
        RECT 10.645 165.600 796.410 175.760 ;
        RECT 10.645 164.200 795.600 165.600 ;
        RECT 10.645 154.040 796.410 164.200 ;
        RECT 10.645 152.640 795.600 154.040 ;
        RECT 10.645 142.480 796.410 152.640 ;
        RECT 10.645 141.080 795.600 142.480 ;
        RECT 10.645 130.920 796.410 141.080 ;
        RECT 10.645 129.520 795.600 130.920 ;
        RECT 10.645 119.360 796.410 129.520 ;
        RECT 10.645 117.960 795.600 119.360 ;
        RECT 10.645 107.800 796.410 117.960 ;
        RECT 10.645 106.400 795.600 107.800 ;
        RECT 10.645 96.240 796.410 106.400 ;
        RECT 10.645 94.840 795.600 96.240 ;
        RECT 10.645 84.680 796.410 94.840 ;
        RECT 10.645 83.280 795.600 84.680 ;
        RECT 10.645 73.120 796.410 83.280 ;
        RECT 10.645 71.720 795.600 73.120 ;
        RECT 10.645 61.560 796.410 71.720 ;
        RECT 10.645 60.160 795.600 61.560 ;
        RECT 10.645 50.000 796.410 60.160 ;
        RECT 10.645 48.600 795.600 50.000 ;
        RECT 10.645 38.440 796.410 48.600 ;
        RECT 10.645 37.040 795.600 38.440 ;
        RECT 10.645 26.880 796.410 37.040 ;
        RECT 10.645 25.480 795.600 26.880 ;
        RECT 10.645 15.320 796.410 25.480 ;
        RECT 10.645 13.920 795.600 15.320 ;
        RECT 10.645 10.715 796.410 13.920 ;
      LAYER met4 ;
        RECT 15.935 28.735 19.720 527.505 ;
        RECT 22.120 28.735 96.520 527.505 ;
        RECT 98.920 28.735 173.320 527.505 ;
        RECT 175.720 28.735 250.120 527.505 ;
        RECT 252.520 28.735 326.920 527.505 ;
        RECT 329.320 28.735 403.720 527.505 ;
        RECT 406.120 28.735 480.520 527.505 ;
        RECT 482.920 28.735 557.320 527.505 ;
        RECT 559.720 28.735 634.120 527.505 ;
        RECT 636.520 28.735 710.920 527.505 ;
        RECT 713.320 28.735 779.865 527.505 ;
  END
END RAM256
END LIBRARY

