* NGSPICE file created from digital_pll.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_2 abstract view
.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_8 abstract view
.subckt sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_4 abstract view
.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_1 abstract view
.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

.subckt digital_pll VGND VPWR clockp[0] clockp[1] dco div[0] div[1] div[2] div[3]
+ div[4] enable ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14]
+ ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20]
+ ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3]
+ ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_363_ _348_/X ext_trim[2] _398_/B _362_/Y VGND VGND VPWR VPWR _363_/X sky130_fd_sc_hd__a211o_2
X_432_ _437_/A _433_/B VGND VGND VPWR VPWR _432_/Y sky130_fd_sc_hd__nor2_2
X_294_ _397_/A _325_/A VGND VGND VPWR VPWR _313_/A sky130_fd_sc_hd__xnor2_2
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_346_ _346_/A VGND VGND VPWR VPWR _456_/D sky130_fd_sc_hd__buf_2
X_415_ _376_/A _370_/A _468_/Q VGND VGND VPWR VPWR _416_/B sky130_fd_sc_hd__o21ai_2
X_277_ _420_/B _302_/A VGND VGND VPWR VPWR _278_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_329_ _463_/Q _291_/X _328_/Y VGND VGND VPWR VPWR _463_/D sky130_fd_sc_hd__o21a_2
Xringosc.dstage\[11\].id.delayen1 ringosc.dstage\[11\].id.delayen1/A _423_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XANTENNA__392__A2 ext_trim[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__383__A2 ext_trim[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[10\].id.delayenb0 ringosc.dstage\[10\].id.delayenb1/A _385_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[9\].id.delayenb0 ringosc.dstage\[9\].id.delayenb1/A _383_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_431_ _437_/A _433_/B VGND VGND VPWR VPWR _431_/Y sky130_fd_sc_hd__nor2_2
X_293_ _293_/A VGND VGND VPWR VPWR _328_/B sky130_fd_sc_hd__buf_2
X_362_ _397_/A _438_/A VGND VGND VPWR VPWR _362_/Y sky130_fd_sc_hd__nor2_2
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_414_ _406_/B _359_/A _371_/Y _403_/B _413_/X VGND VGND VPWR VPWR _414_/X sky130_fd_sc_hd__o2111a_2
X_345_ _455_/Q _456_/Q _345_/S VGND VGND VPWR VPWR _346_/A sky130_fd_sc_hd__mux2_2
X_276_ _465_/Q VGND VGND VPWR VPWR _302_/A sky130_fd_sc_hd__inv_2
X_259_ _288_/B _288_/C _258_/X VGND VGND VPWR VPWR _259_/X sky130_fd_sc_hd__a21o_2
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_328_ _463_/Q _328_/B VGND VGND VPWR VPWR _328_/Y sky130_fd_sc_hd__nand2_2
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[9\].id.delayenb1 ringosc.dstage\[9\].id.delayenb1/A _421_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[10\].id.delayenb1 ringosc.dstage\[10\].id.delayenb1/A _422_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_361_ _367_/A dco VGND VGND VPWR VPWR _398_/B sky130_fd_sc_hd__nor2_2
X_430_ _437_/A _433_/B VGND VGND VPWR VPWR _430_/Y sky130_fd_sc_hd__nor2_2
X_292_ _397_/A _325_/A _278_/Y _291_/X VGND VGND VPWR VPWR _293_/A sky130_fd_sc_hd__o31a_2
X_275_ _466_/Q VGND VGND VPWR VPWR _420_/B sky130_fd_sc_hd__inv_2
X_413_ _301_/Y _367_/Y _386_/Y _412_/X VGND VGND VPWR VPWR _413_/X sky130_fd_sc_hd__o211a_2
X_344_ _344_/A VGND VGND VPWR VPWR _457_/D sky130_fd_sc_hd__buf_2
XANTENNA__410__A2 ext_trim[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[4\].id.delayen0 ringosc.dstage\[4\].id.delayen0/A _369_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_258_ div[1] _258_/B VGND VGND VPWR VPWR _258_/X sky130_fd_sc_hd__and2_2
X_327_ _327_/A VGND VGND VPWR VPWR _464_/D sky130_fd_sc_hd__buf_2
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[8\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[5\].id.delayenb0 ringosc.dstage\[5\].id.delayenb1/A _373_/X VGND
+ VGND VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvn_8
X_360_ _352_/X ext_trim[1] _403_/A VGND VGND VPWR VPWR _360_/X sky130_fd_sc_hd__a21o_2
X_291_ _285_/X _291_/B _291_/C VGND VGND VPWR VPWR _291_/X sky130_fd_sc_hd__and3b_2
XANTENNA__244__A div[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_412_ _420_/B _283_/B _381_/A _376_/Y VGND VGND VPWR VPWR _412_/X sky130_fd_sc_hd__o22a_2
X_343_ _456_/Q _457_/Q _345_/S VGND VGND VPWR VPWR _344_/A sky130_fd_sc_hd__mux2_2
X_274_ _464_/Q _463_/Q VGND VGND VPWR VPWR _324_/B sky130_fd_sc_hd__and2_2
Xringosc.dstage\[4\].id.delayen1 ringosc.dstage\[4\].id.delayen1/A _409_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_257_ div[0] _257_/B _257_/C VGND VGND VPWR VPWR _288_/C sky130_fd_sc_hd__nand3b_2
X_326_ _464_/Q _325_/X _328_/B VGND VGND VPWR VPWR _327_/A sky130_fd_sc_hd__mux2_2
XANTENNA__252__A div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_309_ _309_/A _309_/B VGND VGND VPWR VPWR _309_/X sky130_fd_sc_hd__and2_2
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[5\].id.delayenb1 ringosc.dstage\[5\].id.delayenb1/A _410_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__350__A ext_trim[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_290_ _266_/X _290_/B _290_/C _290_/D VGND VGND VPWR VPWR _291_/C sky130_fd_sc_hd__nand4b_2
X_411_ _379_/X ext_trim[19] _403_/A _403_/B VGND VGND VPWR VPWR _411_/X sky130_fd_sc_hd__a22o_2
X_342_ _342_/A _347_/B _342_/C VGND VGND VPWR VPWR _458_/D sky130_fd_sc_hd__nand3_2
XFILLER_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_273_ _467_/Q VGND VGND VPWR VPWR _376_/A sky130_fd_sc_hd__buf_2
XFILLER_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_256_ _256_/A VGND VGND VPWR VPWR _257_/C sky130_fd_sc_hd__inv_2
X_325_ _325_/A _325_/B VGND VGND VPWR VPWR _325_/X sky130_fd_sc_hd__xor2_2
X_239_ _262_/A _239_/B VGND VGND VPWR VPWR _240_/C sky130_fd_sc_hd__nand2b_2
X_308_ _420_/A _325_/A VGND VGND VPWR VPWR _309_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__348__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__258__A div[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__422__A2 ext_trim[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[4\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__404__A2 ext_trim[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_410_ _428_/A ext_trim[18] _398_/X VGND VGND VPWR VPWR _410_/X sky130_fd_sc_hd__a21o_2
Xringosc.dstage\[1\].id.delayenb0 ringosc.dstage\[1\].id.delayenb1/A _360_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_341_ _342_/C _340_/Y _347_/B VGND VGND VPWR VPWR _459_/D sky130_fd_sc_hd__a21boi_2
XFILLER_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_272_ _302_/B VGND VGND VPWR VPWR _325_/A sky130_fd_sc_hd__buf_2
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_255_ _342_/A _473_/Q VGND VGND VPWR VPWR _256_/A sky130_fd_sc_hd__nor2_2
X_324_ _324_/A _324_/B VGND VGND VPWR VPWR _325_/B sky130_fd_sc_hd__nor2_2
XANTENNA__266__A div[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_238_ _461_/Q _476_/Q VGND VGND VPWR VPWR _239_/B sky130_fd_sc_hd__nand2_2
X_307_ _313_/A _316_/A _316_/B _398_/A _325_/A VGND VGND VPWR VPWR _309_/A sky130_fd_sc_hd__a32o_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[5\].id.delaybuf1 ringosc.dstage\[5\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[1\].id.delayenb1 ringosc.dstage\[1\].id.delayenb1/A _396_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XANTENNA__361__B dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_340_ _459_/Q _342_/A VGND VGND VPWR VPWR _340_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_271_ _260_/X _266_/X _267_/X _290_/C VGND VGND VPWR VPWR _302_/B sky130_fd_sc_hd__o31a_2
Xringosc.dstage\[1\].id.delayen0 ringosc.dstage\[1\].id.delayen0/A _360_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_469_ _477_/CLK _469_/D _445_/Y VGND VGND VPWR VPWR _469_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__389__A2 ext_trim[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_254_ _342_/A _473_/Q VGND VGND VPWR VPWR _257_/B sky130_fd_sc_hd__nand2_2
X_323_ _328_/B _322_/Y _465_/Q _291_/X VGND VGND VPWR VPWR _465_/D sky130_fd_sc_hd__o2bb2a_2
X_237_ _461_/Q _476_/Q VGND VGND VPWR VPWR _262_/A sky130_fd_sc_hd__nor2_2
X_306_ _401_/B VGND VGND VPWR VPWR _398_/A sky130_fd_sc_hd__inv_2
XANTENNA__289__A1 div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_270_ div[4] _266_/B _268_/Y _269_/Y VGND VGND VPWR VPWR _290_/C sky130_fd_sc_hd__o211a_2
X_399_ _379_/X ext_trim[15] _397_/Y _398_/X VGND VGND VPWR VPWR _399_/X sky130_fd_sc_hd__a22o_2
Xringosc.dstage\[1\].id.delayen1 ringosc.dstage\[1\].id.delayen1/A _396_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_468_ _477_/CLK _468_/D _444_/Y VGND VGND VPWR VPWR _468_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[0\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_322_ _322_/A _322_/B VGND VGND VPWR VPWR _322_/Y sky130_fd_sc_hd__xnor2_2
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_253_ _258_/B _253_/B VGND VGND VPWR VPWR _288_/B sky130_fd_sc_hd__nand2b_2
X_236_ _251_/A _251_/B _247_/B _235_/X VGND VGND VPWR VPWR _240_/B sky130_fd_sc_hd__a211o_2
X_305_ _301_/Y _322_/A _322_/B _406_/C _325_/A VGND VGND VPWR VPWR _316_/B sky130_fd_sc_hd__a32o_2
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ _461_/Q _476_/Q _345_/S VGND VGND VPWR VPWR _220_/A sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[9\].id.delayen0 ringosc.dstage\[9\].id.delayen0/A _383_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_467_ _477_/CLK _467_/D _442_/Y VGND VGND VPWR VPWR _467_/Q sky130_fd_sc_hd__dfrtp_2
X_398_ _398_/A _398_/B VGND VGND VPWR VPWR _398_/X sky130_fd_sc_hd__and2_2
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_252_ div[1] VGND VGND VPWR VPWR _253_/B sky130_fd_sc_hd__inv_2
X_321_ _420_/B _321_/B VGND VGND VPWR VPWR _466_/D sky130_fd_sc_hd__xnor2_2
X_235_ _459_/Q _474_/Q VGND VGND VPWR VPWR _235_/X sky130_fd_sc_hd__and2_2
X_304_ _302_/B _303_/Y _324_/B VGND VGND VPWR VPWR _322_/B sky130_fd_sc_hd__a21o_2
X_218_ _218_/A VGND VGND VPWR VPWR _477_/D sky130_fd_sc_hd__buf_2
Xringosc.dstage\[9\].id.delayen1 ringosc.dstage\[9\].id.delayen1/A _421_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__270__A1 div[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_397_ _397_/A _397_/B VGND VGND VPWR VPWR _397_/Y sky130_fd_sc_hd__nand2_2
X_466_ _477_/CLK _466_/D _441_/Y VGND VGND VPWR VPWR _466_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_251_ _251_/A _251_/B VGND VGND VPWR VPWR _258_/B sky130_fd_sc_hd__xnor2_2
X_320_ _302_/A _322_/B _319_/X _293_/A VGND VGND VPWR VPWR _321_/B sky130_fd_sc_hd__o211a_2
X_449_ _454_/A _451_/B VGND VGND VPWR VPWR _449_/Y sky130_fd_sc_hd__nor2_2
X_234_ _460_/Q _475_/Q VGND VGND VPWR VPWR _247_/B sky130_fd_sc_hd__and2_2
X_303_ _324_/A VGND VGND VPWR VPWR _303_/Y sky130_fd_sc_hd__inv_2
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.iss.reseten0 ringosc.iss.const1/HI _433_/B VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_1
XANTENNA__470__D osc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_217_ _462_/Q _477_/Q _347_/B VGND VGND VPWR VPWR _218_/A sky130_fd_sc_hd__mux2_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_396_ _379_/X ext_trim[14] _372_/X _395_/X VGND VGND VPWR VPWR _396_/X sky130_fd_sc_hd__a22o_2
Xringosc.dstage\[8\].id.delayenb0 ringosc.dstage\[8\].id.delayenb1/A _380_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_465_ _477_/CLK _465_/D _440_/Y VGND VGND VPWR VPWR _465_/Q sky130_fd_sc_hd__dfrtp_2
X_250_ _250_/A _250_/B VGND VGND VPWR VPWR _250_/Y sky130_fd_sc_hd__nand2_2
X_448_ _454_/A _451_/B VGND VGND VPWR VPWR _448_/Y sky130_fd_sc_hd__nor2_2
X_379_ dco VGND VGND VPWR VPWR _379_/X sky130_fd_sc_hd__buf_2
X_233_ _459_/Q _474_/Q VGND VGND VPWR VPWR _251_/B sky130_fd_sc_hd__xor2_2
X_302_ _302_/A _302_/B VGND VGND VPWR VPWR _322_/A sky130_fd_sc_hd__xnor2_2
X_216_ _345_/S VGND VGND VPWR VPWR _347_/B sky130_fd_sc_hd__buf_2
Xringosc.iss.delayint0 ringosc.iss.delayen1/Z VGND VGND VPWR VPWR ringosc.iss.delayen0/A
+ sky130_fd_sc_hd__clkinv_1
XANTENNA__419__A2 ext_trim[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_464_ _477_/CLK _464_/D _439_/Y VGND VGND VPWR VPWR _464_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[8\].id.delayenb1 ringosc.dstage\[8\].id.delayenb1/A _419_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XFILLER_4_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_395_ _376_/B _395_/B _395_/C VGND VGND VPWR VPWR _395_/X sky130_fd_sc_hd__and3b_2
X_378_ _352_/X ext_trim[7] _377_/X VGND VGND VPWR VPWR _378_/X sky130_fd_sc_hd__a21o_2
X_447_ dco VGND VGND VPWR VPWR _454_/A sky130_fd_sc_hd__buf_2
X_301_ _406_/C _381_/A VGND VGND VPWR VPWR _301_/Y sky130_fd_sc_hd__nand2_2
X_232_ _458_/Q _473_/Q VGND VGND VPWR VPWR _251_/A sky130_fd_sc_hd__and2_2
Xringosc.dstage\[6\].id.delayen0 ringosc.dstage\[6\].id.delayen0/A _375_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_215_ _215_/A VGND VGND VPWR VPWR _345_/S sky130_fd_sc_hd__buf_2
XANTENNA__373__A2 ext_trim[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__364__A2 ext_trim[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_463_ _477_/CLK _463_/D _437_/Y VGND VGND VPWR VPWR _463_/Q sky130_fd_sc_hd__dfrtp_2
X_394_ _420_/A _278_/D _420_/C VGND VGND VPWR VPWR _395_/C sky130_fd_sc_hd__o21ai_2
X_377_ _406_/C _376_/Y _403_/A VGND VGND VPWR VPWR _377_/X sky130_fd_sc_hd__o21a_2
X_446_ _446_/A _451_/B VGND VGND VPWR VPWR _446_/Y sky130_fd_sc_hd__nor2_2
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[7\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[4\].id.delayenb0 ringosc.dstage\[4\].id.delayenb1/A _369_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_231_ _460_/Q _231_/B VGND VGND VPWR VPWR _240_/A sky130_fd_sc_hd__nand2b_2
X_300_ _370_/A _465_/Q VGND VGND VPWR VPWR _381_/A sky130_fd_sc_hd__nand2_2
X_429_ _438_/A VGND VGND VPWR VPWR _437_/A sky130_fd_sc_hd__buf_2
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[10\].id.delayen0 ringosc.dstage\[10\].id.delayen0/A _385_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[6\].id.delayen1 ringosc.dstage\[6\].id.delayen1/A _411_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_214_ _472_/D _472_/Q VGND VGND VPWR VPWR _215_/A sky130_fd_sc_hd__xnor2_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_462_ _477_/CLK _462_/D _436_/Y VGND VGND VPWR VPWR _462_/Q sky130_fd_sc_hd__dfrtp_2
X_393_ _468_/Q _406_/C _376_/A _367_/A VGND VGND VPWR VPWR _395_/B sky130_fd_sc_hd__a211o_2
XFILLER_1_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_376_ _376_/A _376_/B VGND VGND VPWR VPWR _376_/Y sky130_fd_sc_hd__nand2_2
X_445_ _446_/A _451_/B VGND VGND VPWR VPWR _445_/Y sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[4\].id.delayenb1 ringosc.dstage\[4\].id.delayenb1/A _409_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_230_ _475_/Q VGND VGND VPWR VPWR _231_/B sky130_fd_sc_hd__inv_2
X_359_ _359_/A _359_/B VGND VGND VPWR VPWR _403_/A sky130_fd_sc_hd__and2_2
X_428_ _428_/A _433_/B VGND VGND VPWR VPWR _428_/Y sky130_fd_sc_hd__nor2_2
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[10\].id.delayen1 ringosc.dstage\[10\].id.delayen1/A _422_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__421__B1 ext_trim[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_392_ _428_/A ext_trim[13] _391_/X VGND VGND VPWR VPWR _392_/X sky130_fd_sc_hd__a21o_2
X_461_ _477_/CLK _461_/D _435_/Y VGND VGND VPWR VPWR _461_/Q sky130_fd_sc_hd__dfrtp_2
X_375_ _352_/X ext_trim[6] _374_/Y VGND VGND VPWR VPWR _375_/X sky130_fd_sc_hd__a21o_2
X_444_ _446_/A _451_/B VGND VGND VPWR VPWR _444_/Y sky130_fd_sc_hd__nor2_2
X_427_ _428_/A _433_/B VGND VGND VPWR VPWR _427_/Y sky130_fd_sc_hd__nor2_2
X_358_ dco _358_/B VGND VGND VPWR VPWR _359_/B sky130_fd_sc_hd__nor2_2
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[3\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_289_ div[3] _242_/Y _249_/X _250_/Y VGND VGND VPWR VPWR _290_/D sky130_fd_sc_hd__o211a_2
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[0\].id.delayenb0 ringosc.dstage\[0\].id.delayenb1/A _351_/Y VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__267__A1 div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__425__A enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_391_ _370_/A _376_/Y _403_/A VGND VGND VPWR VPWR _391_/X sky130_fd_sc_hd__o21a_2
X_460_ _477_/CLK _460_/D _433_/Y VGND VGND VPWR VPWR _460_/Q sky130_fd_sc_hd__dfrtp_2
X_374_ _420_/B _358_/B dco VGND VGND VPWR VPWR _374_/Y sky130_fd_sc_hd__a21oi_2
X_443_ _454_/B VGND VGND VPWR VPWR _451_/B sky130_fd_sc_hd__buf_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[3\].id.delayen0 ringosc.dstage\[3\].id.delayen0/A _364_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ _469_/Q _398_/A VGND VGND VPWR VPWR _358_/B sky130_fd_sc_hd__nor2_2
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_426_ _454_/B VGND VGND VPWR VPWR _433_/B sky130_fd_sc_hd__buf_2
X_288_ _258_/X _288_/B _288_/C _288_/D VGND VGND VPWR VPWR _290_/B sky130_fd_sc_hd__and4b_2
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[0\].id.delayenb1 ringosc.dstage\[0\].id.delayenb1/A _392_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_409_ _405_/Y _407_/X _408_/X ext_trim[17] _348_/X VGND VGND VPWR VPWR _409_/X sky130_fd_sc_hd__a32o_2
XFILLER_21_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.iss.delayenb0 ringosc.iss.delayenb1/A ringosc.iss.ctrlen0/X VGND VGND VPWR
+ VPWR ringosc.ibufp00/A sky130_fd_sc_hd__einvn_8
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__425__B resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_390_ _438_/A VGND VGND VPWR VPWR _428_/A sky130_fd_sc_hd__buf_2
XFILLER_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_373_ _352_/X ext_trim[5] _372_/X VGND VGND VPWR VPWR _373_/X sky130_fd_sc_hd__a21o_2
X_442_ _446_/A _442_/B VGND VGND VPWR VPWR _442_/Y sky130_fd_sc_hd__nor2_2
X_356_ _386_/B _371_/B VGND VGND VPWR VPWR _359_/A sky130_fd_sc_hd__nor2_2
X_287_ _251_/A _256_/A div[0] VGND VGND VPWR VPWR _288_/D sky130_fd_sc_hd__o21ai_2
X_425_ enable resetb VGND VGND VPWR VPWR _454_/B sky130_fd_sc_hd__nand2_2
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[3\].id.delayen1 ringosc.dstage\[3\].id.delayen1/A _404_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ _420_/B _365_/Y _401_/Y _406_/B _403_/B VGND VGND VPWR VPWR _408_/X sky130_fd_sc_hd__o221a_2
X_339_ _339_/A VGND VGND VPWR VPWR _460_/D sky130_fd_sc_hd__buf_2
Xringosc.iss.delayenb1 ringosc.iss.delayenb1/A _424_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.dstage\[0\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XANTENNA__349__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_372_ _301_/Y _367_/Y _359_/B _371_/Y VGND VGND VPWR VPWR _372_/X sky130_fd_sc_hd__o211a_2
X_441_ _446_/A _442_/B VGND VGND VPWR VPWR _441_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__447__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_355_ _367_/A _397_/A _467_/Q VGND VGND VPWR VPWR _371_/B sky130_fd_sc_hd__and3_2
X_286_ _215_/A _455_/Q _457_/Q _456_/Q VGND VGND VPWR VPWR _291_/B sky130_fd_sc_hd__and4b_2
X_424_ _379_/X ext_trim[25] _403_/X _407_/C VGND VGND VPWR VPWR _424_/X sky130_fd_sc_hd__a22o_2
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ _407_/A _407_/B _407_/C VGND VGND VPWR VPWR _407_/X sky130_fd_sc_hd__and3_2
X_338_ _347_/B _338_/B VGND VGND VPWR VPWR _339_/A sky130_fd_sc_hd__and2_2
X_269_ _462_/Q _477_/Q VGND VGND VPWR VPWR _269_/Y sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/A VGND VGND VPWR VPWR ringosc.iss.delayen1/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_371_ _397_/B _371_/B VGND VGND VPWR VPWR _371_/Y sky130_fd_sc_hd__nand2_2
X_440_ _446_/A _442_/B VGND VGND VPWR VPWR _440_/Y sky130_fd_sc_hd__nor2_2
X_354_ _467_/Q _376_/B VGND VGND VPWR VPWR _386_/B sky130_fd_sc_hd__and2b_2
X_285_ _302_/B _285_/B _324_/A VGND VGND VPWR VPWR _285_/X sky130_fd_sc_hd__and3_2
X_423_ _379_/X ext_trim[24] _362_/Y _420_/A VGND VGND VPWR VPWR _423_/X sky130_fd_sc_hd__a22o_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_406_ _401_/Y _406_/B _406_/C VGND VGND VPWR VPWR _407_/C sky130_fd_sc_hd__nand3b_2
X_337_ _331_/B _335_/Y _342_/C VGND VGND VPWR VPWR _338_/B sky130_fd_sc_hd__o21ai_2
X_268_ _268_/A _268_/B VGND VGND VPWR VPWR _268_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__424__A2 ext_trim[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_370_ _370_/A _465_/Q VGND VGND VPWR VPWR _397_/B sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[0\].id.delayen0 ringosc.dstage\[0\].id.delayen0/A _351_/Y VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
X_422_ _428_/A ext_trim[23] _398_/B VGND VGND VPWR VPWR _422_/X sky130_fd_sc_hd__a21o_2
X_284_ _464_/Q _463_/Q VGND VGND VPWR VPWR _324_/A sky130_fd_sc_hd__nor2_2
X_353_ _469_/Q _397_/A VGND VGND VPWR VPWR _376_/B sky130_fd_sc_hd__nor2_2
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[7\].id.delayenb0 ringosc.dstage\[7\].id.delayenb1/A _378_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
X_405_ _420_/A _406_/B _420_/C VGND VGND VPWR VPWR _405_/Y sky130_fd_sc_hd__nand3_2
X_336_ _462_/Q _336_/B VGND VGND VPWR VPWR _342_/C sky130_fd_sc_hd__nand2_2
X_267_ div[3] _242_/Y _249_/X VGND VGND VPWR VPWR _267_/X sky130_fd_sc_hd__o21ba_2
XANTENNA__379__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__409__B1 ext_trim[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__360__A2 ext_trim[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_319_ _465_/Q _324_/A _325_/A VGND VGND VPWR VPWR _319_/X sky130_fd_sc_hd__mux2_2
XANTENNA__260__A1 div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_421_ _407_/X _408_/X _420_/Y ext_trim[22] _348_/X VGND VGND VPWR VPWR _421_/X sky130_fd_sc_hd__a32o_2
Xringosc.dstage\[0\].id.delayen1 ringosc.dstage\[0\].id.delayen1/A _392_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _438_/A VGND VGND VPWR VPWR _352_/X sky130_fd_sc_hd__buf_2
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _298_/A _283_/B VGND VGND VPWR VPWR _285_/B sky130_fd_sc_hd__nor2_2
X_404_ _428_/A ext_trim[16] _403_/X VGND VGND VPWR VPWR _404_/X sky130_fd_sc_hd__a21o_2
Xringosc.dstage\[7\].id.delayenb1 ringosc.dstage\[7\].id.delayenb1/A _417_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
X_335_ _459_/Q _342_/A _460_/Q VGND VGND VPWR VPWR _335_/Y sky130_fd_sc_hd__a21oi_2
X_266_ div[4] _266_/B VGND VGND VPWR VPWR _266_/X sky130_fd_sc_hd__and2_2
X_318_ _318_/A VGND VGND VPWR VPWR _467_/D sky130_fd_sc_hd__buf_2
X_249_ _243_/Y _242_/A _242_/B _250_/A _250_/B VGND VGND VPWR VPWR _249_/X sky130_fd_sc_hd__o32a_2
Xringosc.dstage\[8\].id.delayen0 ringosc.dstage\[8\].id.delayen0/A _380_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
Xclockp_buffer_0 _477_/CLK VGND VGND VPWR VPWR clockp[0] sky130_fd_sc_hd__clkbuf_16
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_420_ _420_/A _420_/B _420_/C VGND VGND VPWR VPWR _420_/Y sky130_fd_sc_hd__nand3_2
X_351_ _348_/X _285_/B _350_/Y VGND VGND VPWR VPWR _351_/Y sky130_fd_sc_hd__o21ai_2
X_282_ _367_/A _401_/B VGND VGND VPWR VPWR _283_/B sky130_fd_sc_hd__nand2_2
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _403_/A _403_/B _407_/B VGND VGND VPWR VPWR _403_/X sky130_fd_sc_hd__and3_2
X_334_ _461_/Q _331_/B _333_/Y _347_/B VGND VGND VPWR VPWR _461_/D sky130_fd_sc_hd__o211a_2
XFILLER_2_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_265_ _268_/A _268_/B VGND VGND VPWR VPWR _266_/B sky130_fd_sc_hd__xnor2_2
X_248_ _248_/A _248_/B VGND VGND VPWR VPWR _250_/B sky130_fd_sc_hd__xnor2_2
X_317_ _376_/A _316_/X _328_/B VGND VGND VPWR VPWR _318_/A sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[6\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[3\].id.delayenb0 ringosc.dstage\[3\].id.delayenb1/A _364_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[8\].id.delayen1 ringosc.dstage\[8\].id.delayen1/A _419_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
Xclockp_buffer_1 ringosc.ibufp11/Y VGND VGND VPWR VPWR clockp[1] sky130_fd_sc_hd__clkbuf_16
XANTENNA__384__A_N ext_trim[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_350_ ext_trim[0] _438_/A VGND VGND VPWR VPWR _350_/Y sky130_fd_sc_hd__nand2_2
X_281_ _468_/Q _467_/Q VGND VGND VPWR VPWR _401_/B sky130_fd_sc_hd__nor2_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__257__A_N div[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_402_ _381_/A _376_/Y _401_/Y _406_/C VGND VGND VPWR VPWR _407_/B sky130_fd_sc_hd__o22a_2
X_333_ _462_/Q _336_/B VGND VGND VPWR VPWR _333_/Y sky130_fd_sc_hd__nand2b_2
X_264_ _262_/Y _240_/A _240_/B _263_/X VGND VGND VPWR VPWR _268_/B sky130_fd_sc_hd__a31o_2
XANTENNA__363__A2 ext_trim[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_247_ _247_/A _247_/B VGND VGND VPWR VPWR _248_/B sky130_fd_sc_hd__nor2_2
X_316_ _316_/A _316_/B VGND VGND VPWR VPWR _316_/X sky130_fd_sc_hd__xor2_2
Xringosc.dstage\[3\].id.delayenb1 ringosc.dstage\[3\].id.delayenb1/A _404_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ _469_/Q VGND VGND VPWR VPWR _367_/A sky130_fd_sc_hd__inv_2
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ _462_/Q _336_/B _347_/B VGND VGND VPWR VPWR _462_/D sky130_fd_sc_hd__o21a_2
X_263_ _461_/Q _476_/Q VGND VGND VPWR VPWR _263_/X sky130_fd_sc_hd__and2_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_401_ _469_/Q _401_/B VGND VGND VPWR VPWR _401_/Y sky130_fd_sc_hd__nand2_2
X_246_ _460_/Q _475_/Q VGND VGND VPWR VPWR _247_/A sky130_fd_sc_hd__nor2_2
X_315_ _315_/A VGND VGND VPWR VPWR _468_/D sky130_fd_sc_hd__buf_2
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229_ _468_/Q VGND VGND VPWR VPWR _397_/A sky130_fd_sc_hd__inv_2
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[2\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_477_ _477_/CLK _477_/D _454_/Y VGND VGND VPWR VPWR _477_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.ibufp10 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.ibufp11/A sky130_fd_sc_hd__clkinv_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_400_ _376_/Y _406_/B VGND VGND VPWR VPWR _403_/B sky130_fd_sc_hd__nand2b_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_262_ _262_/A VGND VGND VPWR VPWR _262_/Y sky130_fd_sc_hd__inv_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _461_/Q _331_/B VGND VGND VPWR VPWR _336_/B sky130_fd_sc_hd__and2_2
X_245_ _251_/A _251_/B _235_/X VGND VGND VPWR VPWR _248_/A sky130_fd_sc_hd__a21oi_2
X_314_ _468_/Q _313_/Y _328_/B VGND VGND VPWR VPWR _315_/A sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[5\].id.delayen0 ringosc.dstage\[5\].id.delayen0/A _373_/X VGND VGND
+ VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvp_2
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_228_ _469_/Q VGND VGND VPWR VPWR _420_/A sky130_fd_sc_hd__buf_2
XFILLER_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_476_ _477_/CLK _476_/D _453_/Y VGND VGND VPWR VPWR _476_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.ibufp00 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.ibufp01/A sky130_fd_sc_hd__clkinv_2
XANTENNA__375__A2 ext_trim[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.ibufp11 ringosc.ibufp11/A VGND VGND VPWR VPWR ringosc.ibufp11/Y sky130_fd_sc_hd__clkinv_8
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _460_/Q _459_/Q _342_/A VGND VGND VPWR VPWR _331_/B sky130_fd_sc_hd__and3_2
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _462_/Q _477_/Q VGND VGND VPWR VPWR _268_/A sky130_fd_sc_hd__xor2_2
X_459_ _477_/CLK _459_/D _432_/Y VGND VGND VPWR VPWR _459_/Q sky130_fd_sc_hd__dfrtp_2
X_244_ div[2] VGND VGND VPWR VPWR _250_/A sky130_fd_sc_hd__inv_2
X_313_ _313_/A _313_/B VGND VGND VPWR VPWR _313_/Y sky130_fd_sc_hd__xnor2_2
Xringosc.dstage\[5\].id.delayen1 ringosc.dstage\[5\].id.delayen1/A _410_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
X_227_ _227_/A VGND VGND VPWR VPWR _473_/D sky130_fd_sc_hd__buf_2
XANTENNA__387__B1 ext_trim[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.ibufp01 ringosc.ibufp01/A VGND VGND VPWR VPWR _477_/CLK sky130_fd_sc_hd__clkinv_8
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_475_ _477_/CLK _475_/D _452_/Y VGND VGND VPWR VPWR _475_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ div[3] _242_/Y _249_/X _250_/Y _259_/X VGND VGND VPWR VPWR _260_/X sky130_fd_sc_hd__o2111a_2
X_389_ _352_/X ext_trim[12] _388_/X VGND VGND VPWR VPWR _389_/X sky130_fd_sc_hd__a21o_2
X_458_ _477_/CLK _458_/D _431_/Y VGND VGND VPWR VPWR _458_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__243__A div[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_243_ div[3] VGND VGND VPWR VPWR _243_/Y sky130_fd_sc_hd__inv_2
X_312_ _316_/A _316_/B _297_/B VGND VGND VPWR VPWR _313_/B sky130_fd_sc_hd__a21oi_2
X_226_ _342_/A _473_/Q _345_/S VGND VGND VPWR VPWR _227_/A sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[11\].id.delayenb0 ringosc.dstage\[11\].id.delayenb1/A _387_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvn_8
XANTENNA__411__A2 ext_trim[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_474_ _477_/CLK _474_/D _451_/Y VGND VGND VPWR VPWR _474_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__287__B1 div[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_388_ _370_/A _367_/Y _359_/B VGND VGND VPWR VPWR _388_/X sky130_fd_sc_hd__o21a_2
X_457_ _477_/CLK _457_/D _430_/Y VGND VGND VPWR VPWR _457_/Q sky130_fd_sc_hd__dfrtp_2
X_311_ _420_/A _328_/B _309_/X _310_/Y VGND VGND VPWR VPWR _469_/D sky130_fd_sc_hd__o22a_2
X_242_ _242_/A _242_/B VGND VGND VPWR VPWR _242_/Y sky130_fd_sc_hd__nor2_2
XFILLER_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_225_ _458_/Q VGND VGND VPWR VPWR _342_/A sky130_fd_sc_hd__buf_2
Xringosc.dstage\[11\].id.delayenb1 ringosc.dstage\[11\].id.delayenb1/A _423_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
XANTENNA__396__A2 ext_trim[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__378__A2 ext_trim[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__369__A2 ext_trim[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_473_ _477_/CLK _473_/D _450_/Y VGND VGND VPWR VPWR _473_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_387_ _367_/Y _359_/B _386_/Y ext_trim[11] _348_/X VGND VGND VPWR VPWR _387_/X sky130_fd_sc_hd__a32o_2
X_456_ _477_/CLK _456_/D _428_/Y VGND VGND VPWR VPWR _456_/Q sky130_fd_sc_hd__dfrtp_2
X_310_ _309_/A _309_/B _328_/B VGND VGND VPWR VPWR _310_/Y sky130_fd_sc_hd__o21ai_2
Xringosc.dstage\[2\].id.delayen0 ringosc.dstage\[2\].id.delayen0/A _363_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
Xringosc.iss.const1 VGND VGND VPWR VPWR ringosc.iss.const1/HI ringosc.iss.const1/LO
+ sky130_fd_sc_hd__conb_1
X_439_ _446_/A _442_/B VGND VGND VPWR VPWR _439_/Y sky130_fd_sc_hd__nor2_2
X_241_ _240_/A _240_/B _240_/C VGND VGND VPWR VPWR _242_/B sky130_fd_sc_hd__a21oi_2
X_224_ _224_/A VGND VGND VPWR VPWR _474_/D sky130_fd_sc_hd__buf_2
Xringosc.dstage\[6\].id.delayenb0 ringosc.dstage\[6\].id.delayenb1/A _375_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[10\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_472_ _477_/CLK _472_/D _449_/Y VGND VGND VPWR VPWR _472_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__358__A dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_386_ _406_/B _386_/B VGND VGND VPWR VPWR _386_/Y sky130_fd_sc_hd__nand2_2
X_455_ _477_/CLK _455_/D _427_/Y VGND VGND VPWR VPWR _455_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[2\].id.delayen1 ringosc.dstage\[2\].id.delayen1/A _399_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XANTENNA__423__A2 ext_trim[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_240_ _240_/A _240_/B _240_/C VGND VGND VPWR VPWR _242_/A sky130_fd_sc_hd__and3_2
X_369_ _352_/X ext_trim[4] _407_/A VGND VGND VPWR VPWR _369_/X sky130_fd_sc_hd__a21o_2
X_438_ _438_/A VGND VGND VPWR VPWR _446_/A sky130_fd_sc_hd__buf_2
X_223_ _459_/Q _474_/Q _345_/S VGND VGND VPWR VPWR _224_/A sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[6\].id.delayenb1 ringosc.dstage\[6\].id.delayenb1/A _411_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_471_ _477_/CLK _471_/D _448_/Y VGND VGND VPWR VPWR _472_/D sky130_fd_sc_hd__dfrtp_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_454_ _454_/A _454_/B VGND VGND VPWR VPWR _454_/Y sky130_fd_sc_hd__nor2_2
Xringosc.iss.delayen0 ringosc.iss.delayen0/A _389_/X VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_2
X_385_ _348_/X _283_/B _278_/D _384_/Y VGND VGND VPWR VPWR _385_/X sky130_fd_sc_hd__o31a_2
XANTENNA__417__B1 ext_trim[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_368_ _370_/A _365_/Y _367_/Y _359_/B VGND VGND VPWR VPWR _407_/A sky130_fd_sc_hd__o211a_2
X_437_ _437_/A _442_/B VGND VGND VPWR VPWR _437_/Y sky130_fd_sc_hd__nor2_2
X_299_ _466_/Q VGND VGND VPWR VPWR _370_/A sky130_fd_sc_hd__buf_2
X_222_ _222_/A VGND VGND VPWR VPWR _475_/D sky130_fd_sc_hd__buf_2
XANTENNA__399__A2 ext_trim[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[2\].id.delayenb0 ringosc.dstage\[2\].id.delayenb1/A _363_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.dstage\[6\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_470_ _477_/CLK osc _446_/Y VGND VGND VPWR VPWR _471_/D sky130_fd_sc_hd__dfrtp_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_384_ ext_trim[10] _438_/A VGND VGND VPWR VPWR _384_/Y sky130_fd_sc_hd__nand2b_2
Xringosc.iss.delayen1 ringosc.iss.delayen1/A _424_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvp_2
X_453_ _454_/A _454_/B VGND VGND VPWR VPWR _453_/Y sky130_fd_sc_hd__nor2_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_367_ _367_/A _420_/C VGND VGND VPWR VPWR _367_/Y sky130_fd_sc_hd__nand2_2
X_436_ _437_/A _442_/B VGND VGND VPWR VPWR _436_/Y sky130_fd_sc_hd__nor2_2
X_298_ _298_/A VGND VGND VPWR VPWR _406_/C sky130_fd_sc_hd__buf_2
X_221_ _460_/Q _475_/Q _345_/S VGND VGND VPWR VPWR _222_/A sky130_fd_sc_hd__mux2_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_419_ _428_/A ext_trim[21] _418_/X VGND VGND VPWR VPWR _419_/X sky130_fd_sc_hd__a21o_2
XFILLER_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[2\].id.delayenb1 ringosc.dstage\[2\].id.delayenb1/A _399_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ _379_/X ext_trim[9] _372_/X _382_/X VGND VGND VPWR VPWR _383_/X sky130_fd_sc_hd__a22o_2
X_452_ _454_/A _454_/B VGND VGND VPWR VPWR _452_/Y sky130_fd_sc_hd__nor2_2
X_435_ _437_/A _442_/B VGND VGND VPWR VPWR _435_/Y sky130_fd_sc_hd__nor2_2
X_297_ _297_/A _297_/B VGND VGND VPWR VPWR _316_/A sky130_fd_sc_hd__nor2_2
X_366_ _397_/A _376_/A VGND VGND VPWR VPWR _420_/C sky130_fd_sc_hd__and2_2
X_220_ _220_/A VGND VGND VPWR VPWR _476_/D sky130_fd_sc_hd__buf_2
X_418_ _370_/A _302_/A _401_/Y _403_/X VGND VGND VPWR VPWR _418_/X sky130_fd_sc_hd__o31a_2
X_349_ dco VGND VGND VPWR VPWR _438_/A sky130_fd_sc_hd__buf_2
Xringosc.iss.ctrlen0 _433_/B _389_/X VGND VGND VPWR VPWR ringosc.iss.ctrlen0/X sky130_fd_sc_hd__or2_2
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[1\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__380__A2 ext_trim[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_382_ _406_/C _365_/Y _367_/Y _406_/B VGND VGND VPWR VPWR _382_/X sky130_fd_sc_hd__o22a_2
X_451_ _454_/A _451_/B VGND VGND VPWR VPWR _451_/Y sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_365_ _386_/B VGND VGND VPWR VPWR _365_/Y sky130_fd_sc_hd__inv_2
X_434_ _454_/B VGND VGND VPWR VPWR _442_/B sky130_fd_sc_hd__buf_2
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_296_ _467_/Q _302_/B VGND VGND VPWR VPWR _297_/B sky130_fd_sc_hd__and2_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_417_ _374_/Y _414_/X _416_/Y ext_trim[20] _348_/X VGND VGND VPWR VPWR _417_/X sky130_fd_sc_hd__a32o_2
X_348_ dco VGND VGND VPWR VPWR _348_/X sky130_fd_sc_hd__buf_2
X_279_ _420_/B _302_/A VGND VGND VPWR VPWR _298_/A sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[7\].id.delayen0 ringosc.dstage\[7\].id.delayen0/A _378_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_18_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__374__B1 dco VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_381_ _381_/A VGND VGND VPWR VPWR _406_/B sky130_fd_sc_hd__buf_2
X_450_ _454_/A _451_/B VGND VGND VPWR VPWR _450_/Y sky130_fd_sc_hd__nor2_2
X_433_ _437_/A _433_/B VGND VGND VPWR VPWR _433_/Y sky130_fd_sc_hd__nor2_2
X_364_ _352_/X ext_trim[3] _359_/B VGND VGND VPWR VPWR _364_/X sky130_fd_sc_hd__a21o_2
X_295_ _376_/A _302_/B VGND VGND VPWR VPWR _297_/A sky130_fd_sc_hd__nor2_2
X_347_ _455_/Q _347_/B VGND VGND VPWR VPWR _455_/D sky130_fd_sc_hd__nand2b_2
X_278_ _469_/Q _376_/A _324_/B _278_/D VGND VGND VPWR VPWR _278_/Y sky130_fd_sc_hd__nand4_2
X_416_ _420_/A _416_/B VGND VGND VPWR VPWR _416_/Y sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[11\].id.delayen0 ringosc.dstage\[11\].id.delayen0/A _387_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[7\].id.delayen1 ringosc.dstage\[7\].id.delayen1/A _417_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvp_2
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_380_ _379_/X ext_trim[8] _359_/B _371_/Y VGND VGND VPWR VPWR _380_/X sky130_fd_sc_hd__a22o_2
.ends

