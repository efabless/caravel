magic
tech sky130A
magscale 1 2
timestamp 1665337263
<< metal1 >>
rect 41866 42181 41918 784786
rect 411070 42422 411076 42474
rect 411128 42462 411134 42474
rect 419718 42462 419724 42474
rect 411128 42434 419724 42462
rect 411128 42422 411134 42434
rect 419718 42422 419724 42434
rect 419776 42422 419782 42474
rect 465810 42432 465816 42484
rect 465868 42472 465874 42484
rect 474458 42472 474464 42484
rect 465868 42444 474464 42472
rect 465868 42432 465874 42444
rect 474458 42432 474464 42444
rect 474516 42432 474522 42484
rect 409230 42296 409236 42348
rect 409288 42336 409294 42348
rect 412266 42336 412272 42348
rect 409288 42308 412272 42336
rect 409288 42296 409294 42308
rect 412266 42296 412272 42308
rect 412324 42336 412330 42348
rect 415394 42336 415400 42348
rect 412324 42308 415400 42336
rect 412324 42296 412330 42308
rect 415394 42296 415400 42308
rect 415452 42296 415458 42348
rect 464004 42284 464010 42336
rect 464062 42324 464068 42336
rect 467040 42324 467046 42336
rect 464062 42296 467046 42324
rect 464062 42284 464068 42296
rect 467040 42284 467046 42296
rect 467098 42324 467104 42336
rect 470167 42324 470173 42336
rect 467098 42296 470173 42324
rect 467098 42284 467104 42296
rect 470167 42284 470173 42296
rect 470225 42284 470231 42336
rect 518802 42296 518808 42348
rect 518860 42336 518866 42348
rect 524966 42336 524972 42348
rect 518860 42308 524972 42336
rect 518860 42296 518866 42308
rect 524966 42296 524972 42308
rect 525024 42296 525030 42348
rect 675682 42181 675734 370592
rect 41866 42129 145035 42181
rect 145207 42129 195328 42181
rect 195380 42129 199653 42181
rect 199705 42129 303929 42181
rect 303981 42129 308066 42181
rect 308118 42129 358732 42181
rect 358784 42129 363053 42181
rect 363105 42129 413524 42181
rect 413576 42129 417858 42181
rect 417910 42129 468330 42181
rect 468382 42129 472656 42181
rect 472708 42129 523126 42181
rect 523178 42129 527457 42181
rect 527509 42129 675734 42181
rect 186548 42045 188522 42097
rect 188574 42045 192845 42097
rect 192897 42045 201494 42097
rect 201546 42045 202717 42097
rect 202769 42045 202775 42097
rect 295162 42045 297125 42097
rect 297177 42045 299607 42097
rect 299659 42045 305774 42097
rect 305826 42045 311317 42097
rect 311369 42045 311375 42097
rect 349962 42045 351925 42097
rect 351977 42045 354406 42097
rect 354458 42045 360570 42097
rect 360622 42045 366117 42097
rect 366169 42045 366175 42097
rect 404762 42045 406719 42097
rect 406771 42045 420917 42097
rect 420969 42045 420975 42097
rect 459562 42045 461524 42097
rect 461576 42045 475717 42097
rect 475769 42045 475775 42097
rect 514362 42045 516320 42097
rect 516372 42045 530517 42097
rect 530569 42045 530575 42097
rect 534760 42013 534812 42019
rect 186548 41961 189163 42013
rect 189215 41961 191003 42013
rect 191055 41961 192202 42013
rect 192254 41961 193489 42013
rect 193541 41961 196528 42013
rect 196580 41961 197170 42013
rect 197222 41961 197813 42013
rect 197865 41961 198368 42013
rect 198420 41961 200206 42013
rect 200258 41961 200857 42013
rect 200909 41961 205926 42013
rect 205978 41961 205984 42013
rect 295162 41961 297768 42013
rect 297820 41961 300804 42013
rect 300856 41961 301451 42013
rect 301503 41961 302094 42013
rect 302146 41961 302643 42013
rect 302695 41961 305133 42013
rect 305185 41961 306418 42013
rect 306470 41961 308809 42013
rect 308861 41961 309452 42013
rect 309504 41961 315536 42013
rect 315588 41961 315594 42013
rect 349962 41961 352568 42013
rect 352620 41961 355600 42013
rect 355652 41961 356246 42013
rect 356298 41961 356889 42013
rect 356941 41961 357444 42013
rect 357496 41961 359928 42013
rect 359980 41961 361217 42013
rect 361269 41961 363607 42013
rect 363659 41961 364252 42013
rect 364304 41961 370328 42013
rect 370380 41961 370386 42013
rect 404762 41961 407367 42013
rect 407419 41961 410398 42013
rect 410450 41961 411691 42013
rect 411743 41961 414725 42013
rect 414777 41961 416013 42013
rect 416065 41961 418404 42013
rect 418456 41961 419045 42013
rect 419097 41961 425174 42013
rect 425226 41961 425232 42013
rect 459562 41961 462162 42013
rect 462214 41961 465201 42013
rect 465253 41961 466488 42013
rect 466540 41961 469522 42013
rect 469574 41961 470810 42013
rect 470862 41961 473201 42013
rect 473253 41961 473849 42013
rect 473901 41961 479956 42013
rect 480008 41961 480014 42013
rect 514362 41961 516969 42013
rect 517021 41961 520004 42013
rect 520056 41961 521293 42013
rect 521345 41961 524328 42013
rect 524380 41961 525615 42013
rect 525667 41961 528009 42013
rect 528061 41961 528652 42013
rect 528704 41961 534760 42013
rect 534760 41955 534812 41961
rect 186548 41877 187968 41929
rect 188020 41877 195973 41929
rect 196025 41877 202162 41929
rect 295162 41877 296576 41929
rect 296628 41877 304577 41929
rect 304629 41877 310827 41929
rect 349962 41877 351375 41929
rect 351427 41877 359374 41929
rect 359426 41877 365627 41929
rect 404762 41877 406170 41929
rect 406222 41877 414174 41929
rect 414226 41877 420427 41929
rect 459562 41877 460971 41929
rect 461023 41877 468967 41929
rect 469019 41877 475227 41929
rect 514362 41877 515772 41929
rect 515824 41877 523773 41929
rect 523825 41877 530027 41929
rect 186548 41793 186683 41845
rect 186735 41793 194688 41845
rect 194740 41793 199012 41845
rect 199064 41793 202162 41845
rect 295162 41793 295283 41845
rect 295335 41793 303290 41845
rect 303342 41793 307616 41845
rect 307668 41793 310827 41845
rect 349962 41793 350086 41845
rect 350138 41793 358090 41845
rect 358142 41793 362412 41845
rect 362464 41793 365627 41845
rect 404762 41793 404877 41845
rect 404929 41793 412888 41845
rect 412940 41793 417210 41845
rect 417262 41793 420427 41845
rect 459562 41793 459678 41845
rect 459730 41793 467684 41845
rect 467736 41793 472010 41845
rect 472062 41793 475227 41845
rect 514362 41793 514487 41845
rect 514539 41793 522486 41845
rect 522538 41793 526810 41845
rect 526862 41793 530027 41845
rect 140990 40029 140996 40081
rect 141048 40074 141054 40081
rect 141986 40074 141992 40081
rect 141048 40036 141992 40074
rect 141048 40029 141054 40036
rect 141986 40029 141992 40036
rect 142044 40074 142050 40081
rect 143062 40074 143068 40081
rect 142044 40036 143068 40074
rect 142044 40029 142050 40036
rect 143062 40029 143068 40036
rect 143120 40074 143126 40081
rect 143401 40074 143407 40081
rect 143120 40036 143407 40074
rect 143120 40029 143126 40036
rect 143401 40029 143407 40036
rect 143519 40074 143525 40081
rect 144597 40074 144603 40081
rect 143519 40036 144603 40074
rect 143519 40029 143525 40036
rect 144597 40029 144603 40036
rect 144655 40029 144661 40081
<< via1 >>
rect 411076 42422 411128 42474
rect 419724 42422 419776 42474
rect 465816 42432 465868 42484
rect 474464 42432 474516 42484
rect 409236 42296 409288 42348
rect 412272 42296 412324 42348
rect 415400 42296 415452 42348
rect 464010 42284 464062 42336
rect 467046 42284 467098 42336
rect 470173 42284 470225 42336
rect 518808 42296 518860 42348
rect 524972 42296 525024 42348
rect 145035 42129 145207 42181
rect 195328 42129 195380 42181
rect 199653 42129 199705 42181
rect 303929 42129 303981 42181
rect 308066 42129 308118 42181
rect 358732 42129 358784 42181
rect 363053 42129 363105 42181
rect 413524 42129 413576 42181
rect 417858 42129 417910 42181
rect 468330 42129 468382 42181
rect 472656 42129 472708 42181
rect 523126 42129 523178 42181
rect 527457 42129 527509 42181
rect 188522 42045 188574 42097
rect 192845 42045 192897 42097
rect 201494 42045 201546 42097
rect 202717 42045 202769 42097
rect 297125 42045 297177 42097
rect 299607 42045 299659 42097
rect 305774 42045 305826 42097
rect 311317 42045 311369 42097
rect 351925 42045 351977 42097
rect 354406 42045 354458 42097
rect 360570 42045 360622 42097
rect 366117 42045 366169 42097
rect 406719 42045 406771 42097
rect 420917 42045 420969 42097
rect 461524 42045 461576 42097
rect 475717 42045 475769 42097
rect 516320 42045 516372 42097
rect 530517 42045 530569 42097
rect 189163 41961 189215 42013
rect 191003 41961 191055 42013
rect 192202 41961 192254 42013
rect 193489 41961 193541 42013
rect 196528 41961 196580 42013
rect 197170 41961 197222 42013
rect 197813 41961 197865 42013
rect 198368 41961 198420 42013
rect 200206 41961 200258 42013
rect 200857 41961 200909 42013
rect 205926 41961 205978 42013
rect 297768 41961 297820 42013
rect 300804 41961 300856 42013
rect 301451 41961 301503 42013
rect 302094 41961 302146 42013
rect 302643 41961 302695 42013
rect 305133 41961 305185 42013
rect 306418 41961 306470 42013
rect 308809 41961 308861 42013
rect 309452 41961 309504 42013
rect 315536 41961 315588 42013
rect 352568 41961 352620 42013
rect 355600 41961 355652 42013
rect 356246 41961 356298 42013
rect 356889 41961 356941 42013
rect 357444 41961 357496 42013
rect 359928 41961 359980 42013
rect 361217 41961 361269 42013
rect 363607 41961 363659 42013
rect 364252 41961 364304 42013
rect 370328 41961 370380 42013
rect 407367 41961 407419 42013
rect 410398 41961 410450 42013
rect 411691 41961 411743 42013
rect 414725 41961 414777 42013
rect 416013 41961 416065 42013
rect 418404 41961 418456 42013
rect 419045 41961 419097 42013
rect 425174 41961 425226 42013
rect 462162 41961 462214 42013
rect 465201 41961 465253 42013
rect 466488 41961 466540 42013
rect 469522 41961 469574 42013
rect 470810 41961 470862 42013
rect 473201 41961 473253 42013
rect 473849 41961 473901 42013
rect 479956 41961 480008 42013
rect 516969 41961 517021 42013
rect 520004 41961 520056 42013
rect 521293 41961 521345 42013
rect 524328 41961 524380 42013
rect 525615 41961 525667 42013
rect 528009 41961 528061 42013
rect 528652 41961 528704 42013
rect 534760 41961 534812 42013
rect 187968 41877 188020 41929
rect 195973 41877 196025 41929
rect 296576 41877 296628 41929
rect 304577 41877 304629 41929
rect 351375 41877 351427 41929
rect 359374 41877 359426 41929
rect 406170 41877 406222 41929
rect 414174 41877 414226 41929
rect 460971 41877 461023 41929
rect 468967 41877 469019 41929
rect 515772 41877 515824 41929
rect 523773 41877 523825 41929
rect 186683 41793 186735 41845
rect 194688 41793 194740 41845
rect 199012 41793 199064 41845
rect 295283 41793 295335 41845
rect 303290 41793 303342 41845
rect 307616 41793 307668 41845
rect 350086 41793 350138 41845
rect 358090 41793 358142 41845
rect 362412 41793 362464 41845
rect 404877 41793 404929 41845
rect 412888 41793 412940 41845
rect 417210 41793 417262 41845
rect 459678 41793 459730 41845
rect 467684 41793 467736 41845
rect 472010 41793 472062 41845
rect 514487 41793 514539 41845
rect 522486 41793 522538 41845
rect 526810 41793 526862 41845
rect 140996 40029 141048 40081
rect 141992 40029 142044 40081
rect 143068 40029 143120 40081
rect 143407 40029 143519 40081
rect 144603 40029 144655 40081
<< metal2 >>
rect 230499 997600 235279 998010
rect 240478 997600 245258 1002732
rect 283099 997600 287879 998010
rect 293078 997600 297858 1002732
rect 384899 997600 389679 998010
rect 394878 997600 399658 1002732
rect 675407 878047 675887 878103
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867651 675887 867707
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675407 864523 675887 864579
rect 675407 863327 675887 863383
rect 41713 799417 42193 799473
rect 41713 798221 42193 798277
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 795093 42193 795149
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 675407 788847 675887 788903
rect 41713 788377 42193 788433
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 675407 785167 675887 785223
rect 41713 784697 42193 784753
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 778451 675887 778507
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675407 775323 675887 775379
rect 675407 774127 675887 774183
rect 41713 756217 42193 756273
rect 41713 755021 42193 755077
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751893 42193 751949
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 675407 743847 675887 743903
rect 41713 743337 42193 743393
rect 675407 743295 675887 743351
rect 41713 742693 42193 742749
rect 675407 742651 675887 742707
rect 41713 742049 42193 742105
rect 675407 742007 675887 742063
rect 41713 741497 42193 741553
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 733451 675887 733507
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675407 730323 675887 730379
rect 675407 729127 675887 729183
rect 41713 713017 42193 713073
rect 41713 711821 42193 711877
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708693 42193 708749
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 675407 698847 675887 698903
rect 41713 698297 42193 698353
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 688451 675887 688507
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675407 685323 675887 685379
rect 675407 684127 675887 684183
rect 41713 669817 42193 669873
rect 41713 668621 42193 668677
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 665493 42193 665549
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 41713 655097 42193 655153
rect 675407 653647 675887 653703
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 643251 675887 643307
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675407 640123 675887 640179
rect 675407 638927 675887 638983
rect 41713 626617 42193 626673
rect 41713 625421 42193 625477
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 622293 42193 622349
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 41713 611897 42193 611953
rect 675407 608647 675887 608703
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 598251 675887 598307
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675407 595123 675887 595179
rect 675407 593927 675887 593983
rect 41713 583417 42193 583473
rect 41713 582221 42193 582277
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 579093 42193 579149
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 41713 568697 42193 568753
rect 675407 563447 675887 563503
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 553051 675887 553107
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675407 549923 675887 549979
rect 675407 548727 675887 548783
rect 41713 540217 42193 540273
rect 41713 539021 42193 539077
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535893 42193 535949
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 41713 525497 42193 525553
rect 41713 412617 42193 412673
rect 41713 411421 42193 411477
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 408293 42193 408349
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 41713 397897 42193 397953
rect 675407 386247 675887 386303
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675407 372723 675887 372779
rect 675407 371527 675887 371583
rect 41713 369417 42193 369473
rect 41713 368221 42193 368277
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 365093 42193 365149
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 41713 354697 42193 354753
rect 675407 341047 675887 341103
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675407 327523 675887 327579
rect 675407 326327 675887 326383
rect 41713 326217 42193 326273
rect 41713 325021 42193 325077
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321893 42193 321949
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 41713 311497 42193 311553
rect 675407 296047 675887 296103
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 41713 283017 42193 283073
rect 675407 282523 675887 282579
rect 41713 281821 42193 281877
rect 675407 281327 675887 281383
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278693 42193 278749
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 41713 268297 42193 268353
rect 675407 251047 675887 251103
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 41713 239817 42193 239873
rect 41713 238621 42193 238677
rect 675407 238167 675887 238223
rect 41713 237977 42193 238033
rect 675407 237523 675887 237579
rect 675407 236327 675887 236383
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 41713 225097 42193 225153
rect 675407 205847 675887 205903
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 41713 196617 42193 196673
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 41713 195421 42193 195477
rect 41713 194777 42193 194833
rect 675407 194807 675887 194863
rect 41713 192937 42193 192993
rect 675407 192967 675887 193023
rect 675407 192323 675887 192379
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 675407 191127 675887 191183
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 41713 181897 42193 181953
rect 675407 160847 675887 160903
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675407 147323 675887 147379
rect 675407 146127 675887 146183
rect 675407 115647 675887 115703
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675407 102123 675887 102179
rect 675407 100927 675887 100983
rect 465816 42484 465868 42490
rect 411076 42474 411128 42480
rect 411076 42416 411128 42422
rect 419724 42474 419776 42480
rect 465816 42426 465868 42432
rect 474464 42484 474516 42490
rect 474464 42426 474516 42432
rect 419724 42416 419776 42422
rect 409236 42348 409288 42354
rect 409236 42290 409288 42296
rect 145035 42181 145207 42187
rect 145035 42123 145207 42129
rect 140996 40081 141048 40087
rect 141992 40081 142044 40087
rect 140996 39946 141048 40029
rect 141986 40029 141992 40076
rect 143068 40081 143120 40087
rect 142044 40029 142050 40076
rect 141667 39934 141813 40000
rect 141986 39954 142050 40029
rect 143407 40081 143519 40087
rect 144603 40081 144655 40087
rect 143068 39952 143120 40029
rect 143398 39990 143407 40046
rect 143519 39990 143528 40046
rect 144603 39946 144655 40029
rect 145106 39946 145136 42123
rect 186683 41845 186735 41851
rect 186683 41787 186735 41793
rect 187327 41713 187383 42193
rect 188522 42097 188574 42103
rect 188522 42039 188574 42045
rect 192845 42097 192897 42103
rect 192845 42039 192897 42045
rect 189163 42013 189215 42019
rect 189163 41955 189215 41961
rect 191003 42013 191055 42019
rect 191003 41955 191055 41961
rect 192202 42013 192254 42019
rect 192202 41955 192254 41961
rect 193489 42013 193541 42019
rect 193489 41955 193541 41961
rect 187968 41929 188020 41935
rect 187968 41871 188020 41877
rect 194043 41713 194099 42193
rect 195331 42187 195387 42198
rect 199655 42187 199711 42199
rect 303931 42187 303987 42196
rect 195328 42181 195387 42187
rect 195380 42129 195387 42181
rect 195328 42123 195387 42129
rect 199653 42181 199711 42187
rect 199705 42129 199711 42181
rect 199653 42123 199711 42129
rect 303929 42181 303987 42187
rect 303981 42129 303987 42181
rect 303929 42123 303987 42129
rect 195331 42093 195387 42123
rect 199655 42093 199711 42123
rect 201494 42097 201546 42103
rect 201494 42039 201546 42045
rect 202717 42097 202769 42103
rect 196528 42013 196580 42019
rect 196528 41955 196580 41961
rect 197170 42013 197222 42019
rect 197170 41955 197222 41961
rect 197813 42013 197865 42019
rect 197813 41955 197865 41961
rect 198368 42013 198420 42019
rect 198368 41955 198420 41961
rect 200206 42013 200258 42019
rect 200206 41955 200258 41961
rect 200857 42013 200909 42019
rect 200857 41955 200909 41961
rect 195973 41929 196025 41935
rect 195973 41871 196025 41877
rect 194688 41845 194740 41851
rect 194688 41787 194740 41793
rect 199012 41845 199064 41851
rect 199012 41787 199064 41793
rect 202717 40938 202769 42045
rect 297125 42097 297177 42103
rect 297125 42039 297177 42045
rect 299607 42097 299659 42103
rect 299607 42039 299659 42045
rect 205926 42013 205978 42019
rect 145830 40930 145888 40937
rect 145828 40928 145888 40930
rect 145828 40872 145830 40928
rect 145886 40872 145888 40928
rect 145828 40859 145888 40872
rect 202713 40929 202773 40938
rect 205926 40927 205978 41961
rect 297768 42013 297820 42019
rect 297768 41955 297820 41961
rect 300804 42013 300856 42019
rect 300804 41955 300856 41961
rect 301451 42013 301503 42019
rect 301451 41955 301503 41961
rect 302094 42013 302146 42019
rect 302094 41955 302146 41961
rect 302643 42013 302699 42112
rect 303931 42093 303987 42123
rect 305774 42097 305826 42103
rect 305774 42039 305826 42045
rect 302695 41961 302699 42013
rect 296576 41929 296628 41935
rect 302643 41920 302699 41961
rect 305133 42013 305185 42019
rect 305133 41955 305185 41961
rect 306418 42013 306470 42019
rect 306418 41955 306470 41961
rect 304577 41929 304629 41935
rect 296576 41871 296628 41877
rect 304577 41871 304629 41877
rect 295283 41845 295335 41851
rect 295283 41787 295335 41793
rect 303290 41845 303342 41851
rect 303290 41787 303342 41793
rect 306967 41713 307023 42193
rect 308065 42181 308121 42204
rect 308065 42129 308066 42181
rect 308118 42129 308121 42181
rect 308065 42085 308121 42129
rect 308255 42085 308311 42226
rect 308065 42029 308311 42085
rect 307616 41845 307668 41851
rect 307616 41787 307668 41793
rect 308255 41746 308311 42029
rect 308809 42013 308861 42019
rect 308809 41955 308861 41961
rect 309452 42013 309504 42019
rect 309452 41955 309504 41961
rect 310095 41713 310151 42193
rect 358731 42181 358787 42196
rect 358731 42129 358732 42181
rect 358784 42129 358787 42181
rect 311317 42097 311369 42103
rect 311317 40938 311369 42045
rect 351925 42097 351977 42103
rect 351925 42039 351977 42045
rect 354406 42097 354458 42103
rect 358731 42093 358787 42129
rect 360570 42097 360622 42103
rect 354406 42039 354458 42045
rect 360570 42039 360622 42045
rect 315536 42013 315588 42019
rect 311313 40929 311373 40938
rect 315536 40937 315588 41961
rect 352568 42013 352620 42019
rect 352568 41955 352620 41961
rect 355600 42013 355652 42019
rect 355600 41955 355652 41961
rect 356246 42013 356298 42019
rect 356246 41955 356298 41961
rect 356889 42013 356941 42019
rect 356889 41955 356941 41961
rect 357444 42013 357496 42019
rect 357444 41955 357496 41961
rect 359928 42013 359980 42019
rect 359928 41955 359980 41961
rect 361217 42013 361269 42019
rect 361217 41955 361269 41961
rect 351375 41929 351427 41935
rect 351375 41871 351427 41877
rect 359374 41929 359426 41935
rect 359374 41871 359426 41877
rect 350086 41845 350138 41851
rect 350086 41787 350138 41793
rect 358090 41845 358142 41851
rect 358090 41787 358142 41793
rect 361767 41713 361823 42193
rect 363055 42187 363111 42196
rect 363053 42181 363111 42187
rect 363105 42129 363111 42181
rect 363053 42123 363111 42129
rect 363055 42093 363111 42123
rect 363607 42013 363659 42019
rect 363607 41955 363659 41961
rect 364252 42013 364304 42019
rect 364252 41955 364304 41961
rect 362412 41845 362464 41851
rect 362412 41787 362464 41793
rect 364895 41713 364951 42193
rect 366117 42097 366169 42103
rect 366117 40938 366169 42045
rect 370328 42013 370380 42019
rect 202713 40860 202773 40869
rect 205922 40918 205982 40927
rect 145852 40090 145888 40859
rect 311313 40860 311373 40869
rect 315532 40928 315592 40937
rect 315532 40859 315592 40868
rect 366113 40929 366173 40938
rect 370328 40931 370380 41961
rect 404877 41845 404929 41851
rect 404877 41787 404929 41793
rect 405527 41713 405583 42193
rect 406719 42097 406771 42103
rect 406719 42039 406771 42045
rect 407367 42013 407419 42019
rect 407367 41955 407419 41961
rect 406170 41929 406222 41935
rect 406170 41871 406222 41877
rect 409248 41776 409276 42290
rect 410398 42013 410450 42019
rect 410398 41955 410450 41961
rect 411088 41776 411116 42416
rect 412272 42348 412324 42354
rect 412272 42290 412324 42296
rect 415400 42348 415452 42354
rect 415400 42290 415452 42296
rect 412284 42193 412312 42290
rect 411691 42013 411743 42019
rect 411691 41955 411743 41961
rect 412243 41776 412312 42193
rect 413531 42187 413587 42196
rect 413524 42181 413587 42187
rect 413576 42129 413587 42181
rect 413524 42123 413587 42129
rect 413531 42091 413587 42123
rect 414725 42013 414777 42019
rect 414725 41955 414777 41961
rect 414174 41929 414226 41935
rect 414174 41871 414226 41877
rect 412888 41845 412940 41851
rect 412888 41787 412940 41793
rect 415412 41776 415440 42290
rect 419736 42193 419764 42416
rect 464010 42336 464062 42342
rect 416013 42013 416065 42019
rect 416013 41955 416065 41961
rect 412243 41713 412299 41776
rect 416567 41713 416623 42193
rect 417855 42181 417911 42192
rect 417855 42129 417858 42181
rect 417910 42129 417911 42181
rect 417855 42093 417911 42129
rect 418404 42013 418456 42019
rect 418404 41955 418456 41961
rect 419045 42013 419097 42019
rect 419045 41955 419097 41961
rect 417210 41845 417262 41851
rect 417210 41787 417262 41793
rect 419695 41776 419764 42193
rect 420917 42097 420969 42103
rect 419695 41713 419751 41776
rect 420917 40938 420969 42045
rect 425174 42013 425226 42019
rect 425174 40939 425226 41961
rect 459678 41845 459730 41851
rect 459678 41787 459730 41793
rect 460327 41713 460383 42193
rect 464010 42136 464062 42284
rect 461524 42097 461576 42103
rect 461524 42039 461576 42045
rect 462162 42013 462214 42019
rect 462162 41955 462214 41961
rect 465201 42013 465253 42019
rect 465201 41955 465253 41961
rect 460971 41929 461023 41935
rect 460971 41871 461023 41877
rect 465828 41790 465856 42426
rect 467046 42336 467098 42342
rect 467046 42193 467098 42284
rect 470173 42336 470225 42342
rect 466488 42013 466540 42019
rect 466488 41955 466540 41961
rect 465828 41762 465875 41790
rect 467043 41713 467099 42193
rect 468331 42187 468387 42201
rect 468330 42181 468387 42187
rect 468382 42129 468387 42181
rect 470173 42137 470225 42284
rect 474476 42193 474504 42426
rect 518808 42348 518860 42354
rect 518808 42290 518860 42296
rect 524972 42348 525024 42354
rect 524972 42290 525024 42296
rect 468330 42123 468387 42129
rect 468331 42091 468387 42123
rect 469522 42013 469574 42019
rect 469522 41955 469574 41961
rect 470810 42013 470862 42019
rect 470810 41955 470862 41961
rect 468967 41929 469019 41935
rect 468967 41871 469019 41877
rect 467684 41845 467736 41851
rect 467684 41787 467736 41793
rect 471367 41713 471423 42193
rect 472655 42181 472711 42191
rect 472655 42129 472656 42181
rect 472708 42129 472711 42181
rect 472655 42088 472711 42129
rect 473201 42013 473253 42019
rect 473201 41955 473253 41961
rect 473849 42013 473901 42019
rect 473849 41955 473901 41961
rect 472010 41845 472062 41851
rect 472010 41787 472062 41793
rect 474476 41762 474551 42193
rect 474495 41713 474551 41762
rect 475717 42097 475769 42103
rect 366113 40860 366173 40869
rect 370324 40922 370384 40931
rect 205922 40849 205982 40858
rect 370324 40853 370384 40862
rect 420913 40929 420973 40938
rect 420913 40860 420973 40869
rect 425170 40930 425230 40939
rect 475717 40938 475769 42045
rect 479956 42013 480008 42019
rect 479956 40941 480008 41961
rect 514487 41845 514539 41851
rect 514487 41787 514539 41793
rect 515127 41713 515183 42193
rect 516320 42097 516372 42103
rect 516320 42039 516372 42045
rect 516969 42013 517021 42019
rect 516969 41955 517021 41961
rect 515772 41929 515824 41935
rect 515772 41871 515824 41877
rect 518820 41776 518848 42290
rect 524984 42226 525012 42290
rect 520004 42013 520056 42019
rect 520004 41955 520056 41961
rect 520647 41713 520703 42193
rect 521293 42013 521345 42019
rect 521293 41955 521345 41961
rect 521843 41713 521899 42193
rect 523131 42187 523187 42207
rect 523126 42181 523187 42187
rect 523178 42129 523187 42181
rect 523126 42123 523187 42129
rect 523131 42084 523187 42123
rect 524328 42013 524380 42019
rect 524328 41955 524380 41961
rect 523773 41929 523825 41935
rect 523773 41871 523825 41877
rect 522486 41845 522538 41851
rect 522486 41787 522538 41793
rect 524971 41746 525027 42226
rect 525615 42013 525667 42019
rect 525615 41955 525667 41961
rect 526167 41713 526223 42193
rect 527455 42181 527511 42205
rect 527455 42129 527457 42181
rect 527509 42129 527511 42181
rect 527455 42076 527511 42129
rect 528009 42013 528061 42019
rect 528009 41955 528061 41961
rect 528652 42013 528704 42019
rect 528652 41955 528704 41961
rect 526810 41845 526862 41851
rect 526810 41787 526862 41793
rect 529295 41713 529351 42193
rect 530517 42097 530569 42103
rect 425170 40861 425230 40870
rect 475713 40929 475773 40938
rect 475713 40860 475773 40869
rect 479952 40932 480012 40941
rect 530517 40938 530569 42045
rect 534754 41961 534760 42013
rect 534812 41961 534818 42013
rect 479952 40863 480012 40872
rect 530513 40929 530573 40938
rect 534760 40937 534812 41961
rect 530513 40860 530573 40869
rect 534756 40928 534816 40937
rect 534756 40859 534816 40868
rect 145828 40030 145837 40090
rect 145897 40030 145906 40090
<< via2 >>
rect 143407 40029 143519 40046
rect 143407 39990 143519 40029
rect 145830 40872 145886 40928
rect 202713 40869 202773 40929
rect 205922 40858 205982 40918
rect 311313 40869 311373 40929
rect 315532 40868 315592 40928
rect 366113 40869 366173 40929
rect 370324 40862 370384 40922
rect 420913 40869 420973 40929
rect 425170 40870 425230 40930
rect 475713 40869 475773 40929
rect 479952 40872 480012 40932
rect 530513 40869 530573 40929
rect 534756 40868 534816 40928
rect 145837 40030 145897 40090
<< metal3 >>
rect 82144 997600 87144 1014070
rect 133544 997600 138544 1014070
rect 184944 997600 189944 1014070
rect 240478 997600 254800 1000736
rect 293078 997600 307400 1000736
rect 394878 997600 409200 1000736
rect 478744 997600 483744 1014070
rect 530144 997600 535144 1014070
rect 631944 997600 636944 1014070
rect 23530 960144 40000 965144
rect 677600 956656 694070 961656
rect 40694 926816 46822 926940
rect 40694 922264 44296 926816
rect 46674 922264 46822 926816
rect 40694 922151 46822 922264
rect 670760 922500 676441 922502
rect 670760 922396 676562 922500
rect 40694 921722 46782 921852
rect 40694 917302 41102 921722
rect 43472 917302 46782 921722
rect 670760 917842 674136 922396
rect 676462 917842 676562 922396
rect 670760 917700 676562 917842
rect 40694 917190 46782 917302
rect 670760 917278 676562 917410
rect 41076 916786 46822 916900
rect 41076 912234 44314 916786
rect 46692 912234 46822 916786
rect 670760 912888 670948 917278
rect 673286 912888 676562 917278
rect 670760 912748 676562 912888
rect 41076 912100 46822 912234
rect 670760 912340 676562 912449
rect 670760 907786 674164 912340
rect 676490 907786 676562 912340
rect 670760 907660 676562 907786
rect 670728 474598 676620 474700
rect 670728 469994 670920 474598
rect 673278 469994 676620 474598
rect 670728 469900 676620 469994
rect 670728 469476 676620 469600
rect 670728 465070 674138 469476
rect 676502 465070 676620 469476
rect 670728 464949 676620 465070
rect 670728 464530 676620 464649
rect 670728 460006 670960 464530
rect 673300 460006 676620 464530
rect 670728 459860 676620 460006
rect 40940 455628 46824 455740
rect 40940 451068 41108 455628
rect 43494 451068 46824 455628
rect 40940 450951 46824 451068
rect 40940 450534 46824 450651
rect 40940 446104 44290 450534
rect 46656 446104 46824 450534
rect 40940 446000 46824 446104
rect 34233 440900 39600 445700
rect 40940 445574 46824 445700
rect 40940 441014 41100 445574
rect 43486 441014 46824 445574
rect 40940 440900 46824 441014
rect 479947 40936 480017 40937
rect 145825 40930 145891 40933
rect 145825 40928 148252 40930
rect 145825 40872 145830 40928
rect 145886 40872 148252 40928
rect 145825 40870 148252 40872
rect 202708 40929 202778 40934
rect 311308 40929 311378 40934
rect 145825 40867 145891 40870
rect 202708 40869 202713 40929
rect 202773 40869 203064 40929
rect 205917 40922 205987 40923
rect 205764 40918 205988 40922
rect 202708 40864 202778 40869
rect 205764 40862 205922 40918
rect 205917 40858 205922 40862
rect 205982 40862 205988 40918
rect 311308 40869 311313 40929
rect 311373 40869 312684 40929
rect 315527 40928 315597 40933
rect 315527 40926 315532 40928
rect 311308 40864 311378 40869
rect 315382 40868 315532 40926
rect 315592 40926 315597 40928
rect 366108 40929 366178 40934
rect 420908 40929 420978 40934
rect 425165 40930 425235 40935
rect 315592 40868 315600 40926
rect 315382 40866 315600 40868
rect 366108 40869 366113 40929
rect 366173 40869 367484 40929
rect 370319 40924 370389 40927
rect 370156 40922 370389 40924
rect 315527 40863 315597 40866
rect 366108 40864 366178 40869
rect 370156 40864 370324 40922
rect 370319 40862 370324 40864
rect 370384 40862 370389 40922
rect 420908 40869 420913 40929
rect 420973 40869 422262 40929
rect 425165 40928 425170 40930
rect 424966 40870 425170 40928
rect 425230 40928 425235 40930
rect 475708 40929 475778 40934
rect 479766 40932 480018 40936
rect 425230 40870 425236 40928
rect 420908 40864 420978 40869
rect 424966 40868 425236 40870
rect 475708 40869 475713 40929
rect 475773 40869 477055 40929
rect 479766 40876 479952 40932
rect 479947 40872 479952 40876
rect 480012 40876 480018 40932
rect 530508 40929 530578 40934
rect 480012 40872 480017 40876
rect 425165 40865 425235 40868
rect 475708 40864 475778 40869
rect 479947 40867 480017 40872
rect 530508 40869 530513 40929
rect 530573 40869 531856 40929
rect 534751 40928 534821 40933
rect 534751 40924 534756 40928
rect 530508 40864 530578 40869
rect 534576 40868 534756 40924
rect 534816 40924 534821 40928
rect 534816 40868 534822 40924
rect 534576 40864 534822 40868
rect 534751 40863 534821 40864
rect 205982 40858 205987 40862
rect 205917 40853 205987 40858
rect 370319 40857 370389 40862
rect 133094 40114 144010 40174
rect 133094 39940 133154 40114
rect 143407 40051 143519 40053
rect 143402 40046 143524 40051
rect 143402 39990 143407 40046
rect 143519 39990 143524 40046
rect 143402 39948 143524 39990
rect 143950 39940 144010 40114
rect 145832 40090 145902 40104
rect 145832 40030 145837 40090
rect 145897 40030 145902 40090
rect 145832 39938 145902 40030
rect 148901 40012 149351 40022
rect 148901 39694 149144 40012
rect 149304 39694 149351 40012
rect 148901 31556 149351 39694
rect 149537 40010 149918 40022
rect 149537 39692 149644 40010
rect 149804 39692 149918 40010
rect 149537 38109 149918 39692
rect 149537 37328 149563 38109
rect 149891 37328 149918 38109
rect 149537 37296 149918 37328
rect 203701 40012 204151 40022
rect 203701 39694 203944 40012
rect 204104 39694 204151 40012
rect 148901 30799 148940 31556
rect 149305 30799 149351 31556
rect 148901 30762 149351 30799
rect 203701 31556 204151 39694
rect 204337 40010 204718 40022
rect 204337 39692 204444 40010
rect 204604 39692 204718 40010
rect 204337 38109 204718 39692
rect 204337 37328 204363 38109
rect 204691 37328 204718 38109
rect 204337 37296 204718 37328
rect 313301 40012 313751 40022
rect 313301 39694 313544 40012
rect 313704 39694 313751 40012
rect 203701 30799 203740 31556
rect 204105 30799 204151 31556
rect 203701 30762 204151 30799
rect 313301 31556 313751 39694
rect 313937 40010 314318 40022
rect 313937 39692 314044 40010
rect 314204 39692 314318 40010
rect 313937 38109 314318 39692
rect 313937 37328 313963 38109
rect 314291 37328 314318 38109
rect 313937 37296 314318 37328
rect 368101 40012 368551 40022
rect 368101 39694 368344 40012
rect 368504 39694 368551 40012
rect 313301 30799 313340 31556
rect 313705 30799 313751 31556
rect 313301 30762 313751 30799
rect 368101 31556 368551 39694
rect 368737 40010 369118 40022
rect 368737 39692 368844 40010
rect 369004 39692 369118 40010
rect 368737 38109 369118 39692
rect 368737 37328 368763 38109
rect 369091 37328 369118 38109
rect 368737 37296 369118 37328
rect 422901 40012 423351 40022
rect 422901 39694 423144 40012
rect 423304 39694 423351 40012
rect 368101 30799 368140 31556
rect 368505 30799 368551 31556
rect 368101 30762 368551 30799
rect 422901 31556 423351 39694
rect 423537 40010 423918 40022
rect 423537 39692 423644 40010
rect 423804 39692 423918 40010
rect 423537 38109 423918 39692
rect 423537 37328 423563 38109
rect 423891 37328 423918 38109
rect 423537 37296 423918 37328
rect 477701 40012 478151 40022
rect 477701 39694 477944 40012
rect 478104 39694 478151 40012
rect 422901 30799 422940 31556
rect 423305 30799 423351 31556
rect 422901 30762 423351 30799
rect 477701 31556 478151 39694
rect 478337 40010 478718 40022
rect 478337 39692 478444 40010
rect 478604 39692 478718 40010
rect 478337 38109 478718 39692
rect 478337 37328 478363 38109
rect 478691 37328 478718 38109
rect 478337 37296 478718 37328
rect 532501 40012 532951 40022
rect 532501 39694 532744 40012
rect 532904 39694 532951 40012
rect 477701 30799 477740 31556
rect 478105 30799 478151 31556
rect 477701 30762 478151 30799
rect 532501 31556 532951 39694
rect 533137 40010 533518 40022
rect 533137 39692 533244 40010
rect 533404 39692 533518 40010
rect 533137 38109 533518 39692
rect 533137 37328 533163 38109
rect 533491 37328 533518 38109
rect 533137 37296 533518 37328
rect 532501 30799 532540 31556
rect 532905 30799 532951 31556
rect 532501 30762 532951 30799
<< via3 >>
rect 44296 922264 46674 926816
rect 41102 917302 43472 921722
rect 674136 917842 676462 922396
rect 44314 912234 46692 916786
rect 670948 912888 673286 917278
rect 674164 907786 676490 912340
rect 670920 469994 673278 474598
rect 674138 465070 676502 469476
rect 670960 460006 673300 464530
rect 41108 451068 43494 455628
rect 44290 446104 46656 450534
rect 41100 441014 43486 445574
rect 149144 39694 149304 40012
rect 149644 39692 149804 40010
rect 149563 37328 149891 38109
rect 203944 39694 204104 40012
rect 148940 30799 149305 31556
rect 204444 39692 204604 40010
rect 204363 37328 204691 38109
rect 313544 39694 313704 40012
rect 203740 30799 204105 31556
rect 314044 39692 314204 40010
rect 313963 37328 314291 38109
rect 368344 39694 368504 40012
rect 313340 30799 313705 31556
rect 368844 39692 369004 40010
rect 368763 37328 369091 38109
rect 423144 39694 423304 40012
rect 368140 30799 368505 31556
rect 423644 39692 423804 40010
rect 423563 37328 423891 38109
rect 477944 39694 478104 40012
rect 422940 30799 423305 31556
rect 478444 39692 478604 40010
rect 478363 37328 478691 38109
rect 532744 39694 532904 40012
rect 477740 30799 478105 31556
rect 533244 39692 533404 40010
rect 533163 37328 533491 38109
rect 532540 30799 532905 31556
<< metal4 >>
rect 44190 926816 46788 926944
rect 44190 922264 44296 926816
rect 46674 922264 46788 926816
rect 44190 922166 46788 922264
rect 674010 922396 676620 922516
rect 41004 921722 43602 921846
rect 41004 917302 41102 921722
rect 43472 917302 43602 921722
rect 674010 917842 674136 922396
rect 676462 917842 676620 922396
rect 674010 917694 676620 917842
rect 41004 917210 43602 917302
rect 670818 917278 673422 917402
rect 44198 916786 46796 916896
rect 44198 912234 44314 916786
rect 46692 912234 46796 916786
rect 670818 912888 670948 917278
rect 673286 912888 673422 917278
rect 670818 912752 673422 912888
rect 44198 912118 46796 912234
rect 674026 912340 676636 912478
rect 674026 907786 674164 912340
rect 676490 907786 676636 912340
rect 674026 907656 676636 907786
rect 670810 474598 673416 474704
rect 670810 469994 670920 474598
rect 673278 469994 673416 474598
rect 670810 469900 673416 469994
rect 674020 469476 676628 469600
rect 674020 465070 674138 469476
rect 676502 465070 676628 469476
rect 674020 464944 676628 465070
rect 670818 464530 673420 464664
rect 670818 460006 670960 464530
rect 673300 460006 673420 464530
rect 670818 459860 673420 460006
rect 680587 459800 681277 459992
rect 688881 459800 688947 474800
rect 28653 440800 28719 455800
rect 36323 455607 37013 455799
rect 40998 455628 43584 455724
rect 40998 451068 41108 455628
rect 43494 451068 43584 455628
rect 40998 450948 43584 451068
rect 44190 450534 46796 450646
rect 44190 446104 44290 450534
rect 46656 446104 46796 450534
rect 44190 446010 46796 446104
rect 40992 445574 43578 445690
rect 40992 441014 41100 445574
rect 43486 441014 43578 445574
rect 40992 440914 43578 441014
rect 149134 40012 149314 40108
rect 149134 39694 149144 40012
rect 149304 39694 149314 40012
rect 149134 39682 149314 39694
rect 149634 40010 149814 40108
rect 149634 39692 149644 40010
rect 149804 39692 149814 40010
rect 149634 39682 149814 39692
rect 203934 40012 204114 40104
rect 203934 39694 203944 40012
rect 204104 39694 204114 40012
rect 203934 39682 204114 39694
rect 204434 40010 204614 40104
rect 204434 39692 204444 40010
rect 204604 39692 204614 40010
rect 204434 39682 204614 39692
rect 313534 40012 313714 40104
rect 313534 39694 313544 40012
rect 313704 39694 313714 40012
rect 313534 39682 313714 39694
rect 314034 40010 314214 40104
rect 314034 39692 314044 40010
rect 314204 39692 314214 40010
rect 314034 39682 314214 39692
rect 368334 40012 368514 40104
rect 368334 39694 368344 40012
rect 368504 39694 368514 40012
rect 368334 39682 368514 39694
rect 368834 40010 369014 40104
rect 368834 39692 368844 40010
rect 369004 39692 369014 40010
rect 368834 39682 369014 39692
rect 423134 40012 423314 40104
rect 423134 39694 423144 40012
rect 423304 39694 423314 40012
rect 423134 39682 423314 39694
rect 423634 40010 423814 40104
rect 423634 39692 423644 40010
rect 423804 39692 423814 40010
rect 423634 39682 423814 39692
rect 477934 40012 478114 40104
rect 477934 39694 477944 40012
rect 478104 39694 478114 40012
rect 477934 39682 478114 39694
rect 478434 40010 478614 40104
rect 478434 39692 478444 40010
rect 478604 39692 478614 40010
rect 478434 39682 478614 39692
rect 532734 40012 532914 40104
rect 532734 39694 532744 40012
rect 532904 39694 532914 40012
rect 532734 39682 532914 39694
rect 533234 40010 533414 40104
rect 533234 39692 533244 40010
rect 533404 39692 533414 40010
rect 533234 39682 533414 39692
rect 132600 36323 132792 37013
<< via4 >>
rect 44296 922264 46674 926816
rect 41102 917302 43472 921722
rect 674136 917842 676462 922396
rect 44314 912234 46692 916786
rect 670948 912888 673286 917278
rect 674164 907786 676490 912340
rect 670920 469994 673278 474598
rect 674138 465070 676502 469476
rect 670960 460006 673300 464530
rect 41108 451068 43494 455628
rect 44290 446104 46656 450534
rect 41100 441014 43486 445574
<< metal5 >>
rect 78610 1018624 90778 1030788
rect 130010 1018624 142178 1030788
rect 181410 1018624 193578 1030788
rect 231810 1018624 243978 1030788
rect 284410 1018624 296578 1030788
rect 334810 1018624 346978 1030788
rect 386210 1018624 398378 1030788
rect 475210 1018624 487378 1030788
rect 526610 1018624 538778 1030788
rect 577010 1018624 589178 1030788
rect 628410 1018624 640578 1030788
rect 6811 956610 18975 968778
rect 698624 953022 710788 965190
rect 6167 914054 19619 924934
rect 40996 921722 43596 927224
rect 40996 917302 41102 921722
rect 43472 917302 43596 921722
rect 6811 871210 18975 883378
rect 6811 829010 18975 841178
rect 6598 786640 19088 799160
rect 6598 743440 19088 755960
rect 6598 700240 19088 712760
rect 6598 657040 19088 669560
rect 6598 613840 19088 626360
rect 6598 570640 19088 583160
rect 6598 527440 19088 539960
rect 6811 484410 18975 496578
rect 40996 455628 43596 917302
rect 6167 442854 19619 453734
rect 40996 451068 41108 455628
rect 43494 451068 43596 455628
rect 40996 445574 43596 451068
rect 40996 441014 41100 445574
rect 43486 441014 43596 445574
rect 6598 399840 19088 412360
rect 6598 356640 19088 369160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 6598 227040 19088 239560
rect 6598 183840 19088 196360
rect 40996 178428 43596 441014
rect 44196 926816 46796 927224
rect 44196 922264 44296 926816
rect 46674 922264 46796 926816
rect 44196 916786 46796 922264
rect 44196 912234 44314 916786
rect 46692 912234 46796 916786
rect 44196 450534 46796 912234
rect 44196 446104 44290 450534
rect 46656 446104 46796 450534
rect 44196 178428 46796 446104
rect 670820 917278 673420 922706
rect 670820 912888 670948 917278
rect 673286 912888 673420 917278
rect 670820 474598 673420 912888
rect 670820 469994 670920 474598
rect 673278 469994 673420 474598
rect 670820 464530 673420 469994
rect 670820 460006 670960 464530
rect 673300 460006 673420 464530
rect 670820 134576 673420 460006
rect 674020 922396 676620 922706
rect 674020 917842 674136 922396
rect 676462 917842 676620 922396
rect 674020 912340 676620 917842
rect 674020 907786 674164 912340
rect 676490 907786 676620 912340
rect 697980 909666 711432 920546
rect 674020 469476 676620 907786
rect 698512 863640 711002 876160
rect 698624 819822 710788 831990
rect 698512 774440 711002 786960
rect 698512 729440 711002 741960
rect 698512 684440 711002 696960
rect 698512 639240 711002 651760
rect 698512 594240 711002 606760
rect 698512 549040 711002 561560
rect 698624 505222 710788 517390
rect 674020 465070 674138 469476
rect 676502 465070 676620 469476
rect 674020 134576 676620 465070
rect 697980 461866 711432 472746
rect 698624 417022 710788 429190
rect 698512 371840 711002 384360
rect 698512 326640 711002 339160
rect 698512 281640 711002 294160
rect 698512 236640 711002 249160
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 28653 124946 30453 125266
rect 31983 124946 32633 125266
rect 36343 125007 36993 125327
rect 6811 111610 18975 123778
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use sky130_ef_io__com_bus_slice_20um  FILLER_5 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1663859327
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1663859327
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1663859327
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1663859327
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1663859327
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1663859327
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1663859327
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_13
timestamp 1663859327
transform 1 0 72800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_14 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 76800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15
timestamp 1663859327
transform 1 0 77000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_17
timestamp 1663859327
transform 1 0 92200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1663859327
transform 1 0 96200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1663859327
transform 1 0 100200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1663859327
transform 1 0 104200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1663859327
transform 1 0 108200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1663859327
transform 1 0 112200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1663859327
transform 1 0 116200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1663859327
transform 1 0 120200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1663859327
transform 1 0 124200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_26
timestamp 1663859327
transform 1 0 128200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_27
timestamp 1663859327
transform 1 0 128400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_29
timestamp 1663859327
transform 1 0 143600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_30
timestamp 1663859327
transform 1 0 147600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1663859327
transform 1 0 151600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1663859327
transform 1 0 155600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1663859327
transform 1 0 159600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1663859327
transform 1 0 163600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1663859327
transform 1 0 167600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1663859327
transform 1 0 171600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1663859327
transform 1 0 175600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_38
timestamp 1663859327
transform 1 0 179600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_39
timestamp 1663859327
transform 1 0 179800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_41
timestamp 1663859327
transform 1 0 195000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_42
timestamp 1663859327
transform 1 0 199000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_43
timestamp 1663859327
transform 1 0 203000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1663859327
transform 1 0 207000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1663859327
transform 1 0 211000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1663859327
transform 1 0 215000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_47 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 219000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1663859327
transform 1 0 254800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1663859327
transform 1 0 258800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1663859327
transform 1 0 262800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_52
timestamp 1663859327
transform 1 0 266800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_53 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 270800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1663859327
transform 1 0 271800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1663859327
transform 1 0 272000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_56
timestamp 1663859327
transform 1 0 272200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_57
timestamp 1663859327
transform 1 0 272400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1663859327
transform 1 0 310400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1663859327
transform 1 0 314400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1663859327
transform 1 0 318400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1663859327
transform 1 0 322400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1663859327
transform 1 0 326400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_65
timestamp 1663859327
transform 1 0 330400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_66
timestamp 1663859327
transform 1 0 332400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_68
timestamp 1663859327
transform 1 0 348400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_69
timestamp 1663859327
transform 1 0 352400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_70
timestamp 1663859327
transform 1 0 356400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1663859327
transform 1 0 360400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1663859327
transform 1 0 364400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1663859327
transform 1 0 368400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1663859327
transform 1 0 412200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_79
timestamp 1663859327
transform 1 0 416200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_80
timestamp 1663859327
transform 1 0 420200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_81
timestamp 1663859327
transform 1 0 424200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_82
timestamp 1663859327
transform 1 0 428200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_83
timestamp 1663859327
transform 1 0 432200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_84
timestamp 1663859327
transform 1 0 436200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_85
timestamp 1663859327
transform 1 0 440200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1663859327
transform 1 0 444200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1663859327
transform 1 0 448200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1663859327
transform 1 0 452200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1663859327
transform 1 0 456200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1663859327
transform 1 0 460200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1663859327
transform 1 0 464200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_92
timestamp 1663859327
transform 1 0 468200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_93
timestamp 1663859327
transform 1 0 472200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_94
timestamp 1663859327
transform 1 0 473200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1663859327
transform 1 0 473400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_96
timestamp 1663859327
transform 1 0 473600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_98
timestamp 1663859327
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_99
timestamp 1663859327
transform 1 0 492800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1663859327
transform 1 0 496800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1663859327
transform 1 0 500800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1663859327
transform 1 0 504800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1663859327
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1663859327
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_105
timestamp 1663859327
transform 1 0 516800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_106
timestamp 1663859327
transform 1 0 520800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_107
timestamp 1663859327
transform 1 0 524800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_108
timestamp 1663859327
transform 1 0 525000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_110
timestamp 1663859327
transform 1 0 540200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1663859327
transform 1 0 544200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1663859327
transform 1 0 548200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1663859327
transform 1 0 552200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1663859327
transform 1 0 556200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1663859327
transform 1 0 560200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_116
timestamp 1663859327
transform 1 0 564200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_117
timestamp 1663859327
transform 1 0 568200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_118
timestamp 1663859327
transform 1 0 572200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_119
timestamp 1663859327
transform 1 0 574200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_120
timestamp 1663859327
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_121
timestamp 1663859327
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_123
timestamp 1663859327
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_124
timestamp 1663859327
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1663859327
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_126
timestamp 1663859327
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_127
timestamp 1663859327
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_128
timestamp 1663859327
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_129
timestamp 1663859327
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_130
timestamp 1663859327
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1663859327
transform 1 0 622600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_132
timestamp 1663859327
transform 1 0 626600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_133
timestamp 1663859327
transform 1 0 626800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_135
timestamp 1663859327
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_136
timestamp 1663859327
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_137
timestamp 1663859327
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_138
timestamp 1663859327
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_139
timestamp 1663859327
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_140
timestamp 1663859327
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_141
timestamp 1663859327
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_142
timestamp 1663859327
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_143
timestamp 1663859327
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_144
timestamp 1663859327
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_145
timestamp 1663859327
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_146
timestamp 1663859327
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_147
timestamp 1663859327
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_148
timestamp 1663859327
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_149
timestamp 1663859327
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_150
timestamp 1663859327
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_151
timestamp 1663859327
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_152
timestamp 1663859327
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_159
timestamp 1663859327
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_160
timestamp 1663859327
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_161
timestamp 1663859327
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_162
timestamp 1663859327
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_163
timestamp 1663859327
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_165
timestamp 1663859327
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_166
timestamp 1663859327
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_167
timestamp 1663859327
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_168
timestamp 1663859327
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_169
timestamp 1663859327
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_176
timestamp 1663859327
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_177
timestamp 1663859327
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_178
timestamp 1663859327
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_179
timestamp 1663859327
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_180
timestamp 1663859327
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_182
timestamp 1663859327
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_183
timestamp 1663859327
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_184
timestamp 1663859327
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_185
timestamp 1663859327
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_186
timestamp 1663859327
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_193
timestamp 1663859327
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_194
timestamp 1663859327
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_195
timestamp 1663859327
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_196
timestamp 1663859327
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_197
timestamp 1663859327
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_199
timestamp 1663859327
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_200
timestamp 1663859327
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_201
timestamp 1663859327
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_202
timestamp 1663859327
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_203
timestamp 1663859327
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_210
timestamp 1663859327
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_211
timestamp 1663859327
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_212
timestamp 1663859327
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_213
timestamp 1663859327
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_214
timestamp 1663859327
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_216
timestamp 1663859327
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_217
timestamp 1663859327
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_218
timestamp 1663859327
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_219
timestamp 1663859327
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_220
timestamp 1663859327
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_227
timestamp 1663859327
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_228
timestamp 1663859327
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_229
timestamp 1663859327
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_230
timestamp 1663859327
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_231
timestamp 1663859327
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_233
timestamp 1663859327
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_234
timestamp 1663859327
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_235
timestamp 1663859327
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_236
timestamp 1663859327
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_237
timestamp 1663859327
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_244
timestamp 1663859327
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_245
timestamp 1663859327
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_246
timestamp 1663859327
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_247
timestamp 1663859327
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_248
timestamp 1663859327
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_250
timestamp 1663859327
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_251
timestamp 1663859327
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_252
timestamp 1663859327
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_253
timestamp 1663859327
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_254
timestamp 1663859327
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_261
timestamp 1663859327
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_262
timestamp 1663859327
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_263
timestamp 1663859327
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_264
timestamp 1663859327
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_265
timestamp 1663859327
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_267
timestamp 1663859327
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_268
timestamp 1663859327
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_269
timestamp 1663859327
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_270
timestamp 1663859327
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_271
timestamp 1663859327
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_278
timestamp 1663859327
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_279
timestamp 1663859327
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_280
timestamp 1663859327
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_281
timestamp 1663859327
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_282
timestamp 1663859327
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_284
timestamp 1663859327
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_285
timestamp 1663859327
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_286
timestamp 1663859327
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_287
timestamp 1663859327
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_288
timestamp 1663859327
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_295
timestamp 1663859327
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_296
timestamp 1663859327
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_297
timestamp 1663859327
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_298
timestamp 1663859327
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_299
timestamp 1663859327
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_301
timestamp 1663859327
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_302
timestamp 1663859327
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_303
timestamp 1663859327
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_304
timestamp 1663859327
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_305
timestamp 1663859327
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_312
timestamp 1663859327
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_313
timestamp 1663859327
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_314
timestamp 1663859327
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_315
timestamp 1663859327
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_316
timestamp 1663859327
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_318
timestamp 1663859327
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_319
timestamp 1663859327
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_320
timestamp 1663859327
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_321
timestamp 1663859327
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_322
timestamp 1663859327
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_329
timestamp 1663859327
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_330
timestamp 1663859327
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_331
timestamp 1663859327
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_332
timestamp 1663859327
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_333
timestamp 1663859327
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_335
timestamp 1663859327
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_336
timestamp 1663859327
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_337
timestamp 1663859327
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_338
timestamp 1663859327
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_339
timestamp 1663859327
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_346
timestamp 1663859327
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_347
timestamp 1663859327
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_348
timestamp 1663859327
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_349
timestamp 1663859327
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_350
timestamp 1663859327
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_351
timestamp 1663859327
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_352
timestamp 1663859327
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_353
timestamp 1663859327
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_354
timestamp 1663859327
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_355
timestamp 1663859327
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_356
timestamp 1663859327
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_357
timestamp 1663859327
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_358
timestamp 1663859327
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_359
timestamp 1663859327
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_360
timestamp 1663859327
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_362
timestamp 1663859327
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_363
timestamp 1663859327
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_364
timestamp 1663859327
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_365
timestamp 1663859327
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_366
timestamp 1663859327
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_367
timestamp 1663859327
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_368
timestamp 1663859327
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_369
timestamp 1663859327
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_370
timestamp 1663859327
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_374
timestamp 1663859327
transform 0 -1 39593 1 0 127200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1663859327
transform 0 -1 39593 1 0 131200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_376
timestamp 1663859327
transform 0 -1 39593 1 0 135200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_377
timestamp 1663859327
transform 0 -1 39593 1 0 139200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_378
timestamp 1663859327
transform 0 -1 39593 1 0 143200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_379
timestamp 1663859327
transform 0 -1 39593 1 0 147200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_380
timestamp 1663859327
transform 0 -1 39593 1 0 151200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_381
timestamp 1663859327
transform 0 -1 39593 1 0 155200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_382
timestamp 1663859327
transform 0 -1 39593 1 0 159200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_383
timestamp 1663859327
transform 0 -1 39593 1 0 163200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1663859327
transform 0 -1 39593 1 0 167200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_385
timestamp 1663859327
transform 0 -1 39593 1 0 171200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_386
timestamp 1663859327
transform 0 -1 39593 1 0 175200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_387
timestamp 1663859327
transform 0 -1 39593 1 0 179200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_388
timestamp 1663859327
transform 0 -1 39593 1 0 181200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_389
timestamp 1663859327
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_391
timestamp 1663859327
transform 0 -1 39593 1 0 197600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_392
timestamp 1663859327
transform 0 -1 39593 1 0 201600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_393
timestamp 1663859327
transform 0 -1 39593 1 0 205600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1663859327
transform 0 -1 39593 1 0 209600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_395
timestamp 1663859327
transform 0 -1 39593 1 0 213600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_396
timestamp 1663859327
transform 0 -1 39593 1 0 217600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_397
timestamp 1663859327
transform 0 -1 39593 1 0 221600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_398
timestamp 1663859327
transform 0 -1 39593 1 0 223600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_399
timestamp 1663859327
transform 0 -1 39593 1 0 224600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_401
timestamp 1663859327
transform 0 -1 39593 1 0 240800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_402
timestamp 1663859327
transform 0 -1 39593 1 0 244800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_403
timestamp 1663859327
transform 0 -1 39593 1 0 248800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_404
timestamp 1663859327
transform 0 -1 39593 1 0 252800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1663859327
transform 0 -1 39593 1 0 256800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_406
timestamp 1663859327
transform 0 -1 39593 1 0 260800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_407
timestamp 1663859327
transform 0 -1 39593 1 0 264800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_408
timestamp 1663859327
transform 0 -1 39593 1 0 266800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_409
timestamp 1663859327
transform 0 -1 39593 1 0 267800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_411
timestamp 1663859327
transform 0 -1 39593 1 0 284000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_412
timestamp 1663859327
transform 0 -1 39593 1 0 288000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_413
timestamp 1663859327
transform 0 -1 39593 1 0 292000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_414
timestamp 1663859327
transform 0 -1 39593 1 0 296000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1663859327
transform 0 -1 39593 1 0 300000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1663859327
transform 0 -1 39593 1 0 304000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_417
timestamp 1663859327
transform 0 -1 39593 1 0 308000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_418
timestamp 1663859327
transform 0 -1 39593 1 0 310000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_419
timestamp 1663859327
transform 0 -1 39593 1 0 311000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_421
timestamp 1663859327
transform 0 -1 39593 1 0 327200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_422
timestamp 1663859327
transform 0 -1 39593 1 0 331200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_423
timestamp 1663859327
transform 0 -1 39593 1 0 335200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_424
timestamp 1663859327
transform 0 -1 39593 1 0 339200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1663859327
transform 0 -1 39593 1 0 343200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1663859327
transform 0 -1 39593 1 0 347200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_427
timestamp 1663859327
transform 0 -1 39593 1 0 351200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_428
timestamp 1663859327
transform 0 -1 39593 1 0 353200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_429
timestamp 1663859327
transform 0 -1 39593 1 0 354200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_431
timestamp 1663859327
transform 0 -1 39593 1 0 370400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_432
timestamp 1663859327
transform 0 -1 39593 1 0 374400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_433
timestamp 1663859327
transform 0 -1 39593 1 0 378400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_434
timestamp 1663859327
transform 0 -1 39593 1 0 382400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1663859327
transform 0 -1 39593 1 0 386400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1663859327
transform 0 -1 39593 1 0 390400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_437
timestamp 1663859327
transform 0 -1 39593 1 0 394400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_438
timestamp 1663859327
transform 0 -1 39593 1 0 396400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_439
timestamp 1663859327
transform 0 -1 39593 1 0 397400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_441
timestamp 1663859327
transform 0 -1 39593 1 0 413600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_442
timestamp 1663859327
transform 0 -1 39593 1 0 417600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_443
timestamp 1663859327
transform 0 -1 39593 1 0 421600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_444
timestamp 1663859327
transform 0 -1 39593 1 0 425600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1663859327
transform 0 -1 39593 1 0 429600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1663859327
transform 0 -1 39593 1 0 433600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_447
timestamp 1663859327
transform 0 -1 39593 1 0 437600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_448
timestamp 1663859327
transform 0 -1 39593 1 0 439600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_449
timestamp 1663859327
transform 0 -1 39593 1 0 440600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_451
timestamp 1663859327
transform 0 -1 39593 1 0 455800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_452
timestamp 1663859327
transform 0 -1 39593 1 0 459800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_453
timestamp 1663859327
transform 0 -1 39593 1 0 463800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_454
timestamp 1663859327
transform 0 -1 39593 1 0 467800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1663859327
transform 0 -1 39593 1 0 471800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1663859327
transform 0 -1 39593 1 0 475800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_457
timestamp 1663859327
transform 0 -1 39593 1 0 479800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_458
timestamp 1663859327
transform 0 -1 39593 1 0 481800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_459
timestamp 1663859327
transform 0 -1 39593 1 0 482800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_461
timestamp 1663859327
transform 0 -1 39593 1 0 498000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_462
timestamp 1663859327
transform 0 -1 39593 1 0 502000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_463
timestamp 1663859327
transform 0 -1 39593 1 0 506000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_464
timestamp 1663859327
transform 0 -1 39593 1 0 510000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1663859327
transform 0 -1 39593 1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1663859327
transform 0 -1 39593 1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_467
timestamp 1663859327
transform 0 -1 39593 1 0 522000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_468
timestamp 1663859327
transform 0 -1 39593 1 0 524000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_469
timestamp 1663859327
transform 0 -1 39593 1 0 525000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_471
timestamp 1663859327
transform 0 -1 39593 1 0 541200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_472
timestamp 1663859327
transform 0 -1 39593 1 0 545200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_473
timestamp 1663859327
transform 0 -1 39593 1 0 549200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_474
timestamp 1663859327
transform 0 -1 39593 1 0 553200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1663859327
transform 0 -1 39593 1 0 557200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1663859327
transform 0 -1 39593 1 0 561200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_477
timestamp 1663859327
transform 0 -1 39593 1 0 565200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_478
timestamp 1663859327
transform 0 -1 39593 1 0 567200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_479
timestamp 1663859327
transform 0 -1 39593 1 0 568200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_481
timestamp 1663859327
transform 0 -1 39593 1 0 584400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_482
timestamp 1663859327
transform 0 -1 39593 1 0 588400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_483
timestamp 1663859327
transform 0 -1 39593 1 0 592400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_484
timestamp 1663859327
transform 0 -1 39593 1 0 596400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1663859327
transform 0 -1 39593 1 0 600400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1663859327
transform 0 -1 39593 1 0 604400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_487
timestamp 1663859327
transform 0 -1 39593 1 0 608400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_488
timestamp 1663859327
transform 0 -1 39593 1 0 610400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_489
timestamp 1663859327
transform 0 -1 39593 1 0 611400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_491
timestamp 1663859327
transform 0 -1 39593 1 0 627600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_492
timestamp 1663859327
transform 0 -1 39593 1 0 631600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_493
timestamp 1663859327
transform 0 -1 39593 1 0 635600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_494
timestamp 1663859327
transform 0 -1 39593 1 0 639600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1663859327
transform 0 -1 39593 1 0 643600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1663859327
transform 0 -1 39593 1 0 647600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_497
timestamp 1663859327
transform 0 -1 39593 1 0 651600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_498
timestamp 1663859327
transform 0 -1 39593 1 0 653600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_499
timestamp 1663859327
transform 0 -1 39593 1 0 654600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_501
timestamp 1663859327
transform 0 -1 39593 1 0 670800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_502
timestamp 1663859327
transform 0 -1 39593 1 0 674800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_503
timestamp 1663859327
transform 0 -1 39593 1 0 678800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_504
timestamp 1663859327
transform 0 -1 39593 1 0 682800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1663859327
transform 0 -1 39593 1 0 686800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1663859327
transform 0 -1 39593 1 0 690800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_507
timestamp 1663859327
transform 0 -1 39593 1 0 694800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_508
timestamp 1663859327
transform 0 -1 39593 1 0 696800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_509
timestamp 1663859327
transform 0 -1 39593 1 0 697800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_511
timestamp 1663859327
transform 0 -1 39593 1 0 714000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_512
timestamp 1663859327
transform 0 -1 39593 1 0 718000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_513
timestamp 1663859327
transform 0 -1 39593 1 0 722000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_514
timestamp 1663859327
transform 0 -1 39593 1 0 726000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1663859327
transform 0 -1 39593 1 0 730000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1663859327
transform 0 -1 39593 1 0 734000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_517
timestamp 1663859327
transform 0 -1 39593 1 0 738000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_518
timestamp 1663859327
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_519
timestamp 1663859327
transform 0 -1 39593 1 0 741000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_521
timestamp 1663859327
transform 0 -1 39593 1 0 757200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_522
timestamp 1663859327
transform 0 -1 39593 1 0 761200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_523
timestamp 1663859327
transform 0 -1 39593 1 0 765200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_524
timestamp 1663859327
transform 0 -1 39593 1 0 769200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1663859327
transform 0 -1 39593 1 0 773200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1663859327
transform 0 -1 39593 1 0 777200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_527
timestamp 1663859327
transform 0 -1 39593 1 0 781200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_528
timestamp 1663859327
transform 0 -1 39593 1 0 783200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_529
timestamp 1663859327
transform 0 -1 39593 1 0 784200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_531
timestamp 1663859327
transform 0 -1 39593 1 0 800400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_532
timestamp 1663859327
transform 0 -1 39593 1 0 804400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_533
timestamp 1663859327
transform 0 -1 39593 1 0 808400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_534
timestamp 1663859327
transform 0 -1 39593 1 0 812400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1663859327
transform 0 -1 39593 1 0 816400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1663859327
transform 0 -1 39593 1 0 820400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_537
timestamp 1663859327
transform 0 -1 39593 1 0 824400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_538
timestamp 1663859327
transform 0 -1 39593 1 0 826400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_539
timestamp 1663859327
transform 0 -1 39593 1 0 827400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_541
timestamp 1663859327
transform 0 -1 39593 1 0 842600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_542
timestamp 1663859327
transform 0 -1 39593 1 0 846600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_543
timestamp 1663859327
transform 0 -1 39593 1 0 850600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_544
timestamp 1663859327
transform 0 -1 39593 1 0 854600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1663859327
transform 0 -1 39593 1 0 858600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1663859327
transform 0 -1 39593 1 0 862600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_547
timestamp 1663859327
transform 0 -1 39593 1 0 866600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_548
timestamp 1663859327
transform 0 -1 39593 1 0 868600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_549
timestamp 1663859327
transform 0 -1 39593 1 0 869600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_551
timestamp 1663859327
transform 0 -1 39593 1 0 884800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_552
timestamp 1663859327
transform 0 -1 39593 1 0 888800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_553
timestamp 1663859327
transform 0 -1 39593 1 0 892800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_554
timestamp 1663859327
transform 0 -1 39593 1 0 896800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1663859327
transform 0 -1 39593 1 0 900800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1663859327
transform 0 -1 39593 1 0 904800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_557
timestamp 1663859327
transform 0 -1 39593 1 0 908800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_558
timestamp 1663859327
transform 0 -1 39593 1 0 910800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_559
timestamp 1663859327
transform 0 -1 39593 1 0 911800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_561
timestamp 1663859327
transform 0 -1 39593 1 0 927000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_562
timestamp 1663859327
transform 0 -1 39593 1 0 931000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_563
timestamp 1663859327
transform 0 -1 39593 1 0 935000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_564
timestamp 1663859327
transform 0 -1 39593 1 0 939000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1663859327
transform 0 -1 39593 1 0 943000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1663859327
transform 0 -1 39593 1 0 947000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1663859327
transform 0 -1 39593 1 0 951000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_568
timestamp 1663859327
transform 0 -1 39593 1 0 955000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_570
timestamp 1663859327
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_571
timestamp 1663859327
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_572
timestamp 1663859327
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_573
timestamp 1663859327
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_574
timestamp 1663859327
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1663859327
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_576
timestamp 1663859327
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_577
timestamp 1663859327
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_578
timestamp 1663859327
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_579
timestamp 1663859327
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_580
timestamp 1663859327
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_581
timestamp 1663859327
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_582
timestamp 1663859327
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_583
timestamp 1663859327
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_584
timestamp 1663859327
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1663859327
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1663859327
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_587
timestamp 1663859327
transform 0 1 678007 -1 0 69000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_590
timestamp 1663859327
transform 0 1 678007 -1 0 75000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_591
timestamp 1663859327
transform 0 1 678007 -1 0 79000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_592
timestamp 1663859327
transform 0 1 678007 -1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_593
timestamp 1663859327
transform 0 1 678007 -1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_594
timestamp 1663859327
transform 0 1 678007 -1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1663859327
transform 0 1 678007 -1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1663859327
transform 0 1 678007 -1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_597
timestamp 1663859327
transform 0 1 678007 -1 0 100000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_599
timestamp 1663859327
transform 0 1 678007 -1 0 120000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_600
timestamp 1663859327
transform 0 1 678007 -1 0 124000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_601
timestamp 1663859327
transform 0 1 678007 -1 0 128000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_602
timestamp 1663859327
transform 0 1 678007 -1 0 132000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_603
timestamp 1663859327
transform 0 1 678007 -1 0 136000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_604
timestamp 1663859327
transform 0 1 678007 -1 0 140000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1663859327
transform 0 1 678007 -1 0 144000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_606
timestamp 1663859327
transform 0 1 678007 -1 0 145000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_607
timestamp 1663859327
transform 0 1 678007 -1 0 145200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_609
timestamp 1663859327
transform 0 1 678007 -1 0 165200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_610
timestamp 1663859327
transform 0 1 678007 -1 0 169200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_611
timestamp 1663859327
transform 0 1 678007 -1 0 173200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_612
timestamp 1663859327
transform 0 1 678007 -1 0 177200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_613
timestamp 1663859327
transform 0 1 678007 -1 0 181200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_614
timestamp 1663859327
transform 0 1 678007 -1 0 185200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1663859327
transform 0 1 678007 -1 0 189200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_616
timestamp 1663859327
transform 0 1 678007 -1 0 190200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1663859327
transform 0 1 678007 -1 0 210200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_619
timestamp 1663859327
transform 0 1 678007 -1 0 214200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_620
timestamp 1663859327
transform 0 1 678007 -1 0 218200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_621
timestamp 1663859327
transform 0 1 678007 -1 0 222200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_622
timestamp 1663859327
transform 0 1 678007 -1 0 226200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_623
timestamp 1663859327
transform 0 1 678007 -1 0 230200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1663859327
transform 0 1 678007 -1 0 234200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_625
timestamp 1663859327
transform 0 1 678007 -1 0 235200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_626
timestamp 1663859327
transform 0 1 678007 -1 0 235400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1663859327
transform 0 1 678007 -1 0 255400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_629
timestamp 1663859327
transform 0 1 678007 -1 0 259400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_630
timestamp 1663859327
transform 0 1 678007 -1 0 263400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_631
timestamp 1663859327
transform 0 1 678007 -1 0 267400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_632
timestamp 1663859327
transform 0 1 678007 -1 0 271400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_633
timestamp 1663859327
transform 0 1 678007 -1 0 275400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1663859327
transform 0 1 678007 -1 0 279400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_635
timestamp 1663859327
transform 0 1 678007 -1 0 280400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1663859327
transform 0 1 678007 -1 0 300400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_638
timestamp 1663859327
transform 0 1 678007 -1 0 304400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_639
timestamp 1663859327
transform 0 1 678007 -1 0 308400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_640
timestamp 1663859327
transform 0 1 678007 -1 0 312400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_641
timestamp 1663859327
transform 0 1 678007 -1 0 316400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_642
timestamp 1663859327
transform 0 1 678007 -1 0 320400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1663859327
transform 0 1 678007 -1 0 324400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_644
timestamp 1663859327
transform 0 1 678007 -1 0 325400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1663859327
transform 0 1 678007 -1 0 345400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_647
timestamp 1663859327
transform 0 1 678007 -1 0 349400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_648
timestamp 1663859327
transform 0 1 678007 -1 0 353400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_649
timestamp 1663859327
transform 0 1 678007 -1 0 357400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_650
timestamp 1663859327
transform 0 1 678007 -1 0 361400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_651
timestamp 1663859327
transform 0 1 678007 -1 0 365400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_652
timestamp 1663859327
transform 0 1 678007 -1 0 369400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_653
timestamp 1663859327
transform 0 1 678007 -1 0 370400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_654
timestamp 1663859327
transform 0 1 678007 -1 0 370600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1663859327
transform 0 1 678007 -1 0 390600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_657
timestamp 1663859327
transform 0 1 678007 -1 0 394600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_658
timestamp 1663859327
transform 0 1 678007 -1 0 398600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_659
timestamp 1663859327
transform 0 1 678007 -1 0 402600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_660
timestamp 1663859327
transform 0 1 678007 -1 0 406600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_661
timestamp 1663859327
transform 0 1 678007 -1 0 410600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1663859327
transform 0 1 678007 -1 0 414600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_663
timestamp 1663859327
transform 0 1 678007 -1 0 415600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1663859327
transform 0 1 678007 -1 0 434600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1663859327
transform 0 1 678007 -1 0 438600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_667
timestamp 1663859327
transform 0 1 678007 -1 0 442600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_668
timestamp 1663859327
transform 0 1 678007 -1 0 446600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_669
timestamp 1663859327
transform 0 1 678007 -1 0 450600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_670
timestamp 1663859327
transform 0 1 678007 -1 0 454600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1663859327
transform 0 1 678007 -1 0 458600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_672
timestamp 1663859327
transform 0 1 678007 -1 0 459600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_673
timestamp 1663859327
transform 0 1 678007 -1 0 459800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1663859327
transform 0 1 678007 -1 0 478800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_676
timestamp 1663859327
transform 0 1 678007 -1 0 482800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_677
timestamp 1663859327
transform 0 1 678007 -1 0 486800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_678
timestamp 1663859327
transform 0 1 678007 -1 0 490800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_679
timestamp 1663859327
transform 0 1 678007 -1 0 494800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_680
timestamp 1663859327
transform 0 1 678007 -1 0 498800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1663859327
transform 0 1 678007 -1 0 502800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_682
timestamp 1663859327
transform 0 1 678007 -1 0 503800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1663859327
transform 0 1 678007 -1 0 522800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_685
timestamp 1663859327
transform 0 1 678007 -1 0 526800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_686
timestamp 1663859327
transform 0 1 678007 -1 0 530800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_687
timestamp 1663859327
transform 0 1 678007 -1 0 534800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_688
timestamp 1663859327
transform 0 1 678007 -1 0 538800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_689
timestamp 1663859327
transform 0 1 678007 -1 0 542800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1663859327
transform 0 1 678007 -1 0 546800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_691
timestamp 1663859327
transform 0 1 678007 -1 0 547800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1663859327
transform 0 1 678007 -1 0 567800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1663859327
transform 0 1 678007 -1 0 571800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_695
timestamp 1663859327
transform 0 1 678007 -1 0 575800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_696
timestamp 1663859327
transform 0 1 678007 -1 0 579800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_697
timestamp 1663859327
transform 0 1 678007 -1 0 583800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_698
timestamp 1663859327
transform 0 1 678007 -1 0 587800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_699
timestamp 1663859327
transform 0 1 678007 -1 0 591800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_700
timestamp 1663859327
transform 0 1 678007 -1 0 592800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_701
timestamp 1663859327
transform 0 1 678007 -1 0 593000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1663859327
transform 0 1 678007 -1 0 613000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_704
timestamp 1663859327
transform 0 1 678007 -1 0 617000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_705
timestamp 1663859327
transform 0 1 678007 -1 0 621000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_706
timestamp 1663859327
transform 0 1 678007 -1 0 625000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_707
timestamp 1663859327
transform 0 1 678007 -1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_708
timestamp 1663859327
transform 0 1 678007 -1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1663859327
transform 0 1 678007 -1 0 637000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_710
timestamp 1663859327
transform 0 1 678007 -1 0 638000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1663859327
transform 0 1 678007 -1 0 658000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1663859327
transform 0 1 678007 -1 0 662000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_714
timestamp 1663859327
transform 0 1 678007 -1 0 666000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_715
timestamp 1663859327
transform 0 1 678007 -1 0 670000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_716
timestamp 1663859327
transform 0 1 678007 -1 0 674000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_717
timestamp 1663859327
transform 0 1 678007 -1 0 678000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1663859327
transform 0 1 678007 -1 0 682000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_719
timestamp 1663859327
transform 0 1 678007 -1 0 683000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_720
timestamp 1663859327
transform 0 1 678007 -1 0 683200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1663859327
transform 0 1 678007 -1 0 703200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_723
timestamp 1663859327
transform 0 1 678007 -1 0 707200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_724
timestamp 1663859327
transform 0 1 678007 -1 0 711200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_725
timestamp 1663859327
transform 0 1 678007 -1 0 715200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_726
timestamp 1663859327
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_727
timestamp 1663859327
transform 0 1 678007 -1 0 723200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1663859327
transform 0 1 678007 -1 0 727200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_729
timestamp 1663859327
transform 0 1 678007 -1 0 728200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1663859327
transform 0 1 678007 -1 0 748200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_732
timestamp 1663859327
transform 0 1 678007 -1 0 752200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_733
timestamp 1663859327
transform 0 1 678007 -1 0 756200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_734
timestamp 1663859327
transform 0 1 678007 -1 0 760200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_735
timestamp 1663859327
transform 0 1 678007 -1 0 764200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_736
timestamp 1663859327
transform 0 1 678007 -1 0 768200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1663859327
transform 0 1 678007 -1 0 772200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_738
timestamp 1663859327
transform 0 1 678007 -1 0 773200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1663859327
transform 0 1 678007 -1 0 793200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1663859327
transform 0 1 678007 -1 0 797200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_742
timestamp 1663859327
transform 0 1 678007 -1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_743
timestamp 1663859327
transform 0 1 678007 -1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_744
timestamp 1663859327
transform 0 1 678007 -1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_745
timestamp 1663859327
transform 0 1 678007 -1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_746
timestamp 1663859327
transform 0 1 678007 -1 0 817200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_747
timestamp 1663859327
transform 0 1 678007 -1 0 818200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_748
timestamp 1663859327
transform 0 1 678007 -1 0 818400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1663859327
transform 0 1 678007 -1 0 837400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_751
timestamp 1663859327
transform 0 1 678007 -1 0 841400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_752
timestamp 1663859327
transform 0 1 678007 -1 0 845400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_753
timestamp 1663859327
transform 0 1 678007 -1 0 849400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_754
timestamp 1663859327
transform 0 1 678007 -1 0 853400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_755
timestamp 1663859327
transform 0 1 678007 -1 0 857400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1663859327
transform 0 1 678007 -1 0 861400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_757
timestamp 1663859327
transform 0 1 678007 -1 0 862400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1663859327
transform 0 1 678007 -1 0 882400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1663859327
transform 0 1 678007 -1 0 886400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_761
timestamp 1663859327
transform 0 1 678007 -1 0 890400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_762
timestamp 1663859327
transform 0 1 678007 -1 0 894400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_763
timestamp 1663859327
transform 0 1 678007 -1 0 898400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_764
timestamp 1663859327
transform 0 1 678007 -1 0 902400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1663859327
transform 0 1 678007 -1 0 906400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_766
timestamp 1663859327
transform 0 1 678007 -1 0 907400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_767
timestamp 1663859327
transform 0 1 678007 -1 0 907600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1663859327
transform 0 1 678007 -1 0 926600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_770
timestamp 1663859327
transform 0 1 678007 -1 0 930600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_771
timestamp 1663859327
transform 0 1 678007 -1 0 934600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_772
timestamp 1663859327
transform 0 1 678007 -1 0 938600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_773
timestamp 1663859327
transform 0 1 678007 -1 0 942600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_774
timestamp 1663859327
transform 0 1 678007 -1 0 946600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1663859327
transform 0 1 678007 -1 0 950600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_776
timestamp 1663859327
transform 0 1 678007 -1 0 968600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_777
timestamp 1663859327
transform 0 1 678007 -1 0 951600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_779
timestamp 1663859327
transform 0 1 678007 -1 0 972600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_780
timestamp 1663859327
transform 0 1 678007 -1 0 976600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_781
timestamp 1663859327
transform 0 1 678007 -1 0 980600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_782
timestamp 1663859327
transform 0 1 678007 -1 0 984600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_783
timestamp 1663859327
transform 0 1 678007 -1 0 988600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1663859327
transform 0 1 678007 -1 0 992600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1663859327
transform 0 1 678007 -1 0 996600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_786
timestamp 1663859327
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB1
timestamp 1663859327
transform 0 1 678007 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB2
timestamp 1663859327
transform 0 -1 39593 1 0 126200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB3
timestamp 1663859327
transform 1 0 373400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1663859327
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3
timestamp 1663859327
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1663859327
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1663859327
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1663859327
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1663859327
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1663859327
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1663859327
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1663859327
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1663859327
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1663859327
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1663859327
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1663859327
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1663859327
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1663859327
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1663859327
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1663859327
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1663859327
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1663859327
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1663859327
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1663859327
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1663859327
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1663859327
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1663859327
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1663859327
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1663859327
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1663859327
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1663859327
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1663859327
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1663859327
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1663859327
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1663859327
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1663859327
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1663859327
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1663859327
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1663859327
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1663859327
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1663859327
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1663859327
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1663859327
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1663859327
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1663859327
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1663859327
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1663859327
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1663859327
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1663859327
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1663859327
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1663859327
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1663859327
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1663859327
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1663859327
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1663859327
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1663859327
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1663859327
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1663859327
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1663859327
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1663859327
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1663859327
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1663859327
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1663859327
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1663859327
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1663859327
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1663859327
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1663859327
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1663859327
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1663859327
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1663859327
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1663859327
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1663859327
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1663859327
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1663859327
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use chip_io_gpio_connects  chip_io_gpio_connects_0
timestamp 1665336875
transform 1 0 0 0 1 0
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_1
timestamp 1665336875
transform 1 0 0 0 1 45200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_2
timestamp 1665336875
transform 1 0 0 0 1 90200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_3
timestamp 1665336875
transform 1 0 0 0 1 135400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_4
timestamp 1665336875
transform 1 0 0 0 1 180400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_5
timestamp 1665336875
transform 1 0 0 0 1 225400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_6
timestamp 1665336875
transform 1 0 0 0 1 270600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_7
timestamp 1665336875
transform 1 0 0 0 1 447800
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_8
timestamp 1665336875
transform 1 0 0 0 1 493000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_9
timestamp 1665336875
transform 1 0 0 0 1 538000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_10
timestamp 1665336875
transform 1 0 0 0 1 583200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_11
timestamp 1665336875
transform 1 0 0 0 1 628200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_12
timestamp 1665336875
transform 1 0 0 0 1 673200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_13
timestamp 1665336875
transform 1 0 0 0 1 762400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_15
timestamp 1665336875
transform -1 0 717600 0 -1 297600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_27
timestamp 1665336875
transform -1 0 717600 0 -1 900400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_28
timestamp 1665336875
transform -1 0 717600 0 -1 857200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_29
timestamp 1665336875
transform -1 0 717600 0 -1 814000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_30
timestamp 1665336875
transform -1 0 717600 0 -1 770800
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_31
timestamp 1665336875
transform -1 0 717600 0 -1 727600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_32
timestamp 1665336875
transform -1 0 717600 0 -1 684400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_33
timestamp 1665336875
transform -1 0 717600 0 -1 641200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_34
timestamp 1665336875
transform -1 0 717600 0 -1 513600
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_35
timestamp 1665336875
transform -1 0 717600 0 -1 470400
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_36
timestamp 1665336875
transform -1 0 717600 0 -1 427200
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_37
timestamp 1665336875
transform -1 0 717600 0 -1 384000
box 675407 99896 675887 115709
use chip_io_gpio_connects  chip_io_gpio_connects_38
timestamp 1665336875
transform -1 0 717600 0 -1 340800
box 675407 99896 675887 115709
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 202400 0 -1 42193
box -32 0 16032 42193
use constant_block  constant_block_0 ../maglef
timestamp 1665254081
transform -1 0 151016 0 1 39608
box 0 496 2800 2224
use constant_block  constant_block_1
timestamp 1665254081
transform -1 0 205816 0 1 39608
box 0 496 2800 2224
use constant_block  constant_block_2
timestamp 1665254081
transform -1 0 315416 0 1 39608
box 0 496 2800 2224
use constant_block  constant_block_3
timestamp 1665254081
transform -1 0 370216 0 1 39608
box 0 496 2800 2224
use constant_block  constant_block_4
timestamp 1665254081
transform -1 0 425016 0 1 39608
box 0 496 2800 2224
use constant_block  constant_block_5
timestamp 1665254081
transform -1 0 479816 0 1 39608
box 0 496 2800 2224
use constant_block  constant_block_6
timestamp 1665254081
transform -1 0 534616 0 1 39608
box 0 496 2800 2224
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 372400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1
timestamp 1663859327
transform 0 1 678007 -1 0 70000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1663859327
transform 0 -1 39593 1 0 125200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1663859327
transform -1 0 365800 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1663859327
transform -1 0 311000 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1663859327
transform -1 0 420600 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1663859327
transform -1 0 475400 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1663859327
transform -1 0 530200 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__corner_pad  mgmt_corner\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1663859327
transform 0 1 676800 -1 0 40000
box 0 0 40000 40800
use sky130_ef_io__vccd_lvc_clamped_pad  mgmt_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 0 -1 39593 1 0 68000
box 0 -2107 17239 39593
use sky130_ef_io__vdda_hvc_clamped_pad  mgmt_vdda_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1663859327
transform 0 -1 39593 1 0 869800
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  mgmt_vssa_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 93800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped_pad  mgmt_vssd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 256200 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 584000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[1\]
timestamp 1663859327
transform 1 0 333400 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[0\]
timestamp 1663859327
transform 0 1 675407 -1 0 116000
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[1\]
timestamp 1663859327
transform 0 1 675407 -1 0 161200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[2\]
timestamp 1663859327
transform 0 1 675407 -1 0 206200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[3\]
timestamp 1663859327
transform 0 1 675407 -1 0 251400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[4\]
timestamp 1663859327
transform 0 1 675407 -1 0 296400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[5\]
timestamp 1663859327
transform 0 1 675407 -1 0 341400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[6\]
timestamp 1663859327
transform 0 1 675407 -1 0 386600
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[7\]
timestamp 1663859327
transform 0 1 675407 -1 0 563800
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[8\]
timestamp 1663859327
transform 0 1 675407 -1 0 609000
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[9\]
timestamp 1663859327
transform 0 1 675407 -1 0 654000
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[10\]
timestamp 1663859327
transform 0 1 675407 -1 0 699200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[11\]
timestamp 1663859327
transform 0 1 675407 -1 0 744200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[12\]
timestamp 1663859327
transform 0 1 675407 -1 0 789200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[13\]
timestamp 1663859327
transform 0 1 675407 -1 0 878400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[0\]
timestamp 1663859327
transform 0 -1 42193 1 0 784400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[1\]
timestamp 1663859327
transform 0 -1 42193 1 0 741200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[2\]
timestamp 1663859327
transform 0 -1 42193 1 0 698000
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[3\]
timestamp 1663859327
transform 0 -1 42193 1 0 654800
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[4\]
timestamp 1663859327
transform 0 -1 42193 1 0 611600
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[5\]
timestamp 1663859327
transform 0 -1 42193 1 0 568400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[6\]
timestamp 1663859327
transform 0 -1 42193 1 0 525200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[7\]
timestamp 1663859327
transform 0 -1 42193 1 0 397600
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[8\]
timestamp 1663859327
transform 0 -1 42193 1 0 354400
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[9\]
timestamp 1663859327
transform 0 -1 42193 1 0 311200
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[10\]
timestamp 1663859327
transform 0 -1 42193 1 0 268000
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[11\]
timestamp 1663859327
transform 0 -1 42193 1 0 224800
box -32 0 16032 42193
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[12\]
timestamp 1663859327
transform 0 -1 42193 1 0 181600
box -32 0 16032 42193
use sky130_fd_io__top_xres4v2  resetb_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform -1 0 147600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_0
timestamp 1663859327
transform 1 0 374400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_1
timestamp 1663859327
transform 1 0 409200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_2
timestamp 1663859327
transform 1 0 272600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_3
timestamp 1663859327
transform 1 0 307400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_0
timestamp 1663859327
transform 1 0 410200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_1
timestamp 1663859327
transform 1 0 308400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__analog_pad  user1_analog_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 627000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__analog_pad  user1_analog_pad\[1\]
timestamp 1663859327
transform 1 0 525200 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__analog_pad  user1_analog_pad\[2\]
timestamp 1663859327
transform 1 0 473800 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__analog_pad  user1_analog_pad\[3\]
timestamp 1663859327
transform 0 1 677600 -1 0 966600
box 0 0 15000 40000
use sky130_ef_io__top_power_hvc  user1_analog_pad_with_clamp $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 1 0 375400 0 1 998007
box 0 -407 33800 39593
use sky130_ef_io__corner_pad  user1_corner
timestamp 1663859327
transform 1 0 677600 0 1 996800
box 0 0 40000 40800
use sky130_ef_io__vccd_lvc_clamped3_pad  user1_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 0 1 678007 -1 0 922600
box 0 -2177 17187 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1663859327
transform 0 1 678007 -1 0 833400
box 0 -407 15000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1663859327
transform 0 1 678007 -1 0 518800
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1663859327
transform 1 0 575600 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1663859327
transform 0 1 678007 -1 0 430600
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  user1_vssd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1663859327
transform 0 1 678007 -1 0 474800
box 0 -2177 17187 39593
use sky130_ef_io__analog_pad  user2_analog_pad\[0\]
timestamp 1663859327
transform 1 0 180000 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__analog_pad  user2_analog_pad\[1\]
timestamp 1663859327
transform 1 0 128600 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__analog_pad  user2_analog_pad\[2\]
timestamp 1663859327
transform 1 0 77200 0 1 997600
box 0 0 15000 40000
use sky130_ef_io__analog_pad  user2_analog_pad\[3\]
timestamp 1663859327
transform 0 -1 40000 1 0 955200
box 0 0 15000 40000
use sky130_ef_io__top_power_hvc  user2_analog_pad_with_clamp\[0\]
timestamp 1663859327
transform 1 0 273600 0 1 998007
box 0 -407 33800 39593
use sky130_ef_io__top_power_hvc  user2_analog_pad_with_clamp\[1\]
timestamp 1663859327
transform 1 0 221000 0 1 998007
box 0 -407 33800 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1663859327
transform 0 -1 40800 1 0 997600
box 0 0 40000 40800
use sky130_ef_io__vccd_lvc_clamped3_pad  user2_vccd_lvclamp_pad
timestamp 1663859327
transform 0 -1 39593 1 0 912000
box 0 -2177 17187 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user2_vdda_hvclamp_pad
timestamp 1663859327
transform 0 -1 39593 1 0 483000
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user2_vssa_hvclamp_pad
timestamp 1663859327
transform 0 -1 39593 1 0 827600
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  user2_vssd_lvclamp_pad
timestamp 1663859327
transform 0 -1 39593 1 0 440800
box 0 -2177 17187 39593
<< labels >>
flabel metal5 s 187640 6598 200180 19088 6 FreeSans 320 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363580 19088 6 FreeSans 320 0 0 0 flash_clk
port 3 nsew signal tristate
flabel metal5 s 296240 6598 308780 19088 6 FreeSans 320 0 0 0 flash_csb
port 7 nsew signal tristate
flabel metal5 s 405840 6598 418380 19088 6 FreeSans 320 0 0 0 flash_io0
port 11 nsew signal bidirectional
flabel metal5 s 460640 6598 473180 19088 6 FreeSans 320 0 0 0 flash_io1
port 16 nsew signal bidirectional
flabel metal5 s 515440 6598 527980 19088 6 FreeSans 320 0 0 0 gpio
port 21 nsew signal bidirectional
flabel metal5 s 6167 70054 19619 80934 6 FreeSans 320 0 0 0 vccd_pad
port 28 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18975 6 FreeSans 320 0 0 0 vdda_pad
port 29 nsew signal bidirectional
flabel metal5 s 6811 111610 18975 123778 6 FreeSans 320 0 0 0 vddio_pad
port 30 nsew signal bidirectional
flabel metal5 s 6811 871210 18975 883378 6 FreeSans 320 0 0 0 vddio_pad2
port 31 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18975 6 FreeSans 320 0 0 0 vssa_pad
port 32 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19619 6 FreeSans 320 0 0 0 vssd_pad
port 33 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18975 6 FreeSans 320 0 0 0 vssio_pad
port 34 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030788 6 FreeSans 320 0 0 0 vssio_pad2
port 35 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113780 6 FreeSans 320 0 0 0 mprj_io[0]
port 36 nsew signal bidirectional
flabel metal2 s 675407 105803 675887 105859 0 FreeSans 320 0 0 0 mprj_io_analog_en[0]
port 37 nsew signal input
flabel metal2 s 675407 107091 675887 107147 0 FreeSans 320 0 0 0 mprj_io_analog_pol[0]
port 38 nsew signal input
flabel metal2 s 675407 110127 675887 110183 0 FreeSans 320 0 0 0 mprj_io_analog_sel[0]
port 39 nsew signal input
flabel metal2 s 675407 106447 675887 106503 0 FreeSans 320 0 0 0 mprj_io_dm[0]
port 40 nsew signal input
flabel metal2 s 675407 104607 675887 104663 0 FreeSans 320 0 0 0 mprj_io_dm[1]
port 41 nsew signal input
flabel metal2 s 675407 110771 675887 110827 0 FreeSans 320 0 0 0 mprj_io_dm[2]
port 42 nsew signal input
flabel metal2 s 675407 111415 675887 111471 0 FreeSans 320 0 0 0 mprj_io_holdover[0]
port 43 nsew signal input
flabel metal2 s 675407 114451 675887 114507 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[0]
port 44 nsew signal input
flabel metal2 s 675407 107643 675887 107699 0 FreeSans 320 0 0 0 mprj_io_inp_dis[0]
port 45 nsew signal input
flabel metal2 s 675407 115095 675887 115151 0 FreeSans 320 0 0 0 mprj_io_oeb[0]
port 46 nsew signal input
flabel metal2 s 675407 111967 675887 112023 0 FreeSans 320 0 0 0 mprj_io_out[0]
port 47 nsew signal input
flabel metal2 s 675407 102767 675887 102823 0 FreeSans 320 0 0 0 mprj_io_slow_sel[0]
port 48 nsew signal input
flabel metal2 s 675407 113807 675887 113863 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[0]
port 49 nsew signal input
flabel metal2 s 675407 100927 675887 100983 0 FreeSans 320 0 0 0 mprj_io_in[0]
port 50 nsew signal tristate
flabel metal2 s 675407 115647 675887 115703 0 FreeSans 320 0 0 0 mprj_io_in_3v3[0]
port 51 nsew signal tristate
flabel metal2 s 675407 686611 675887 686667 0 FreeSans 320 0 0 0 mprj_gpio_analog[3]
port 52 nsew signal bidirectional
flabel metal2 s 675407 688451 675887 688507 0 FreeSans 320 0 0 0 mprj_gpio_noesd[3]
port 53 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696980 6 FreeSans 320 0 0 0 mprj_io[10]
port 54 nsew signal bidirectional
flabel metal2 s 675407 689003 675887 689059 0 FreeSans 320 0 0 0 mprj_io_analog_en[10]
port 55 nsew signal input
flabel metal2 s 675407 690291 675887 690347 0 FreeSans 320 0 0 0 mprj_io_analog_pol[10]
port 56 nsew signal input
flabel metal2 s 675407 693327 675887 693383 0 FreeSans 320 0 0 0 mprj_io_analog_sel[10]
port 57 nsew signal input
flabel metal2 s 675407 689647 675887 689703 0 FreeSans 320 0 0 0 mprj_io_dm[30]
port 58 nsew signal input
flabel metal2 s 675407 687807 675887 687863 0 FreeSans 320 0 0 0 mprj_io_dm[31]
port 59 nsew signal input
flabel metal2 s 675407 693971 675887 694027 0 FreeSans 320 0 0 0 mprj_io_dm[32]
port 60 nsew signal input
flabel metal2 s 675407 694615 675887 694671 0 FreeSans 320 0 0 0 mprj_io_holdover[10]
port 61 nsew signal input
flabel metal2 s 675407 697651 675887 697707 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[10]
port 62 nsew signal input
flabel metal2 s 675407 690843 675887 690899 0 FreeSans 320 0 0 0 mprj_io_inp_dis[10]
port 63 nsew signal input
flabel metal2 s 675407 698295 675887 698351 0 FreeSans 320 0 0 0 mprj_io_oeb[10]
port 64 nsew signal input
flabel metal2 s 675407 695167 675887 695223 0 FreeSans 320 0 0 0 mprj_io_out[10]
port 65 nsew signal input
flabel metal2 s 675407 685967 675887 686023 0 FreeSans 320 0 0 0 mprj_io_slow_sel[10]
port 66 nsew signal input
flabel metal2 s 675407 697007 675887 697063 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[10]
port 67 nsew signal input
flabel metal2 s 675407 684127 675887 684183 0 FreeSans 320 0 0 0 mprj_io_in[10]
port 68 nsew signal tristate
flabel metal2 s 675407 698847 675887 698903 0 FreeSans 320 0 0 0 mprj_io_in_3v3[10]
port 69 nsew signal tristate
flabel metal2 s 675407 731611 675887 731667 0 FreeSans 320 0 0 0 mprj_gpio_analog[4]
port 70 nsew signal bidirectional
flabel metal2 s 675407 733451 675887 733507 0 FreeSans 320 0 0 0 mprj_gpio_noesd[4]
port 71 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741980 6 FreeSans 320 0 0 0 mprj_io[11]
port 72 nsew signal bidirectional
flabel metal2 s 675407 734003 675887 734059 0 FreeSans 320 0 0 0 mprj_io_analog_en[11]
port 73 nsew signal input
flabel metal2 s 675407 735291 675887 735347 0 FreeSans 320 0 0 0 mprj_io_analog_pol[11]
port 74 nsew signal input
flabel metal2 s 675407 738327 675887 738383 0 FreeSans 320 0 0 0 mprj_io_analog_sel[11]
port 75 nsew signal input
flabel metal2 s 675407 734647 675887 734703 0 FreeSans 320 0 0 0 mprj_io_dm[33]
port 76 nsew signal input
flabel metal2 s 675407 732807 675887 732863 0 FreeSans 320 0 0 0 mprj_io_dm[34]
port 77 nsew signal input
flabel metal2 s 675407 738971 675887 739027 0 FreeSans 320 0 0 0 mprj_io_dm[35]
port 78 nsew signal input
flabel metal2 s 675407 739615 675887 739671 0 FreeSans 320 0 0 0 mprj_io_holdover[11]
port 79 nsew signal input
flabel metal2 s 675407 742651 675887 742707 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[11]
port 80 nsew signal input
flabel metal2 s 675407 735843 675887 735899 0 FreeSans 320 0 0 0 mprj_io_inp_dis[11]
port 81 nsew signal input
flabel metal2 s 675407 743295 675887 743351 0 FreeSans 320 0 0 0 mprj_io_oeb[11]
port 82 nsew signal input
flabel metal2 s 675407 740167 675887 740223 0 FreeSans 320 0 0 0 mprj_io_out[11]
port 83 nsew signal input
flabel metal2 s 675407 730967 675887 731023 0 FreeSans 320 0 0 0 mprj_io_slow_sel[11]
port 84 nsew signal input
flabel metal2 s 675407 742007 675887 742063 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[11]
port 85 nsew signal input
flabel metal2 s 675407 729127 675887 729183 0 FreeSans 320 0 0 0 mprj_io_in[11]
port 86 nsew signal tristate
flabel metal2 s 675407 743847 675887 743903 0 FreeSans 320 0 0 0 mprj_io_in_3v3[11]
port 87 nsew signal tristate
flabel metal2 s 675407 776611 675887 776667 0 FreeSans 320 0 0 0 mprj_gpio_analog[5]
port 88 nsew signal bidirectional
flabel metal2 s 675407 778451 675887 778507 0 FreeSans 320 0 0 0 mprj_gpio_noesd[5]
port 89 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786980 6 FreeSans 320 0 0 0 mprj_io[12]
port 90 nsew signal bidirectional
flabel metal2 s 675407 779003 675887 779059 0 FreeSans 320 0 0 0 mprj_io_analog_en[12]
port 91 nsew signal input
flabel metal2 s 675407 780291 675887 780347 0 FreeSans 320 0 0 0 mprj_io_analog_pol[12]
port 92 nsew signal input
flabel metal2 s 675407 783327 675887 783383 0 FreeSans 320 0 0 0 mprj_io_analog_sel[12]
port 93 nsew signal input
flabel metal2 s 675407 779647 675887 779703 0 FreeSans 320 0 0 0 mprj_io_dm[36]
port 94 nsew signal input
flabel metal2 s 675407 777807 675887 777863 0 FreeSans 320 0 0 0 mprj_io_dm[37]
port 95 nsew signal input
flabel metal2 s 675407 783971 675887 784027 0 FreeSans 320 0 0 0 mprj_io_dm[38]
port 96 nsew signal input
flabel metal2 s 675407 784615 675887 784671 0 FreeSans 320 0 0 0 mprj_io_holdover[12]
port 97 nsew signal input
flabel metal2 s 675407 787651 675887 787707 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[12]
port 98 nsew signal input
flabel metal2 s 675407 780843 675887 780899 0 FreeSans 320 0 0 0 mprj_io_inp_dis[12]
port 99 nsew signal input
flabel metal2 s 675407 788295 675887 788351 0 FreeSans 320 0 0 0 mprj_io_oeb[12]
port 100 nsew signal input
flabel metal2 s 675407 785167 675887 785223 0 FreeSans 320 0 0 0 mprj_io_out[12]
port 101 nsew signal input
flabel metal2 s 675407 775967 675887 776023 0 FreeSans 320 0 0 0 mprj_io_slow_sel[12]
port 102 nsew signal input
flabel metal2 s 675407 787007 675887 787063 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[12]
port 103 nsew signal input
flabel metal2 s 675407 774127 675887 774183 0 FreeSans 320 0 0 0 mprj_io_in[12]
port 104 nsew signal tristate
flabel metal2 s 675407 788847 675887 788903 0 FreeSans 320 0 0 0 mprj_io_in_3v3[12]
port 105 nsew signal tristate
flabel metal2 s 675407 865811 675887 865867 0 FreeSans 320 0 0 0 mprj_gpio_analog[6]
port 106 nsew signal bidirectional
flabel metal2 s 675407 867651 675887 867707 0 FreeSans 320 0 0 0 mprj_gpio_noesd[6]
port 107 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876180 6 FreeSans 320 0 0 0 mprj_io[13]
port 108 nsew signal bidirectional
flabel metal2 s 675407 868203 675887 868259 0 FreeSans 320 0 0 0 mprj_io_analog_en[13]
port 109 nsew signal input
flabel metal2 s 675407 869491 675887 869547 0 FreeSans 320 0 0 0 mprj_io_analog_pol[13]
port 110 nsew signal input
flabel metal2 s 675407 872527 675887 872583 0 FreeSans 320 0 0 0 mprj_io_analog_sel[13]
port 111 nsew signal input
flabel metal2 s 675407 868847 675887 868903 0 FreeSans 320 0 0 0 mprj_io_dm[39]
port 112 nsew signal input
flabel metal2 s 675407 867007 675887 867063 0 FreeSans 320 0 0 0 mprj_io_dm[40]
port 113 nsew signal input
flabel metal2 s 675407 873171 675887 873227 0 FreeSans 320 0 0 0 mprj_io_dm[41]
port 114 nsew signal input
flabel metal2 s 675407 873815 675887 873871 0 FreeSans 320 0 0 0 mprj_io_holdover[13]
port 115 nsew signal input
flabel metal2 s 675407 876851 675887 876907 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[13]
port 116 nsew signal input
flabel metal2 s 675407 870043 675887 870099 0 FreeSans 320 0 0 0 mprj_io_inp_dis[13]
port 117 nsew signal input
flabel metal2 s 675407 877495 675887 877551 0 FreeSans 320 0 0 0 mprj_io_oeb[13]
port 118 nsew signal input
flabel metal2 s 675407 874367 675887 874423 0 FreeSans 320 0 0 0 mprj_io_out[13]
port 119 nsew signal input
flabel metal2 s 675407 865167 675887 865223 0 FreeSans 320 0 0 0 mprj_io_slow_sel[13]
port 120 nsew signal input
flabel metal2 s 675407 876207 675887 876263 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[13]
port 121 nsew signal input
flabel metal2 s 675407 863327 675887 863383 0 FreeSans 320 0 0 0 mprj_io_in[13]
port 122 nsew signal tristate
flabel metal2 s 675407 878047 675887 878103 0 FreeSans 320 0 0 0 mprj_io_in_3v3[13]
port 123 nsew signal tristate
flabel metal5 s 698512 146440 711002 158980 6 FreeSans 320 0 0 0 mprj_io[1]
port 124 nsew signal bidirectional
flabel metal2 s 675407 151003 675887 151059 0 FreeSans 320 0 0 0 mprj_io_analog_en[1]
port 125 nsew signal input
flabel metal2 s 675407 152291 675887 152347 0 FreeSans 320 0 0 0 mprj_io_analog_pol[1]
port 126 nsew signal input
flabel metal2 s 675407 155327 675887 155383 0 FreeSans 320 0 0 0 mprj_io_analog_sel[1]
port 127 nsew signal input
flabel metal2 s 675407 151647 675887 151703 0 FreeSans 320 0 0 0 mprj_io_dm[3]
port 128 nsew signal input
flabel metal2 s 675407 149807 675887 149863 0 FreeSans 320 0 0 0 mprj_io_dm[4]
port 129 nsew signal input
flabel metal2 s 675407 155971 675887 156027 0 FreeSans 320 0 0 0 mprj_io_dm[5]
port 130 nsew signal input
flabel metal2 s 675407 156615 675887 156671 0 FreeSans 320 0 0 0 mprj_io_holdover[1]
port 131 nsew signal input
flabel metal2 s 675407 159651 675887 159707 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[1]
port 132 nsew signal input
flabel metal2 s 675407 152843 675887 152899 0 FreeSans 320 0 0 0 mprj_io_inp_dis[1]
port 133 nsew signal input
flabel metal2 s 675407 160295 675887 160351 0 FreeSans 320 0 0 0 mprj_io_oeb[1]
port 134 nsew signal input
flabel metal2 s 675407 157167 675887 157223 0 FreeSans 320 0 0 0 mprj_io_out[1]
port 135 nsew signal input
flabel metal2 s 675407 147967 675887 148023 0 FreeSans 320 0 0 0 mprj_io_slow_sel[1]
port 136 nsew signal input
flabel metal2 s 675407 159007 675887 159063 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[1]
port 137 nsew signal input
flabel metal2 s 675407 146127 675887 146183 0 FreeSans 320 0 0 0 mprj_io_in[1]
port 138 nsew signal tristate
flabel metal2 s 675407 160847 675887 160903 0 FreeSans 320 0 0 0 mprj_io_in_3v3[1]
port 139 nsew signal tristate
flabel metal5 s 698512 191440 711002 203980 6 FreeSans 320 0 0 0 mprj_io[2]
port 140 nsew signal bidirectional
flabel metal2 s 675407 196003 675887 196059 0 FreeSans 320 0 0 0 mprj_io_analog_en[2]
port 141 nsew signal input
flabel metal2 s 675407 197291 675887 197347 0 FreeSans 320 0 0 0 mprj_io_analog_pol[2]
port 142 nsew signal input
flabel metal2 s 675407 200327 675887 200383 0 FreeSans 320 0 0 0 mprj_io_analog_sel[2]
port 143 nsew signal input
flabel metal2 s 675407 196647 675887 196703 0 FreeSans 320 0 0 0 mprj_io_dm[6]
port 144 nsew signal input
flabel metal2 s 675407 194807 675887 194863 0 FreeSans 320 0 0 0 mprj_io_dm[7]
port 145 nsew signal input
flabel metal2 s 675407 200971 675887 201027 0 FreeSans 320 0 0 0 mprj_io_dm[8]
port 146 nsew signal input
flabel metal2 s 675407 201615 675887 201671 0 FreeSans 320 0 0 0 mprj_io_holdover[2]
port 147 nsew signal input
flabel metal2 s 675407 204651 675887 204707 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[2]
port 148 nsew signal input
flabel metal2 s 675407 197843 675887 197899 0 FreeSans 320 0 0 0 mprj_io_inp_dis[2]
port 149 nsew signal input
flabel metal2 s 675407 205295 675887 205351 0 FreeSans 320 0 0 0 mprj_io_oeb[2]
port 150 nsew signal input
flabel metal2 s 675407 202167 675887 202223 0 FreeSans 320 0 0 0 mprj_io_out[2]
port 151 nsew signal input
flabel metal2 s 675407 192967 675887 193023 0 FreeSans 320 0 0 0 mprj_io_slow_sel[2]
port 152 nsew signal input
flabel metal2 s 675407 204007 675887 204063 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[2]
port 153 nsew signal input
flabel metal2 s 675407 191127 675887 191183 0 FreeSans 320 0 0 0 mprj_io_in[2]
port 154 nsew signal tristate
flabel metal2 s 675407 205847 675887 205903 0 FreeSans 320 0 0 0 mprj_io_in_3v3[2]
port 155 nsew signal tristate
flabel metal5 s 698512 236640 711002 249180 6 FreeSans 320 0 0 0 mprj_io[3]
port 156 nsew signal bidirectional
flabel metal2 s 675407 241203 675887 241259 0 FreeSans 320 0 0 0 mprj_io_analog_en[3]
port 157 nsew signal input
flabel metal2 s 675407 242491 675887 242547 0 FreeSans 320 0 0 0 mprj_io_analog_pol[3]
port 158 nsew signal input
flabel metal2 s 675407 245527 675887 245583 0 FreeSans 320 0 0 0 mprj_io_analog_sel[3]
port 159 nsew signal input
flabel metal2 s 675407 240007 675887 240063 0 FreeSans 320 0 0 0 mprj_io_dm[10]
port 160 nsew signal input
flabel metal2 s 675407 246171 675887 246227 0 FreeSans 320 0 0 0 mprj_io_dm[11]
port 161 nsew signal input
flabel metal2 s 675407 241847 675887 241903 0 FreeSans 320 0 0 0 mprj_io_dm[9]
port 162 nsew signal input
flabel metal2 s 675407 246815 675887 246871 0 FreeSans 320 0 0 0 mprj_io_holdover[3]
port 163 nsew signal input
flabel metal2 s 675407 249851 675887 249907 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[3]
port 164 nsew signal input
flabel metal2 s 675407 243043 675887 243099 0 FreeSans 320 0 0 0 mprj_io_inp_dis[3]
port 165 nsew signal input
flabel metal2 s 675407 250495 675887 250551 0 FreeSans 320 0 0 0 mprj_io_oeb[3]
port 166 nsew signal input
flabel metal2 s 675407 247367 675887 247423 0 FreeSans 320 0 0 0 mprj_io_out[3]
port 167 nsew signal input
flabel metal2 s 675407 238167 675887 238223 0 FreeSans 320 0 0 0 mprj_io_slow_sel[3]
port 168 nsew signal input
flabel metal2 s 675407 249207 675887 249263 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[3]
port 169 nsew signal input
flabel metal2 s 675407 236327 675887 236383 0 FreeSans 320 0 0 0 mprj_io_in[3]
port 170 nsew signal tristate
flabel metal2 s 675407 251047 675887 251103 0 FreeSans 320 0 0 0 mprj_io_in_3v3[3]
port 171 nsew signal tristate
flabel metal5 s 698512 281640 711002 294180 6 FreeSans 320 0 0 0 mprj_io[4]
port 172 nsew signal bidirectional
flabel metal2 s 675407 286203 675887 286259 0 FreeSans 320 0 0 0 mprj_io_analog_en[4]
port 173 nsew signal input
flabel metal2 s 675407 287491 675887 287547 0 FreeSans 320 0 0 0 mprj_io_analog_pol[4]
port 174 nsew signal input
flabel metal2 s 675407 290527 675887 290583 0 FreeSans 320 0 0 0 mprj_io_analog_sel[4]
port 175 nsew signal input
flabel metal2 s 675407 286847 675887 286903 0 FreeSans 320 0 0 0 mprj_io_dm[12]
port 176 nsew signal input
flabel metal2 s 675407 285007 675887 285063 0 FreeSans 320 0 0 0 mprj_io_dm[13]
port 177 nsew signal input
flabel metal2 s 675407 291171 675887 291227 0 FreeSans 320 0 0 0 mprj_io_dm[14]
port 178 nsew signal input
flabel metal2 s 675407 291815 675887 291871 0 FreeSans 320 0 0 0 mprj_io_holdover[4]
port 179 nsew signal input
flabel metal2 s 675407 294851 675887 294907 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[4]
port 180 nsew signal input
flabel metal2 s 675407 288043 675887 288099 0 FreeSans 320 0 0 0 mprj_io_inp_dis[4]
port 181 nsew signal input
flabel metal2 s 675407 295495 675887 295551 0 FreeSans 320 0 0 0 mprj_io_oeb[4]
port 182 nsew signal input
flabel metal2 s 675407 292367 675887 292423 0 FreeSans 320 0 0 0 mprj_io_out[4]
port 183 nsew signal input
flabel metal2 s 675407 283167 675887 283223 0 FreeSans 320 0 0 0 mprj_io_slow_sel[4]
port 184 nsew signal input
flabel metal2 s 675407 294207 675887 294263 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[4]
port 185 nsew signal input
flabel metal2 s 675407 281327 675887 281383 0 FreeSans 320 0 0 0 mprj_io_in[4]
port 186 nsew signal tristate
flabel metal2 s 675407 296047 675887 296103 0 FreeSans 320 0 0 0 mprj_io_in_3v3[4]
port 187 nsew signal tristate
flabel metal5 s 698512 326640 711002 339180 6 FreeSans 320 0 0 0 mprj_io[5]
port 188 nsew signal bidirectional
flabel metal2 s 675407 331203 675887 331259 0 FreeSans 320 0 0 0 mprj_io_analog_en[5]
port 189 nsew signal input
flabel metal2 s 675407 332491 675887 332547 0 FreeSans 320 0 0 0 mprj_io_analog_pol[5]
port 190 nsew signal input
flabel metal2 s 675407 335527 675887 335583 0 FreeSans 320 0 0 0 mprj_io_analog_sel[5]
port 191 nsew signal input
flabel metal2 s 675407 331847 675887 331903 0 FreeSans 320 0 0 0 mprj_io_dm[15]
port 192 nsew signal input
flabel metal2 s 675407 330007 675887 330063 0 FreeSans 320 0 0 0 mprj_io_dm[16]
port 193 nsew signal input
flabel metal2 s 675407 336171 675887 336227 0 FreeSans 320 0 0 0 mprj_io_dm[17]
port 194 nsew signal input
flabel metal2 s 675407 336815 675887 336871 0 FreeSans 320 0 0 0 mprj_io_holdover[5]
port 195 nsew signal input
flabel metal2 s 675407 339851 675887 339907 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[5]
port 196 nsew signal input
flabel metal2 s 675407 333043 675887 333099 0 FreeSans 320 0 0 0 mprj_io_inp_dis[5]
port 197 nsew signal input
flabel metal2 s 675407 340495 675887 340551 0 FreeSans 320 0 0 0 mprj_io_oeb[5]
port 198 nsew signal input
flabel metal2 s 675407 337367 675887 337423 0 FreeSans 320 0 0 0 mprj_io_out[5]
port 199 nsew signal input
flabel metal2 s 675407 328167 675887 328223 0 FreeSans 320 0 0 0 mprj_io_slow_sel[5]
port 200 nsew signal input
flabel metal2 s 675407 339207 675887 339263 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[5]
port 201 nsew signal input
flabel metal2 s 675407 326327 675887 326383 0 FreeSans 320 0 0 0 mprj_io_in[5]
port 202 nsew signal tristate
flabel metal2 s 675407 341047 675887 341103 0 FreeSans 320 0 0 0 mprj_io_in_3v3[5]
port 203 nsew signal tristate
flabel metal5 s 698512 371840 711002 384380 6 FreeSans 320 0 0 0 mprj_io[6]
port 204 nsew signal bidirectional
flabel metal2 s 675407 376403 675887 376459 0 FreeSans 320 0 0 0 mprj_io_analog_en[6]
port 205 nsew signal input
flabel metal2 s 675407 377691 675887 377747 0 FreeSans 320 0 0 0 mprj_io_analog_pol[6]
port 206 nsew signal input
flabel metal2 s 675407 380727 675887 380783 0 FreeSans 320 0 0 0 mprj_io_analog_sel[6]
port 207 nsew signal input
flabel metal2 s 675407 377047 675887 377103 0 FreeSans 320 0 0 0 mprj_io_dm[18]
port 208 nsew signal input
flabel metal2 s 675407 375207 675887 375263 0 FreeSans 320 0 0 0 mprj_io_dm[19]
port 209 nsew signal input
flabel metal2 s 675407 381371 675887 381427 0 FreeSans 320 0 0 0 mprj_io_dm[20]
port 210 nsew signal input
flabel metal2 s 675407 382015 675887 382071 0 FreeSans 320 0 0 0 mprj_io_holdover[6]
port 211 nsew signal input
flabel metal2 s 675407 385051 675887 385107 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[6]
port 212 nsew signal input
flabel metal2 s 675407 378243 675887 378299 0 FreeSans 320 0 0 0 mprj_io_inp_dis[6]
port 213 nsew signal input
flabel metal2 s 675407 385695 675887 385751 0 FreeSans 320 0 0 0 mprj_io_oeb[6]
port 214 nsew signal input
flabel metal2 s 675407 382567 675887 382623 0 FreeSans 320 0 0 0 mprj_io_out[6]
port 215 nsew signal input
flabel metal2 s 675407 373367 675887 373423 0 FreeSans 320 0 0 0 mprj_io_slow_sel[6]
port 216 nsew signal input
flabel metal2 s 675407 384407 675887 384463 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[6]
port 217 nsew signal input
flabel metal2 s 675407 371527 675887 371583 0 FreeSans 320 0 0 0 mprj_io_in[6]
port 218 nsew signal tristate
flabel metal2 s 675407 386247 675887 386303 0 FreeSans 320 0 0 0 mprj_io_in_3v3[6]
port 219 nsew signal tristate
flabel metal2 s 675407 551211 675887 551267 0 FreeSans 320 0 0 0 mprj_gpio_analog[0]
port 220 nsew signal bidirectional
flabel metal2 s 675407 553051 675887 553107 0 FreeSans 320 0 0 0 mprj_gpio_noesd[0]
port 221 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561580 6 FreeSans 320 0 0 0 mprj_io[7]
port 222 nsew signal bidirectional
flabel metal2 s 675407 553603 675887 553659 0 FreeSans 320 0 0 0 mprj_io_analog_en[7]
port 223 nsew signal input
flabel metal2 s 675407 554891 675887 554947 0 FreeSans 320 0 0 0 mprj_io_analog_pol[7]
port 224 nsew signal input
flabel metal2 s 675407 557927 675887 557983 0 FreeSans 320 0 0 0 mprj_io_analog_sel[7]
port 225 nsew signal input
flabel metal2 s 675407 554247 675887 554303 0 FreeSans 320 0 0 0 mprj_io_dm[21]
port 226 nsew signal input
flabel metal2 s 675407 552407 675887 552463 0 FreeSans 320 0 0 0 mprj_io_dm[22]
port 227 nsew signal input
flabel metal2 s 675407 558571 675887 558627 0 FreeSans 320 0 0 0 mprj_io_dm[23]
port 228 nsew signal input
flabel metal2 s 675407 559215 675887 559271 0 FreeSans 320 0 0 0 mprj_io_holdover[7]
port 229 nsew signal input
flabel metal2 s 675407 562251 675887 562307 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[7]
port 230 nsew signal input
flabel metal2 s 675407 555443 675887 555499 0 FreeSans 320 0 0 0 mprj_io_inp_dis[7]
port 231 nsew signal input
flabel metal2 s 675407 562895 675887 562951 0 FreeSans 320 0 0 0 mprj_io_oeb[7]
port 232 nsew signal input
flabel metal2 s 675407 559767 675887 559823 0 FreeSans 320 0 0 0 mprj_io_out[7]
port 233 nsew signal input
flabel metal2 s 675407 550567 675887 550623 0 FreeSans 320 0 0 0 mprj_io_slow_sel[7]
port 234 nsew signal input
flabel metal2 s 675407 561607 675887 561663 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[7]
port 235 nsew signal input
flabel metal2 s 675407 548727 675887 548783 0 FreeSans 320 0 0 0 mprj_io_in[7]
port 236 nsew signal tristate
flabel metal2 s 675407 563447 675887 563503 0 FreeSans 320 0 0 0 mprj_io_in_3v3[7]
port 237 nsew signal tristate
flabel metal2 s 675407 596411 675887 596467 0 FreeSans 320 0 0 0 mprj_gpio_analog[1]
port 238 nsew signal bidirectional
flabel metal2 s 675407 598251 675887 598307 0 FreeSans 320 0 0 0 mprj_gpio_noesd[1]
port 239 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606780 6 FreeSans 320 0 0 0 mprj_io[8]
port 240 nsew signal bidirectional
flabel metal2 s 675407 598803 675887 598859 0 FreeSans 320 0 0 0 mprj_io_analog_en[8]
port 241 nsew signal input
flabel metal2 s 675407 600091 675887 600147 0 FreeSans 320 0 0 0 mprj_io_analog_pol[8]
port 242 nsew signal input
flabel metal2 s 675407 603127 675887 603183 0 FreeSans 320 0 0 0 mprj_io_analog_sel[8]
port 243 nsew signal input
flabel metal2 s 675407 599447 675887 599503 0 FreeSans 320 0 0 0 mprj_io_dm[24]
port 244 nsew signal input
flabel metal2 s 675407 597607 675887 597663 0 FreeSans 320 0 0 0 mprj_io_dm[25]
port 245 nsew signal input
flabel metal2 s 675407 603771 675887 603827 0 FreeSans 320 0 0 0 mprj_io_dm[26]
port 246 nsew signal input
flabel metal2 s 675407 604415 675887 604471 0 FreeSans 320 0 0 0 mprj_io_holdover[8]
port 247 nsew signal input
flabel metal2 s 675407 607451 675887 607507 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[8]
port 248 nsew signal input
flabel metal2 s 675407 600643 675887 600699 0 FreeSans 320 0 0 0 mprj_io_inp_dis[8]
port 249 nsew signal input
flabel metal2 s 675407 608095 675887 608151 0 FreeSans 320 0 0 0 mprj_io_oeb[8]
port 250 nsew signal input
flabel metal2 s 675407 604967 675887 605023 0 FreeSans 320 0 0 0 mprj_io_out[8]
port 251 nsew signal input
flabel metal2 s 675407 595767 675887 595823 0 FreeSans 320 0 0 0 mprj_io_slow_sel[8]
port 252 nsew signal input
flabel metal2 s 675407 606807 675887 606863 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[8]
port 253 nsew signal input
flabel metal2 s 675407 593927 675887 593983 0 FreeSans 320 0 0 0 mprj_io_in[8]
port 254 nsew signal tristate
flabel metal2 s 675407 608647 675887 608703 0 FreeSans 320 0 0 0 mprj_io_in_3v3[8]
port 255 nsew signal tristate
flabel metal2 s 675407 641411 675887 641467 0 FreeSans 320 0 0 0 mprj_gpio_analog[2]
port 256 nsew signal bidirectional
flabel metal2 s 675407 643251 675887 643307 0 FreeSans 320 0 0 0 mprj_gpio_noesd[2]
port 257 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651780 6 FreeSans 320 0 0 0 mprj_io[9]
port 258 nsew signal bidirectional
flabel metal2 s 675407 643803 675887 643859 0 FreeSans 320 0 0 0 mprj_io_analog_en[9]
port 259 nsew signal input
flabel metal2 s 675407 645091 675887 645147 0 FreeSans 320 0 0 0 mprj_io_analog_pol[9]
port 260 nsew signal input
flabel metal2 s 675407 648127 675887 648183 0 FreeSans 320 0 0 0 mprj_io_analog_sel[9]
port 261 nsew signal input
flabel metal2 s 675407 644447 675887 644503 0 FreeSans 320 0 0 0 mprj_io_dm[27]
port 262 nsew signal input
flabel metal2 s 675407 642607 675887 642663 0 FreeSans 320 0 0 0 mprj_io_dm[28]
port 263 nsew signal input
flabel metal2 s 675407 648771 675887 648827 0 FreeSans 320 0 0 0 mprj_io_dm[29]
port 264 nsew signal input
flabel metal2 s 675407 649415 675887 649471 0 FreeSans 320 0 0 0 mprj_io_holdover[9]
port 265 nsew signal input
flabel metal2 s 675407 652451 675887 652507 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[9]
port 266 nsew signal input
flabel metal2 s 675407 645643 675887 645699 0 FreeSans 320 0 0 0 mprj_io_inp_dis[9]
port 267 nsew signal input
flabel metal2 s 675407 653095 675887 653151 0 FreeSans 320 0 0 0 mprj_io_oeb[9]
port 268 nsew signal input
flabel metal2 s 675407 649967 675887 650023 0 FreeSans 320 0 0 0 mprj_io_out[9]
port 269 nsew signal input
flabel metal2 s 675407 640767 675887 640823 0 FreeSans 320 0 0 0 mprj_io_slow_sel[9]
port 270 nsew signal input
flabel metal2 s 675407 651807 675887 651863 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[9]
port 271 nsew signal input
flabel metal2 s 675407 638927 675887 638983 0 FreeSans 320 0 0 0 mprj_io_in[9]
port 272 nsew signal tristate
flabel metal2 s 675407 653647 675887 653703 0 FreeSans 320 0 0 0 mprj_io_in_3v3[9]
port 273 nsew signal tristate
flabel metal2 s 41713 796933 42193 796989 0 FreeSans 320 0 0 0 mprj_gpio_analog[7]
port 274 nsew signal bidirectional
flabel metal2 s 41713 795093 42193 795149 0 FreeSans 320 0 0 0 mprj_gpio_noesd[7]
port 275 nsew signal bidirectional
flabel metal5 s 6598 786620 19088 799160 6 FreeSans 320 0 0 0 mprj_io[25]
port 276 nsew signal bidirectional
flabel metal2 s 41713 794541 42193 794597 0 FreeSans 320 0 0 0 mprj_io_analog_en[14]
port 277 nsew signal input
flabel metal2 s 41713 793253 42193 793309 0 FreeSans 320 0 0 0 mprj_io_analog_pol[14]
port 278 nsew signal input
flabel metal2 s 41713 790217 42193 790273 0 FreeSans 320 0 0 0 mprj_io_analog_sel[14]
port 279 nsew signal input
flabel metal2 s 41713 793897 42193 793953 0 FreeSans 320 0 0 0 mprj_io_dm[42]
port 280 nsew signal input
flabel metal2 s 41713 795737 42193 795793 0 FreeSans 320 0 0 0 mprj_io_dm[43]
port 281 nsew signal input
flabel metal2 s 41713 789573 42193 789629 0 FreeSans 320 0 0 0 mprj_io_dm[44]
port 282 nsew signal input
flabel metal2 s 41713 788929 42193 788985 0 FreeSans 320 0 0 0 mprj_io_holdover[14]
port 283 nsew signal input
flabel metal2 s 41713 785893 42193 785949 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[14]
port 284 nsew signal input
flabel metal2 s 41713 792701 42193 792757 0 FreeSans 320 0 0 0 mprj_io_inp_dis[14]
port 285 nsew signal input
flabel metal2 s 41713 785249 42193 785305 0 FreeSans 320 0 0 0 mprj_io_oeb[14]
port 286 nsew signal input
flabel metal2 s 41713 788377 42193 788433 0 FreeSans 320 0 0 0 mprj_io_out[14]
port 287 nsew signal input
flabel metal2 s 41713 797577 42193 797633 0 FreeSans 320 0 0 0 mprj_io_slow_sel[14]
port 288 nsew signal input
flabel metal2 s 41713 786537 42193 786593 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[14]
port 289 nsew signal input
flabel metal2 s 41713 799417 42193 799473 0 FreeSans 320 0 0 0 mprj_io_in[14]
port 290 nsew signal tristate
flabel metal2 s 41713 784697 42193 784753 0 FreeSans 320 0 0 0 mprj_io_in_3v3[14]
port 291 nsew signal tristate
flabel metal2 s 41713 280533 42193 280589 0 FreeSans 320 0 0 0 mprj_gpio_analog[17]
port 292 nsew signal bidirectional
flabel metal2 s 41713 278693 42193 278749 0 FreeSans 320 0 0 0 mprj_gpio_noesd[17]
port 293 nsew signal bidirectional
flabel metal5 s 6598 270220 19088 282760 6 FreeSans 320 0 0 0 mprj_io[35]
port 294 nsew signal bidirectional
flabel metal2 s 41713 278141 42193 278197 0 FreeSans 320 0 0 0 mprj_io_analog_en[24]
port 295 nsew signal input
flabel metal2 s 41713 276853 42193 276909 0 FreeSans 320 0 0 0 mprj_io_analog_pol[24]
port 296 nsew signal input
flabel metal2 s 41713 273817 42193 273873 0 FreeSans 320 0 0 0 mprj_io_analog_sel[24]
port 297 nsew signal input
flabel metal2 s 41713 277497 42193 277553 0 FreeSans 320 0 0 0 mprj_io_dm[72]
port 298 nsew signal input
flabel metal2 s 41713 279337 42193 279393 0 FreeSans 320 0 0 0 mprj_io_dm[73]
port 299 nsew signal input
flabel metal2 s 41713 273173 42193 273229 0 FreeSans 320 0 0 0 mprj_io_dm[74]
port 300 nsew signal input
flabel metal2 s 41713 272529 42193 272585 0 FreeSans 320 0 0 0 mprj_io_holdover[24]
port 301 nsew signal input
flabel metal2 s 41713 269493 42193 269549 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[24]
port 302 nsew signal input
flabel metal2 s 41713 276301 42193 276357 0 FreeSans 320 0 0 0 mprj_io_inp_dis[24]
port 303 nsew signal input
flabel metal2 s 41713 268849 42193 268905 0 FreeSans 320 0 0 0 mprj_io_oeb[24]
port 304 nsew signal input
flabel metal2 s 41713 271977 42193 272033 0 FreeSans 320 0 0 0 mprj_io_out[24]
port 305 nsew signal input
flabel metal2 s 41713 281177 42193 281233 0 FreeSans 320 0 0 0 mprj_io_slow_sel[24]
port 306 nsew signal input
flabel metal2 s 41713 270137 42193 270193 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[24]
port 307 nsew signal input
flabel metal2 s 41713 283017 42193 283073 0 FreeSans 320 0 0 0 mprj_io_in[24]
port 308 nsew signal tristate
flabel metal2 s 41713 268297 42193 268353 0 FreeSans 320 0 0 0 mprj_io_in_3v3[24]
port 309 nsew signal tristate
flabel metal5 s 6598 227020 19088 239560 6 FreeSans 320 0 0 0 mprj_io[36]
port 310 nsew signal bidirectional
flabel metal2 s 41713 234941 42193 234997 0 FreeSans 320 0 0 0 mprj_io_analog_en[25]
port 311 nsew signal input
flabel metal2 s 41713 233653 42193 233709 0 FreeSans 320 0 0 0 mprj_io_analog_pol[25]
port 312 nsew signal input
flabel metal2 s 41713 230617 42193 230673 0 FreeSans 320 0 0 0 mprj_io_analog_sel[25]
port 313 nsew signal input
flabel metal2 s 41713 234297 42193 234353 0 FreeSans 320 0 0 0 mprj_io_dm[75]
port 314 nsew signal input
flabel metal2 s 41713 236137 42193 236193 0 FreeSans 320 0 0 0 mprj_io_dm[76]
port 315 nsew signal input
flabel metal2 s 41713 229973 42193 230029 0 FreeSans 320 0 0 0 mprj_io_dm[77]
port 316 nsew signal input
flabel metal2 s 41713 229329 42193 229385 0 FreeSans 320 0 0 0 mprj_io_holdover[25]
port 317 nsew signal input
flabel metal2 s 41713 226293 42193 226349 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[25]
port 318 nsew signal input
flabel metal2 s 41713 233101 42193 233157 0 FreeSans 320 0 0 0 mprj_io_inp_dis[25]
port 319 nsew signal input
flabel metal2 s 41713 225649 42193 225705 0 FreeSans 320 0 0 0 mprj_io_oeb[25]
port 320 nsew signal input
flabel metal2 s 41713 228777 42193 228833 0 FreeSans 320 0 0 0 mprj_io_out[25]
port 321 nsew signal input
flabel metal2 s 41713 237977 42193 238033 0 FreeSans 320 0 0 0 mprj_io_slow_sel[25]
port 322 nsew signal input
flabel metal2 s 41713 226937 42193 226993 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[25]
port 323 nsew signal input
flabel metal2 s 41713 239817 42193 239873 0 FreeSans 320 0 0 0 mprj_io_in[25]
port 324 nsew signal tristate
flabel metal2 s 41713 225097 42193 225153 0 FreeSans 320 0 0 0 mprj_io_in_3v3[25]
port 325 nsew signal tristate
flabel metal5 s 6598 183820 19088 196360 6 FreeSans 320 0 0 0 mprj_io[37]
port 326 nsew signal bidirectional
flabel metal2 s 41713 191741 42193 191797 0 FreeSans 320 0 0 0 mprj_io_analog_en[26]
port 327 nsew signal input
flabel metal2 s 41713 190453 42193 190509 0 FreeSans 320 0 0 0 mprj_io_analog_pol[26]
port 328 nsew signal input
flabel metal2 s 41713 187417 42193 187473 0 FreeSans 320 0 0 0 mprj_io_analog_sel[26]
port 329 nsew signal input
flabel metal2 s 41713 191097 42193 191153 0 FreeSans 320 0 0 0 mprj_io_dm[78]
port 330 nsew signal input
flabel metal2 s 41713 192937 42193 192993 0 FreeSans 320 0 0 0 mprj_io_dm[79]
port 331 nsew signal input
flabel metal2 s 41713 186773 42193 186829 0 FreeSans 320 0 0 0 mprj_io_dm[80]
port 332 nsew signal input
flabel metal2 s 41713 186129 42193 186185 0 FreeSans 320 0 0 0 mprj_io_holdover[26]
port 333 nsew signal input
flabel metal2 s 41713 183093 42193 183149 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[26]
port 334 nsew signal input
flabel metal2 s 41713 189901 42193 189957 0 FreeSans 320 0 0 0 mprj_io_inp_dis[26]
port 335 nsew signal input
flabel metal2 s 41713 182449 42193 182505 0 FreeSans 320 0 0 0 mprj_io_oeb[26]
port 336 nsew signal input
flabel metal2 s 41713 185577 42193 185633 0 FreeSans 320 0 0 0 mprj_io_out[26]
port 337 nsew signal input
flabel metal2 s 41713 194777 42193 194833 0 FreeSans 320 0 0 0 mprj_io_slow_sel[26]
port 338 nsew signal input
flabel metal2 s 41713 183737 42193 183793 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[26]
port 339 nsew signal input
flabel metal2 s 41713 196617 42193 196673 0 FreeSans 320 0 0 0 mprj_io_in[26]
port 340 nsew signal tristate
flabel metal2 s 41713 181897 42193 181953 0 FreeSans 320 0 0 0 mprj_io_in_3v3[26]
port 341 nsew signal tristate
flabel metal2 s 41713 753733 42193 753789 0 FreeSans 320 0 0 0 mprj_gpio_analog[8]
port 342 nsew signal bidirectional
flabel metal2 s 41713 751893 42193 751949 0 FreeSans 320 0 0 0 mprj_gpio_noesd[8]
port 343 nsew signal bidirectional
flabel metal5 s 6598 743420 19088 755960 6 FreeSans 320 0 0 0 mprj_io[26]
port 344 nsew signal bidirectional
flabel metal2 s 41713 751341 42193 751397 0 FreeSans 320 0 0 0 mprj_io_analog_en[15]
port 345 nsew signal input
flabel metal2 s 41713 750053 42193 750109 0 FreeSans 320 0 0 0 mprj_io_analog_pol[15]
port 346 nsew signal input
flabel metal2 s 41713 747017 42193 747073 0 FreeSans 320 0 0 0 mprj_io_analog_sel[15]
port 347 nsew signal input
flabel metal2 s 41713 750697 42193 750753 0 FreeSans 320 0 0 0 mprj_io_dm[45]
port 348 nsew signal input
flabel metal2 s 41713 752537 42193 752593 0 FreeSans 320 0 0 0 mprj_io_dm[46]
port 349 nsew signal input
flabel metal2 s 41713 746373 42193 746429 0 FreeSans 320 0 0 0 mprj_io_dm[47]
port 350 nsew signal input
flabel metal2 s 41713 745729 42193 745785 0 FreeSans 320 0 0 0 mprj_io_holdover[15]
port 351 nsew signal input
flabel metal2 s 41713 742693 42193 742749 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[15]
port 352 nsew signal input
flabel metal2 s 41713 749501 42193 749557 0 FreeSans 320 0 0 0 mprj_io_inp_dis[15]
port 353 nsew signal input
flabel metal2 s 41713 742049 42193 742105 0 FreeSans 320 0 0 0 mprj_io_oeb[15]
port 354 nsew signal input
flabel metal2 s 41713 745177 42193 745233 0 FreeSans 320 0 0 0 mprj_io_out[15]
port 355 nsew signal input
flabel metal2 s 41713 754377 42193 754433 0 FreeSans 320 0 0 0 mprj_io_slow_sel[15]
port 356 nsew signal input
flabel metal2 s 41713 743337 42193 743393 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[15]
port 357 nsew signal input
flabel metal2 s 41713 756217 42193 756273 0 FreeSans 320 0 0 0 mprj_io_in[15]
port 358 nsew signal tristate
flabel metal2 s 41713 741497 42193 741553 0 FreeSans 320 0 0 0 mprj_io_in_3v3[15]
port 359 nsew signal tristate
flabel metal2 s 41713 710533 42193 710589 0 FreeSans 320 0 0 0 mprj_gpio_analog[9]
port 360 nsew signal bidirectional
flabel metal2 s 41713 708693 42193 708749 0 FreeSans 320 0 0 0 mprj_gpio_noesd[9]
port 361 nsew signal bidirectional
flabel metal5 s 6598 700220 19088 712760 6 FreeSans 320 0 0 0 mprj_io[27]
port 362 nsew signal bidirectional
flabel metal2 s 41713 708141 42193 708197 0 FreeSans 320 0 0 0 mprj_io_analog_en[16]
port 363 nsew signal input
flabel metal2 s 41713 706853 42193 706909 0 FreeSans 320 0 0 0 mprj_io_analog_pol[16]
port 364 nsew signal input
flabel metal2 s 41713 703817 42193 703873 0 FreeSans 320 0 0 0 mprj_io_analog_sel[16]
port 365 nsew signal input
flabel metal2 s 41713 707497 42193 707553 0 FreeSans 320 0 0 0 mprj_io_dm[48]
port 366 nsew signal input
flabel metal2 s 41713 709337 42193 709393 0 FreeSans 320 0 0 0 mprj_io_dm[49]
port 367 nsew signal input
flabel metal2 s 41713 703173 42193 703229 0 FreeSans 320 0 0 0 mprj_io_dm[50]
port 368 nsew signal input
flabel metal2 s 41713 702529 42193 702585 0 FreeSans 320 0 0 0 mprj_io_holdover[16]
port 369 nsew signal input
flabel metal2 s 41713 699493 42193 699549 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[16]
port 370 nsew signal input
flabel metal2 s 41713 706301 42193 706357 0 FreeSans 320 0 0 0 mprj_io_inp_dis[16]
port 371 nsew signal input
flabel metal2 s 41713 698849 42193 698905 0 FreeSans 320 0 0 0 mprj_io_oeb[16]
port 372 nsew signal input
flabel metal2 s 41713 701977 42193 702033 0 FreeSans 320 0 0 0 mprj_io_out[16]
port 373 nsew signal input
flabel metal2 s 41713 711177 42193 711233 0 FreeSans 320 0 0 0 mprj_io_slow_sel[16]
port 374 nsew signal input
flabel metal2 s 41713 700137 42193 700193 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[16]
port 375 nsew signal input
flabel metal2 s 41713 713017 42193 713073 0 FreeSans 320 0 0 0 mprj_io_in[16]
port 376 nsew signal tristate
flabel metal2 s 41713 698297 42193 698353 0 FreeSans 320 0 0 0 mprj_io_in_3v3[16]
port 377 nsew signal tristate
flabel metal2 s 41713 667333 42193 667389 0 FreeSans 320 0 0 0 mprj_gpio_analog[10]
port 378 nsew signal bidirectional
flabel metal2 s 41713 665493 42193 665549 0 FreeSans 320 0 0 0 mprj_gpio_noesd[10]
port 379 nsew signal bidirectional
flabel metal5 s 6598 657020 19088 669560 6 FreeSans 320 0 0 0 mprj_io[28]
port 380 nsew signal bidirectional
flabel metal2 s 41713 664941 42193 664997 0 FreeSans 320 0 0 0 mprj_io_analog_en[17]
port 381 nsew signal input
flabel metal2 s 41713 663653 42193 663709 0 FreeSans 320 0 0 0 mprj_io_analog_pol[17]
port 382 nsew signal input
flabel metal2 s 41713 660617 42193 660673 0 FreeSans 320 0 0 0 mprj_io_analog_sel[17]
port 383 nsew signal input
flabel metal2 s 41713 664297 42193 664353 0 FreeSans 320 0 0 0 mprj_io_dm[51]
port 384 nsew signal input
flabel metal2 s 41713 666137 42193 666193 0 FreeSans 320 0 0 0 mprj_io_dm[52]
port 385 nsew signal input
flabel metal2 s 41713 659973 42193 660029 0 FreeSans 320 0 0 0 mprj_io_dm[53]
port 386 nsew signal input
flabel metal2 s 41713 659329 42193 659385 0 FreeSans 320 0 0 0 mprj_io_holdover[17]
port 387 nsew signal input
flabel metal2 s 41713 656293 42193 656349 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[17]
port 388 nsew signal input
flabel metal2 s 41713 663101 42193 663157 0 FreeSans 320 0 0 0 mprj_io_inp_dis[17]
port 389 nsew signal input
flabel metal2 s 41713 655649 42193 655705 0 FreeSans 320 0 0 0 mprj_io_oeb[17]
port 390 nsew signal input
flabel metal2 s 41713 658777 42193 658833 0 FreeSans 320 0 0 0 mprj_io_out[17]
port 391 nsew signal input
flabel metal2 s 41713 667977 42193 668033 0 FreeSans 320 0 0 0 mprj_io_slow_sel[17]
port 392 nsew signal input
flabel metal2 s 41713 656937 42193 656993 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[17]
port 393 nsew signal input
flabel metal2 s 41713 669817 42193 669873 0 FreeSans 320 0 0 0 mprj_io_in[17]
port 394 nsew signal tristate
flabel metal2 s 41713 655097 42193 655153 0 FreeSans 320 0 0 0 mprj_io_in_3v3[17]
port 395 nsew signal tristate
flabel metal2 s 41713 624133 42193 624189 0 FreeSans 320 0 0 0 mprj_gpio_analog[11]
port 396 nsew signal bidirectional
flabel metal2 s 41713 622293 42193 622349 0 FreeSans 320 0 0 0 mprj_gpio_noesd[11]
port 397 nsew signal bidirectional
flabel metal5 s 6598 613820 19088 626360 6 FreeSans 320 0 0 0 mprj_io[29]
port 398 nsew signal bidirectional
flabel metal2 s 41713 621741 42193 621797 0 FreeSans 320 0 0 0 mprj_io_analog_en[18]
port 399 nsew signal input
flabel metal2 s 41713 620453 42193 620509 0 FreeSans 320 0 0 0 mprj_io_analog_pol[18]
port 400 nsew signal input
flabel metal2 s 41713 617417 42193 617473 0 FreeSans 320 0 0 0 mprj_io_analog_sel[18]
port 401 nsew signal input
flabel metal2 s 41713 621097 42193 621153 0 FreeSans 320 0 0 0 mprj_io_dm[54]
port 402 nsew signal input
flabel metal2 s 41713 622937 42193 622993 0 FreeSans 320 0 0 0 mprj_io_dm[55]
port 403 nsew signal input
flabel metal2 s 41713 616773 42193 616829 0 FreeSans 320 0 0 0 mprj_io_dm[56]
port 404 nsew signal input
flabel metal2 s 41713 616129 42193 616185 0 FreeSans 320 0 0 0 mprj_io_holdover[18]
port 405 nsew signal input
flabel metal2 s 41713 613093 42193 613149 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[18]
port 406 nsew signal input
flabel metal2 s 41713 619901 42193 619957 0 FreeSans 320 0 0 0 mprj_io_inp_dis[18]
port 407 nsew signal input
flabel metal2 s 41713 612449 42193 612505 0 FreeSans 320 0 0 0 mprj_io_oeb[18]
port 408 nsew signal input
flabel metal2 s 41713 615577 42193 615633 0 FreeSans 320 0 0 0 mprj_io_out[18]
port 409 nsew signal input
flabel metal2 s 41713 624777 42193 624833 0 FreeSans 320 0 0 0 mprj_io_slow_sel[18]
port 410 nsew signal input
flabel metal2 s 41713 613737 42193 613793 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[18]
port 411 nsew signal input
flabel metal2 s 41713 626617 42193 626673 0 FreeSans 320 0 0 0 mprj_io_in[18]
port 412 nsew signal tristate
flabel metal2 s 41713 611897 42193 611953 0 FreeSans 320 0 0 0 mprj_io_in_3v3[18]
port 413 nsew signal tristate
flabel metal2 s 41713 580933 42193 580989 0 FreeSans 320 0 0 0 mprj_gpio_analog[12]
port 414 nsew signal bidirectional
flabel metal2 s 41713 579093 42193 579149 0 FreeSans 320 0 0 0 mprj_gpio_noesd[12]
port 415 nsew signal bidirectional
flabel metal5 s 6598 570620 19088 583160 6 FreeSans 320 0 0 0 mprj_io[30]
port 416 nsew signal bidirectional
flabel metal2 s 41713 578541 42193 578597 0 FreeSans 320 0 0 0 mprj_io_analog_en[19]
port 417 nsew signal input
flabel metal2 s 41713 577253 42193 577309 0 FreeSans 320 0 0 0 mprj_io_analog_pol[19]
port 418 nsew signal input
flabel metal2 s 41713 574217 42193 574273 0 FreeSans 320 0 0 0 mprj_io_analog_sel[19]
port 419 nsew signal input
flabel metal2 s 41713 577897 42193 577953 0 FreeSans 320 0 0 0 mprj_io_dm[57]
port 420 nsew signal input
flabel metal2 s 41713 579737 42193 579793 0 FreeSans 320 0 0 0 mprj_io_dm[58]
port 421 nsew signal input
flabel metal2 s 41713 573573 42193 573629 0 FreeSans 320 0 0 0 mprj_io_dm[59]
port 422 nsew signal input
flabel metal2 s 41713 572929 42193 572985 0 FreeSans 320 0 0 0 mprj_io_holdover[19]
port 423 nsew signal input
flabel metal2 s 41713 569893 42193 569949 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[19]
port 424 nsew signal input
flabel metal2 s 41713 576701 42193 576757 0 FreeSans 320 0 0 0 mprj_io_inp_dis[19]
port 425 nsew signal input
flabel metal2 s 41713 569249 42193 569305 0 FreeSans 320 0 0 0 mprj_io_oeb[19]
port 426 nsew signal input
flabel metal2 s 41713 572377 42193 572433 0 FreeSans 320 0 0 0 mprj_io_out[19]
port 427 nsew signal input
flabel metal2 s 41713 581577 42193 581633 0 FreeSans 320 0 0 0 mprj_io_slow_sel[19]
port 428 nsew signal input
flabel metal2 s 41713 570537 42193 570593 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[19]
port 429 nsew signal input
flabel metal2 s 41713 583417 42193 583473 0 FreeSans 320 0 0 0 mprj_io_in[19]
port 430 nsew signal tristate
flabel metal2 s 41713 568697 42193 568753 0 FreeSans 320 0 0 0 mprj_io_in_3v3[19]
port 431 nsew signal tristate
flabel metal2 s 41713 537733 42193 537789 0 FreeSans 320 0 0 0 mprj_gpio_analog[13]
port 432 nsew signal bidirectional
flabel metal2 s 41713 535893 42193 535949 0 FreeSans 320 0 0 0 mprj_gpio_noesd[13]
port 433 nsew signal bidirectional
flabel metal5 s 6598 527420 19088 539960 6 FreeSans 320 0 0 0 mprj_io[31]
port 434 nsew signal bidirectional
flabel metal2 s 41713 535341 42193 535397 0 FreeSans 320 0 0 0 mprj_io_analog_en[20]
port 435 nsew signal input
flabel metal2 s 41713 534053 42193 534109 0 FreeSans 320 0 0 0 mprj_io_analog_pol[20]
port 436 nsew signal input
flabel metal2 s 41713 531017 42193 531073 0 FreeSans 320 0 0 0 mprj_io_analog_sel[20]
port 437 nsew signal input
flabel metal2 s 41713 534697 42193 534753 0 FreeSans 320 0 0 0 mprj_io_dm[60]
port 438 nsew signal input
flabel metal2 s 41713 536537 42193 536593 0 FreeSans 320 0 0 0 mprj_io_dm[61]
port 439 nsew signal input
flabel metal2 s 41713 530373 42193 530429 0 FreeSans 320 0 0 0 mprj_io_dm[62]
port 440 nsew signal input
flabel metal2 s 41713 529729 42193 529785 0 FreeSans 320 0 0 0 mprj_io_holdover[20]
port 441 nsew signal input
flabel metal2 s 41713 526693 42193 526749 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[20]
port 442 nsew signal input
flabel metal2 s 41713 533501 42193 533557 0 FreeSans 320 0 0 0 mprj_io_inp_dis[20]
port 443 nsew signal input
flabel metal2 s 41713 526049 42193 526105 0 FreeSans 320 0 0 0 mprj_io_oeb[20]
port 444 nsew signal input
flabel metal2 s 41713 529177 42193 529233 0 FreeSans 320 0 0 0 mprj_io_out[20]
port 445 nsew signal input
flabel metal2 s 41713 538377 42193 538433 0 FreeSans 320 0 0 0 mprj_io_slow_sel[20]
port 446 nsew signal input
flabel metal2 s 41713 527337 42193 527393 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[20]
port 447 nsew signal input
flabel metal2 s 41713 540217 42193 540273 0 FreeSans 320 0 0 0 mprj_io_in[20]
port 448 nsew signal tristate
flabel metal2 s 41713 525497 42193 525553 0 FreeSans 320 0 0 0 mprj_io_in_3v3[20]
port 449 nsew signal tristate
flabel metal2 s 41713 410133 42193 410189 0 FreeSans 320 0 0 0 mprj_gpio_analog[14]
port 450 nsew signal bidirectional
flabel metal2 s 41713 408293 42193 408349 0 FreeSans 320 0 0 0 mprj_gpio_noesd[14]
port 451 nsew signal bidirectional
flabel metal5 s 6598 399820 19088 412360 6 FreeSans 320 0 0 0 mprj_io[32]
port 452 nsew signal bidirectional
flabel metal2 s 41713 407741 42193 407797 0 FreeSans 320 0 0 0 mprj_io_analog_en[21]
port 453 nsew signal input
flabel metal2 s 41713 406453 42193 406509 0 FreeSans 320 0 0 0 mprj_io_analog_pol[21]
port 454 nsew signal input
flabel metal2 s 41713 403417 42193 403473 0 FreeSans 320 0 0 0 mprj_io_analog_sel[21]
port 455 nsew signal input
flabel metal2 s 41713 407097 42193 407153 0 FreeSans 320 0 0 0 mprj_io_dm[63]
port 456 nsew signal input
flabel metal2 s 41713 408937 42193 408993 0 FreeSans 320 0 0 0 mprj_io_dm[64]
port 457 nsew signal input
flabel metal2 s 41713 402773 42193 402829 0 FreeSans 320 0 0 0 mprj_io_dm[65]
port 458 nsew signal input
flabel metal2 s 41713 402129 42193 402185 0 FreeSans 320 0 0 0 mprj_io_holdover[21]
port 459 nsew signal input
flabel metal2 s 41713 399093 42193 399149 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[21]
port 460 nsew signal input
flabel metal2 s 41713 405901 42193 405957 0 FreeSans 320 0 0 0 mprj_io_inp_dis[21]
port 461 nsew signal input
flabel metal2 s 41713 398449 42193 398505 0 FreeSans 320 0 0 0 mprj_io_oeb[21]
port 462 nsew signal input
flabel metal2 s 41713 401577 42193 401633 0 FreeSans 320 0 0 0 mprj_io_out[21]
port 463 nsew signal input
flabel metal2 s 41713 410777 42193 410833 0 FreeSans 320 0 0 0 mprj_io_slow_sel[21]
port 464 nsew signal input
flabel metal2 s 41713 399737 42193 399793 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[21]
port 465 nsew signal input
flabel metal2 s 41713 412617 42193 412673 0 FreeSans 320 0 0 0 mprj_io_in[21]
port 466 nsew signal tristate
flabel metal2 s 41713 397897 42193 397953 0 FreeSans 320 0 0 0 mprj_io_in_3v3[21]
port 467 nsew signal tristate
flabel metal2 s 41713 366933 42193 366989 0 FreeSans 320 0 0 0 mprj_gpio_analog[15]
port 468 nsew signal bidirectional
flabel metal2 s 41713 365093 42193 365149 0 FreeSans 320 0 0 0 mprj_gpio_noesd[15]
port 469 nsew signal bidirectional
flabel metal5 s 6598 356620 19088 369160 6 FreeSans 320 0 0 0 mprj_io[33]
port 470 nsew signal bidirectional
flabel metal2 s 41713 364541 42193 364597 0 FreeSans 320 0 0 0 mprj_io_analog_en[22]
port 471 nsew signal input
flabel metal2 s 41713 363253 42193 363309 0 FreeSans 320 0 0 0 mprj_io_analog_pol[22]
port 472 nsew signal input
flabel metal2 s 41713 360217 42193 360273 0 FreeSans 320 0 0 0 mprj_io_analog_sel[22]
port 473 nsew signal input
flabel metal2 s 41713 363897 42193 363953 0 FreeSans 320 0 0 0 mprj_io_dm[66]
port 474 nsew signal input
flabel metal2 s 41713 365737 42193 365793 0 FreeSans 320 0 0 0 mprj_io_dm[67]
port 475 nsew signal input
flabel metal2 s 41713 359573 42193 359629 0 FreeSans 320 0 0 0 mprj_io_dm[68]
port 476 nsew signal input
flabel metal2 s 41713 358929 42193 358985 0 FreeSans 320 0 0 0 mprj_io_holdover[22]
port 477 nsew signal input
flabel metal2 s 41713 355893 42193 355949 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[22]
port 478 nsew signal input
flabel metal2 s 41713 362701 42193 362757 0 FreeSans 320 0 0 0 mprj_io_inp_dis[22]
port 479 nsew signal input
flabel metal2 s 41713 355249 42193 355305 0 FreeSans 320 0 0 0 mprj_io_oeb[22]
port 480 nsew signal input
flabel metal2 s 41713 358377 42193 358433 0 FreeSans 320 0 0 0 mprj_io_out[22]
port 481 nsew signal input
flabel metal2 s 41713 367577 42193 367633 0 FreeSans 320 0 0 0 mprj_io_slow_sel[22]
port 482 nsew signal input
flabel metal2 s 41713 356537 42193 356593 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[22]
port 483 nsew signal input
flabel metal2 s 41713 369417 42193 369473 0 FreeSans 320 0 0 0 mprj_io_in[22]
port 484 nsew signal tristate
flabel metal2 s 41713 354697 42193 354753 0 FreeSans 320 0 0 0 mprj_io_in_3v3[22]
port 485 nsew signal tristate
flabel metal2 s 41713 323733 42193 323789 0 FreeSans 320 0 0 0 mprj_gpio_analog[16]
port 486 nsew signal bidirectional
flabel metal2 s 41713 321893 42193 321949 0 FreeSans 320 0 0 0 mprj_gpio_noesd[16]
port 487 nsew signal bidirectional
flabel metal5 s 6598 313420 19088 325960 6 FreeSans 320 0 0 0 mprj_io[34]
port 488 nsew signal bidirectional
flabel metal2 s 41713 321341 42193 321397 0 FreeSans 320 0 0 0 mprj_io_analog_en[23]
port 489 nsew signal input
flabel metal2 s 41713 320053 42193 320109 0 FreeSans 320 0 0 0 mprj_io_analog_pol[23]
port 490 nsew signal input
flabel metal2 s 41713 317017 42193 317073 0 FreeSans 320 0 0 0 mprj_io_analog_sel[23]
port 491 nsew signal input
flabel metal2 s 41713 320697 42193 320753 0 FreeSans 320 0 0 0 mprj_io_dm[69]
port 492 nsew signal input
flabel metal2 s 41713 322537 42193 322593 0 FreeSans 320 0 0 0 mprj_io_dm[70]
port 493 nsew signal input
flabel metal2 s 41713 316373 42193 316429 0 FreeSans 320 0 0 0 mprj_io_dm[71]
port 494 nsew signal input
flabel metal2 s 41713 315729 42193 315785 0 FreeSans 320 0 0 0 mprj_io_holdover[23]
port 495 nsew signal input
flabel metal2 s 41713 312693 42193 312749 0 FreeSans 320 0 0 0 mprj_io_ib_mode_sel[23]
port 496 nsew signal input
flabel metal2 s 41713 319501 42193 319557 0 FreeSans 320 0 0 0 mprj_io_inp_dis[23]
port 497 nsew signal input
flabel metal2 s 41713 312049 42193 312105 0 FreeSans 320 0 0 0 mprj_io_oeb[23]
port 498 nsew signal input
flabel metal2 s 41713 315177 42193 315233 0 FreeSans 320 0 0 0 mprj_io_out[23]
port 499 nsew signal input
flabel metal2 s 41713 324377 42193 324433 0 FreeSans 320 0 0 0 mprj_io_slow_sel[23]
port 500 nsew signal input
flabel metal2 s 41713 313337 42193 313393 0 FreeSans 320 0 0 0 mprj_io_vtrip_sel[23]
port 501 nsew signal input
flabel metal2 s 41713 326217 42193 326273 0 FreeSans 320 0 0 0 mprj_io_in[23]
port 502 nsew signal tristate
flabel metal2 s 41713 311497 42193 311553 0 FreeSans 320 0 0 0 mprj_io_in_3v3[23]
port 503 nsew signal tristate
flabel metal5 s 136713 7143 144149 18309 6 FreeSans 320 0 0 0 resetb
port 505 nsew signal input
flabel metal4 s 132600 36323 132792 37013 6 FreeSans 320 0 0 0 vdda
port 507 nsew signal bidirectional
flabel metal5 s 628410 1018624 640578 1030788 6 FreeSans 320 0 0 0 mprj_io[15]
port 511 nsew signal bidirectional
flabel metal5 s 526610 1018624 538778 1030788 6 FreeSans 320 0 0 0 mprj_io[16]
port 513 nsew signal bidirectional
flabel metal5 s 475210 1018624 487378 1030788 6 FreeSans 320 0 0 0 mprj_io[17]
port 515 nsew signal bidirectional
flabel metal5 s 697980 909666 711432 920546 6 FreeSans 320 0 0 0 vccd1_pad
port 522 nsew signal bidirectional
flabel metal5 s 698624 819822 710788 831990 6 FreeSans 320 0 0 0 vdda1_pad
port 523 nsew signal bidirectional
flabel metal5 s 698624 505222 710788 517390 6 FreeSans 320 0 0 0 vdda1_pad2
port 524 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030788 6 FreeSans 320 0 0 0 vssa1_pad
port 525 nsew signal bidirectional
flabel metal5 s 698624 417022 710788 429190 6 FreeSans 320 0 0 0 vssa1_pad2
port 526 nsew signal bidirectional
flabel metal4 s 680587 459800 681277 459992 6 FreeSans 320 0 0 0 vdda1
port 528 nsew signal bidirectional
flabel metal4 s 688881 459800 688947 474800 6 FreeSans 320 0 0 0 vssa1
port 529 nsew signal bidirectional
flabel metal5 s 697980 461866 711432 472746 6 FreeSans 320 0 0 0 vssd1_pad
port 531 nsew signal bidirectional
flabel metal3 s 184944 997600 189944 1014070 6 FreeSans 320 0 0 0 mprj_analog[7]
port 532 nsew signal bidirectional
flabel metal5 s 181410 1018624 193578 1030788 6 FreeSans 320 0 0 0 mprj_io[21]
port 533 nsew signal bidirectional
flabel metal3 s 133544 997600 138544 1014070 6 FreeSans 320 0 0 0 mprj_analog[8]
port 534 nsew signal bidirectional
flabel metal5 s 130010 1018624 142178 1030788 6 FreeSans 320 0 0 0 mprj_io[22]
port 535 nsew signal bidirectional
flabel metal3 s 82144 997600 87144 1014070 6 FreeSans 320 0 0 0 mprj_analog[9]
port 536 nsew signal bidirectional
flabel metal5 s 78610 1018624 90778 1030788 6 FreeSans 320 0 0 0 mprj_io[23]
port 537 nsew signal bidirectional
flabel metal3 s 23530 960144 40000 965144 6 FreeSans 320 0 0 0 mprj_analog[10]
port 538 nsew signal bidirectional
flabel metal5 s 6811 956610 18975 968778 6 FreeSans 320 0 0 0 mprj_io[24]
port 539 nsew signal bidirectional
flabel metal3 s 240478 997600 254800 1000736 6 FreeSans 320 0 0 0 mprj_analog[6]
port 544 nsew signal bidirectional
flabel metal2 s 240478 997600 245258 1002732 6 FreeSans 320 0 0 0 mprj_clamp_high[2]
port 545 nsew signal input
flabel metal2 s 230499 997600 235279 998010 6 FreeSans 320 0 0 0 mprj_clamp_low[2]
port 546 nsew signal input
flabel metal5 s 231810 1018624 243978 1030788 6 FreeSans 320 0 0 0 mprj_io[20]
port 547 nsew signal bidirectional
flabel metal5 s 6167 914054 19619 924934 6 FreeSans 320 0 0 0 vccd2_pad
port 548 nsew signal bidirectional
flabel metal5 s 6811 484410 18975 496578 6 FreeSans 320 0 0 0 vdda2_pad
port 549 nsew signal bidirectional
flabel metal5 s 6811 829010 18975 841178 6 FreeSans 320 0 0 0 vssa2_pad
port 550 nsew signal bidirectional
flabel metal4 s 36323 455607 37013 455799 6 FreeSans 320 0 0 0 vdda2
port 553 nsew signal bidirectional
flabel metal4 s 28653 440800 28719 455800 6 FreeSans 320 0 0 0 vssa2
port 555 nsew signal bidirectional
flabel metal5 s 6167 442854 19619 453734 6 FreeSans 320 0 0 0 vssd2_pad
port 557 nsew signal bidirectional
flabel metal5 s 386210 1018624 398378 1030788 6 FreeSans 320 0 0 0 mprj_io[18]
port 521 nsew signal bidirectional
flabel metal5 s 284410 1018624 296578 1030788 6 FreeSans 320 0 0 0 mprj_io[19]
port 543 nsew signal bidirectional
flabel metal5 s 698624 953022 710788 965190 6 FreeSans 320 0 0 0 mprj_io[14]
port 517 nsew signal bidirectional
flabel metal3 s 293078 997600 307400 1000736 6 FreeSans 320 0 0 0 mprj_analog[5]
port 540 nsew signal bidirectional
flabel metal2 s 293078 997600 297858 1002732 6 FreeSans 320 0 0 0 mprj_clamp_high[1]
port 541 nsew signal input
flabel metal2 s 283099 997600 287879 998010 6 FreeSans 320 0 0 0 mprj_clamp_low[1]
port 542 nsew signal input
flabel metal3 s 394878 997600 409200 1000736 6 FreeSans 320 0 0 0 mprj_analog[4]
port 518 nsew signal bidirectional
flabel metal2 s 394878 997600 399658 1002732 6 FreeSans 320 0 0 0 mprj_clamp_high[0]
port 519 nsew signal input
flabel metal2 s 384899 997600 389679 998010 6 FreeSans 320 0 0 0 mprj_clamp_low[0]
port 520 nsew signal input
flabel metal2 141667 39934 141813 40000 0 FreeSans 320 0 0 0 resetb_core_h
port 506 nsew signal tristate
flabel metal5 44276 178502 46712 179254 0 FreeSans 3200 0 0 0 vccd2
port 552 nsew signal bidirectional
flabel metal5 41056 178502 43492 179254 0 FreeSans 3200 0 0 0 vssd2
port 556 nsew signal bidirectional
flabel metal5 674150 134670 676514 135366 0 FreeSans 3200 0 0 0 vccd1
port 527 nsew signal bidirectional
flabel metal5 670936 134790 673300 135486 0 FreeSans 3200 0 0 0 vssd1
port 530 nsew signal bidirectional
flabel metal3 s 677600 956656 694070 961656 6 FreeSans 320 0 0 0 mprj_analog[0]
port 516 nsew signal bidirectional
flabel metal3 s 631944 997600 636944 1014070 6 FreeSans 320 0 0 0 mprj_analog[1]
port 510 nsew signal bidirectional
flabel metal3 s 530144 997600 535144 1014070 6 FreeSans 320 0 0 0 mprj_analog[2]
port 512 nsew signal bidirectional
flabel metal3 s 478744 997600 483744 1014070 6 FreeSans 320 0 0 0 mprj_analog[3]
port 514 nsew signal bidirectional
flabel metal2 s 521843 41713 521899 42193 0 FreeSans 320 90 0 0 gpio_inenb_core
port 23 nsew signal input
flabel metal2 310095 41713 310151 42193 0 FreeSans 320 90 0 0 flash_csb_oeb_core
port 563 nsew signal input
flabel metal2 361767 41713 361823 42193 0 FreeSans 320 90 0 0 flash_clk_core
port 562 nsew signal input
flabel metal2 364895 41713 364951 42193 0 FreeSans 320 90 0 0 flash_clk_oeb_core
port 561 nsew signal input
flabel metal2 306967 41713 307023 42193 0 FreeSans 320 90 0 0 flash_csb_core
port 559 nsew signal input
flabel metal2 s 529295 41713 529351 42193 0 FreeSans 320 90 0 0 gpio_outenb_core
port 27 nsew signal input
flabel metal2 s 526167 41713 526223 42193 0 FreeSans 320 90 0 0 gpio_out_core
port 26 nsew signal input
flabel metal2 s 520647 41713 520703 42193 0 FreeSans 320 90 0 0 gpio_mode0_core
port 24 nsew signal input
flabel metal2 s 515127 41713 515183 42193 0 FreeSans 320 90 0 0 gpio_in_core
port 22 nsew signal tristate
flabel metal2 s 474495 41713 474551 42193 0 FreeSans 320 90 0 0 flash_io1_oeb_core
port 20 nsew signal input
flabel metal2 s 467043 41713 467099 42193 0 FreeSans 320 90 0 0 flash_io1_ieb_core
port 19 nsew signal input
flabel metal2 s 471367 41713 471423 42193 0 FreeSans 320 90 0 0 flash_io1_do_core
port 18 nsew signal input
flabel metal2 s 460327 41713 460383 42193 0 FreeSans 320 90 0 0 flash_io1_di_core
port 17 nsew signal tristate
flabel metal2 s 419695 41713 419751 42193 0 FreeSans 320 90 0 0 flash_io0_oeb_core
port 15 nsew signal input
flabel metal2 s 412243 41713 412299 42193 0 FreeSans 320 90 0 0 flash_io0_ieb_core
port 14 nsew signal input
flabel metal2 s 416567 41713 416623 42193 0 FreeSans 320 90 0 0 flash_io0_do_core
port 13 nsew signal input
flabel metal2 s 405527 41713 405583 42193 0 FreeSans 320 90 0 0 flash_io0_di_core
port 12 nsew signal tristate
flabel metal2 s 194043 41713 194099 42193 0 FreeSans 320 90 0 0 por
port 2 nsew signal input
flabel metal2 s 187327 41713 187383 42193 0 FreeSans 320 90 0 0 clock_core
port 1 nsew signal tristate
rlabel metal3 140494 40139 140494 40139 1 xresloop
rlabel metal1 142538 40056 142538 40056 1 xres_vss_loop
flabel metal2 s 524971 41746 525027 42226 0 FreeSans 320 90 0 0 gpio_mode1_core
port 592 nsew signal input
flabel metal2 675407 102123 675887 102179 0 FreeSans 320 0 0 0 mprj_io_one[0]
port 564 nsew
flabel metal2 675407 147323 675887 147379 0 FreeSans 320 0 0 0 mprj_io_one[1]
port 565 nsew
flabel metal2 675407 192323 675887 192379 0 FreeSans 320 0 0 0 mprj_io_one[2]
port 566 nsew
flabel metal2 675407 237523 675887 237579 0 FreeSans 320 0 0 0 mprj_io_one[3]
port 567 nsew
flabel metal2 675407 282523 675887 282579 0 FreeSans 320 0 0 0 mprj_io_one[4]
port 568 nsew
flabel metal2 675407 327523 675887 327579 0 FreeSans 320 0 0 0 mprj_io_one[5]
port 569 nsew
flabel metal2 675407 372723 675887 372779 0 FreeSans 320 0 0 0 mprj_io_one[6]
port 570 nsew
flabel metal2 675407 549923 675887 549979 0 FreeSans 320 0 0 0 mprj_io_one[7]
port 571 nsew
flabel metal2 675407 595123 675887 595179 0 FreeSans 320 0 0 0 mprj_io_one[8]
port 572 nsew
flabel metal2 675407 640123 675887 640179 0 FreeSans 320 0 0 0 mprj_io_one[9]
port 573 nsew
flabel metal2 675407 685323 675887 685379 0 FreeSans 320 0 0 0 mprj_io_one[10]
port 574 nsew
flabel metal2 675407 730323 675887 730379 0 FreeSans 320 0 0 0 mprj_io_one[11]
port 575 nsew
flabel metal2 675407 775323 675887 775379 0 FreeSans 320 0 0 0 mprj_io_one[12]
port 576 nsew
flabel metal2 675407 864523 675887 864579 0 FreeSans 320 0 0 0 mprj_io_one[13]
port 577 nsew
flabel metal2 41713 798221 42193 798277 0 FreeSans 320 0 0 0 mprj_io_one[14]
port 578 nsew
flabel metal2 41713 755021 42193 755077 0 FreeSans 320 0 0 0 mprj_io_one[15]
port 579 nsew
flabel metal2 41713 711821 42193 711877 0 FreeSans 320 0 0 0 mprj_io_one[16]
port 580 nsew
flabel metal2 41713 668621 42193 668677 0 FreeSans 320 0 0 0 mprj_io_one[17]
port 581 nsew
flabel metal2 41713 625421 42193 625477 0 FreeSans 320 0 0 0 mprj_io_one[18]
port 582 nsew
flabel metal2 41713 582221 42193 582277 0 FreeSans 320 0 0 0 mprj_io_one[19]
port 583 nsew
flabel metal2 41713 539021 42193 539077 0 FreeSans 320 0 0 0 mprj_io_one[20]
port 584 nsew
flabel metal2 41713 411421 42193 411477 0 FreeSans 320 0 0 0 mprj_io_one[21]
port 585 nsew
flabel metal2 41713 368221 42193 368277 0 FreeSans 320 0 0 0 mprj_io_one[22]
port 586 nsew
flabel metal2 41713 325021 42193 325077 0 FreeSans 320 0 0 0 mprj_io_one[23]
port 587 nsew
flabel metal2 41713 281821 42193 281877 0 FreeSans 320 0 0 0 mprj_io_one[24]
port 588 nsew
flabel metal2 41713 238621 42193 238677 0 FreeSans 320 0 0 0 mprj_io_one[25]
port 589 nsew
flabel metal2 41713 195421 42193 195477 0 FreeSans 320 0 0 0 mprj_io_one[26]
port 590 nsew
flabel metal2 308255 41746 308311 42226 0 FreeSans 320 90 0 0 porb_h
port 591 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
